VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 1.500 -3.500 ;
  SIZE 191.790 BY 435.000 ;
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.000 10.155 159.520 10.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 16.295 159.520 16.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 22.435 159.520 23.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 28.575 159.520 29.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 34.715 159.520 35.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 40.855 159.520 41.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 46.995 159.520 47.695 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 53.135 159.520 53.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 59.275 159.520 59.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 65.415 159.520 66.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 71.555 159.520 72.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 77.695 159.520 78.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 83.835 159.520 84.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 89.975 159.520 90.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 96.115 159.520 96.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 102.255 159.520 102.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 108.395 159.520 109.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 114.535 159.520 115.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 120.675 159.520 121.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 126.815 159.520 127.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 132.955 159.520 133.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 139.095 159.520 139.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 145.235 159.520 145.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 151.375 159.520 152.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 157.515 159.520 158.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 163.655 159.520 164.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 169.795 159.520 170.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 175.935 159.520 176.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 182.075 159.520 182.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 188.215 159.520 188.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 194.355 159.520 195.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 200.495 159.520 201.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 206.635 159.520 207.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 212.775 159.520 213.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 218.915 159.520 219.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 225.055 159.520 225.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 231.195 159.520 231.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 237.335 159.520 238.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 243.475 159.520 244.175 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 249.615 159.520 250.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 255.755 159.520 256.455 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 261.895 159.520 262.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 268.035 159.520 268.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 274.175 159.520 274.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 280.315 159.520 281.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 286.455 159.520 287.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 292.595 159.520 293.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 298.735 159.520 299.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 304.875 159.520 305.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 311.015 159.520 311.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 317.155 159.520 317.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 323.295 159.520 323.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 329.435 159.520 330.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 335.575 159.520 336.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 341.715 159.520 342.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 347.855 159.520 348.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 353.995 159.520 354.695 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 360.135 159.520 360.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 366.275 159.520 366.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 372.415 159.520 373.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 378.555 159.520 379.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 384.695 159.520 385.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 390.835 159.520 391.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 396.975 159.520 397.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 406.915 159.520 407.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 428.615 188.875 430.115 ;
    END
  END VDDA
  PIN VSSA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.000 6.705 159.520 7.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 12.845 159.520 13.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 18.985 159.520 19.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 25.125 159.520 25.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 31.265 159.520 31.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 37.405 159.520 38.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 43.545 159.520 44.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 49.685 159.520 50.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 55.825 159.520 56.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 61.965 159.520 62.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 68.105 159.520 68.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 74.245 159.520 74.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 80.385 159.520 81.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 86.525 159.520 87.225 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 92.665 159.520 93.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 98.805 159.520 99.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 104.945 159.520 105.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 111.085 159.520 111.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 117.225 159.520 117.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 123.365 159.520 124.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 129.505 159.520 130.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 135.645 159.520 136.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 141.785 159.520 142.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 147.925 159.520 148.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 154.065 159.520 154.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 160.205 159.520 160.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 166.345 159.520 167.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 172.485 159.520 173.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 178.625 159.520 179.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 184.765 159.520 185.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 190.905 159.520 191.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 197.045 159.520 197.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 203.185 159.520 203.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 209.325 159.520 210.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 215.465 159.520 216.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 221.605 159.520 222.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 227.745 159.520 228.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 233.885 159.520 234.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 240.025 159.520 240.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 246.165 159.520 246.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 252.305 159.520 253.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 258.445 159.520 259.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 264.585 159.520 265.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 270.725 159.520 271.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 276.865 159.520 277.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 283.005 159.520 283.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 289.145 159.520 289.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 295.285 159.520 295.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 301.425 159.520 302.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 307.565 159.520 308.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 313.705 159.520 314.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 319.845 159.520 320.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 325.985 159.520 326.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 332.125 159.520 332.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 338.265 159.520 338.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 344.405 159.520 345.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 350.545 159.520 351.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 356.685 159.520 357.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 362.825 159.520 363.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 368.965 159.520 369.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 375.105 159.520 375.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 381.245 159.520 381.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 387.385 159.520 388.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 393.525 159.520 394.225 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.000 412.565 159.520 414.065 ;
    END
  END VSSA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.000 400.265 159.520 400.765 ;
    END
  END VCCD
  PIN VSSD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.000 402.565 159.520 403.065 ;
    END
  END VSSD
  PIN VREFH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -2.600 5.000 3.500 5.500 ;
    END
  END VREFH
  PIN Din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.210 408.645 8.410 439.300 ;
    END
  END Din0[0]
  PIN Din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.900 409.095 9.100 439.300 ;
    END
  END Din0[1]
  PIN Din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.580 409.545 9.780 439.300 ;
    END
  END Din0[2]
  PIN Din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.250 409.995 10.450 439.300 ;
    END
  END Din0[3]
  PIN Din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.910 410.455 11.110 439.300 ;
    END
  END Din0[4]
  PIN Din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.570 410.955 11.770 439.300 ;
    END
  END Din0[5]
  PIN Din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.230 411.445 12.430 439.300 ;
    END
  END Din0[6]
  PIN Din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.900 411.985 13.100 439.300 ;
    END
  END Din0[7]
  PIN VOUT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.040 431.140 37.280 439.300 ;
    END
  END VOUT0
  PIN Din1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.840 408.645 47.040 439.300 ;
    END
  END Din1[0]
  PIN Din1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.530 409.095 47.730 439.300 ;
    END
  END Din1[1]
  PIN Din1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.210 409.545 48.410 439.300 ;
    END
  END Din1[2]
  PIN Din1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.880 409.995 49.080 439.300 ;
    END
  END Din1[3]
  PIN Din1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.540 410.455 49.740 439.300 ;
    END
  END Din1[4]
  PIN Din1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.200 410.955 50.400 439.300 ;
    END
  END Din1[5]
  PIN Din1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.860 411.445 51.060 439.300 ;
    END
  END Din1[6]
  PIN Din1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.530 411.985 51.730 439.300 ;
    END
  END Din1[7]
  PIN VOUT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.670 419.115 75.910 439.300 ;
    END
  END VOUT1
  PIN Din2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.470 408.645 85.670 439.300 ;
    END
  END Din2[0]
  PIN Din2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.160 409.095 86.360 439.300 ;
    END
  END Din2[1]
  PIN Din2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.840 409.545 87.040 439.300 ;
    END
  END Din2[2]
  PIN Din2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.510 409.995 87.710 439.300 ;
    END
  END Din2[3]
  PIN Din2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.170 410.455 88.370 439.300 ;
    END
  END Din2[4]
  PIN Din2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.830 410.955 89.030 439.300 ;
    END
  END Din2[5]
  PIN Din2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.490 411.445 89.690 439.300 ;
    END
  END Din2[6]
  PIN Din2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.160 411.985 90.360 439.300 ;
    END
  END Din2[7]
  PIN VOUT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.300 419.115 114.540 439.300 ;
    END
  END VOUT2
  PIN Din3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.100 408.645 124.300 439.300 ;
    END
  END Din3[0]
  PIN Din3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.790 409.095 124.990 439.300 ;
    END
  END Din3[1]
  PIN Din3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.470 409.545 125.670 439.300 ;
    END
  END Din3[2]
  PIN Din3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.140 409.995 126.340 439.300 ;
    END
  END Din3[3]
  PIN Din3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.800 410.455 127.000 439.300 ;
    END
  END Din3[4]
  PIN Din3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.460 410.955 127.660 439.300 ;
    END
  END Din3[5]
  PIN Din3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.120 411.445 128.320 439.300 ;
    END
  END Din3[6]
  PIN Din3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.790 411.985 128.990 439.300 ;
    END
  END Din3[7]
  PIN VOUT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.930 419.115 153.170 439.300 ;
    END
  END VOUT3
  PIN SAMPLE0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.390 432.435 161.560 439.300 ;
    END
  END SAMPLE0
  PIN RESULT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.140 433.430 165.310 439.300 ;
    END
  END RESULT0
  PIN PIN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.655 427.620 166.825 439.300 ;
    END
  END PIN0
  PIN SEL0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.570 426.945 167.740 439.300 ;
    END
  END SEL0
  PIN RESULT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.450 433.835 173.620 439.300 ;
    END
  END RESULT1
  PIN PIN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.110 427.620 174.280 439.300 ;
    END
  END PIN1
  PIN SEL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.010 426.945 175.180 439.300 ;
    END
  END SEL1
  PIN SAMPLE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.890 432.670 176.060 439.300 ;
    END
  END SAMPLE1
  PIN RESULT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.700 433.345 179.870 439.300 ;
    END
  END RESULT2
  PIN SAMPLE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.590 433.375 180.760 439.300 ;
    END
  END SAMPLE2
  PIN PIN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.645 427.620 181.815 439.300 ;
    END
  END PIN2
  PIN SEL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.490 426.945 182.660 439.300 ;
    END
  END SEL2
  PIN RESULT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.440 432.485 186.610 439.300 ;
    END
  END RESULT3
  PIN SAMPLE3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.520 432.320 187.690 439.300 ;
    END
  END SAMPLE3
  PIN PIN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.490 427.620 188.660 439.300 ;
    END
  END PIN3
  PIN SEL3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.415 426.945 189.585 439.300 ;
    END
  END SEL3
  OBS
      LAYER li1 ;
        RECT 7.710 6.210 188.065 437.895 ;
      LAYER met1 ;
        RECT 3.470 5.000 188.735 437.970 ;
      LAYER met2 ;
        RECT 3.500 408.365 7.930 437.940 ;
        RECT 13.380 430.860 36.760 437.940 ;
        RECT 37.560 430.860 46.560 437.940 ;
        RECT 13.380 411.705 46.560 430.860 ;
        RECT 52.010 418.835 75.390 437.940 ;
        RECT 76.190 418.835 85.190 437.940 ;
        RECT 52.010 411.705 85.190 418.835 ;
        RECT 90.640 418.835 114.020 437.940 ;
        RECT 114.820 418.835 123.820 437.940 ;
        RECT 90.640 411.705 123.820 418.835 ;
        RECT 129.270 418.835 152.650 437.940 ;
        RECT 153.450 432.155 161.110 437.940 ;
        RECT 161.840 433.150 164.860 437.940 ;
        RECT 165.590 433.150 166.375 437.940 ;
        RECT 161.840 432.155 166.375 433.150 ;
        RECT 153.450 427.340 166.375 432.155 ;
        RECT 167.105 427.340 167.290 437.940 ;
        RECT 153.450 426.665 167.290 427.340 ;
        RECT 168.020 433.555 173.170 437.940 ;
        RECT 168.020 427.340 173.830 433.555 ;
        RECT 174.560 427.340 174.730 437.940 ;
        RECT 168.020 426.665 174.730 427.340 ;
        RECT 175.460 432.390 175.610 437.940 ;
        RECT 176.340 433.065 179.420 437.940 ;
        RECT 180.150 433.095 180.310 437.940 ;
        RECT 181.040 433.095 181.365 437.940 ;
        RECT 180.150 433.065 181.365 433.095 ;
        RECT 176.340 432.390 181.365 433.065 ;
        RECT 175.460 427.340 181.365 432.390 ;
        RECT 182.095 427.340 182.210 437.940 ;
        RECT 175.460 426.665 182.210 427.340 ;
        RECT 182.940 432.205 186.160 437.940 ;
        RECT 186.890 432.205 187.240 437.940 ;
        RECT 182.940 432.040 187.240 432.205 ;
        RECT 187.970 432.040 188.210 437.940 ;
        RECT 182.940 427.340 188.210 432.040 ;
        RECT 188.940 427.340 189.135 437.940 ;
        RECT 182.940 426.665 189.135 427.340 ;
        RECT 153.450 418.835 189.415 426.665 ;
        RECT 129.270 411.705 189.415 418.835 ;
        RECT 12.710 411.165 46.560 411.705 ;
        RECT 51.340 411.165 85.190 411.705 ;
        RECT 89.970 411.165 123.820 411.705 ;
        RECT 128.600 411.165 189.415 411.705 ;
        RECT 12.050 410.675 46.560 411.165 ;
        RECT 50.680 410.675 85.190 411.165 ;
        RECT 89.310 410.675 123.820 411.165 ;
        RECT 127.940 410.675 189.415 411.165 ;
        RECT 11.390 410.175 46.560 410.675 ;
        RECT 50.020 410.175 85.190 410.675 ;
        RECT 88.650 410.175 123.820 410.675 ;
        RECT 127.280 410.175 189.415 410.675 ;
        RECT 10.730 409.715 46.560 410.175 ;
        RECT 49.360 409.715 85.190 410.175 ;
        RECT 87.990 409.715 123.820 410.175 ;
        RECT 126.620 409.715 189.415 410.175 ;
        RECT 10.060 409.265 46.560 409.715 ;
        RECT 48.690 409.265 85.190 409.715 ;
        RECT 87.320 409.265 123.820 409.715 ;
        RECT 125.950 409.265 189.415 409.715 ;
        RECT 9.380 408.815 46.560 409.265 ;
        RECT 48.010 408.815 85.190 409.265 ;
        RECT 86.640 408.815 123.820 409.265 ;
        RECT 125.270 408.815 189.415 409.265 ;
        RECT 8.690 408.365 46.560 408.815 ;
        RECT 47.320 408.365 85.190 408.815 ;
        RECT 85.950 408.365 123.820 408.815 ;
        RECT 124.580 408.365 189.415 408.815 ;
        RECT 3.500 5.780 189.415 408.365 ;
        RECT 3.780 4.970 189.415 5.780 ;
      LAYER met3 ;
        RECT 14.635 430.515 189.690 436.370 ;
        RECT 189.275 428.215 189.690 430.515 ;
        RECT 14.635 414.465 189.690 428.215 ;
        RECT 159.920 412.165 189.690 414.465 ;
        RECT 14.635 407.815 189.690 412.165 ;
        RECT 159.920 406.515 189.690 407.815 ;
        RECT 14.635 403.465 189.690 406.515 ;
        RECT 159.920 402.165 189.690 403.465 ;
        RECT 14.635 401.165 189.690 402.165 ;
        RECT 159.920 399.865 189.690 401.165 ;
        RECT 14.635 398.075 189.690 399.865 ;
        RECT 159.920 396.575 189.690 398.075 ;
        RECT 14.635 394.625 189.690 396.575 ;
        RECT 159.920 393.125 189.690 394.625 ;
        RECT 14.635 391.935 189.690 393.125 ;
        RECT 159.920 390.435 189.690 391.935 ;
        RECT 14.635 388.485 189.690 390.435 ;
        RECT 159.920 386.985 189.690 388.485 ;
        RECT 14.635 385.795 189.690 386.985 ;
        RECT 159.920 384.295 189.690 385.795 ;
        RECT 14.635 382.345 189.690 384.295 ;
        RECT 159.920 380.845 189.690 382.345 ;
        RECT 14.635 379.655 189.690 380.845 ;
        RECT 159.920 378.155 189.690 379.655 ;
        RECT 14.635 376.205 189.690 378.155 ;
        RECT 159.920 374.705 189.690 376.205 ;
        RECT 14.635 373.515 189.690 374.705 ;
        RECT 159.920 372.015 189.690 373.515 ;
        RECT 14.635 370.065 189.690 372.015 ;
        RECT 159.920 368.565 189.690 370.065 ;
        RECT 14.635 367.375 189.690 368.565 ;
        RECT 159.920 365.875 189.690 367.375 ;
        RECT 14.635 363.925 189.690 365.875 ;
        RECT 159.920 362.425 189.690 363.925 ;
        RECT 14.635 361.235 189.690 362.425 ;
        RECT 159.920 359.735 189.690 361.235 ;
        RECT 14.635 357.785 189.690 359.735 ;
        RECT 159.920 356.285 189.690 357.785 ;
        RECT 14.635 355.095 189.690 356.285 ;
        RECT 159.920 353.595 189.690 355.095 ;
        RECT 14.635 351.645 189.690 353.595 ;
        RECT 159.920 350.145 189.690 351.645 ;
        RECT 14.635 348.955 189.690 350.145 ;
        RECT 159.920 347.455 189.690 348.955 ;
        RECT 14.635 345.505 189.690 347.455 ;
        RECT 159.920 344.005 189.690 345.505 ;
        RECT 14.635 342.815 189.690 344.005 ;
        RECT 159.920 341.315 189.690 342.815 ;
        RECT 14.635 339.365 189.690 341.315 ;
        RECT 159.920 337.865 189.690 339.365 ;
        RECT 14.635 336.675 189.690 337.865 ;
        RECT 159.920 335.175 189.690 336.675 ;
        RECT 14.635 333.225 189.690 335.175 ;
        RECT 159.920 331.725 189.690 333.225 ;
        RECT 14.635 330.535 189.690 331.725 ;
        RECT 159.920 329.035 189.690 330.535 ;
        RECT 14.635 327.085 189.690 329.035 ;
        RECT 159.920 325.585 189.690 327.085 ;
        RECT 14.635 324.395 189.690 325.585 ;
        RECT 159.920 322.895 189.690 324.395 ;
        RECT 14.635 320.945 189.690 322.895 ;
        RECT 159.920 319.445 189.690 320.945 ;
        RECT 14.635 318.255 189.690 319.445 ;
        RECT 159.920 316.755 189.690 318.255 ;
        RECT 14.635 314.805 189.690 316.755 ;
        RECT 159.920 313.305 189.690 314.805 ;
        RECT 14.635 312.115 189.690 313.305 ;
        RECT 159.920 310.615 189.690 312.115 ;
        RECT 14.635 308.665 189.690 310.615 ;
        RECT 159.920 307.165 189.690 308.665 ;
        RECT 14.635 305.975 189.690 307.165 ;
        RECT 159.920 304.475 189.690 305.975 ;
        RECT 14.635 302.525 189.690 304.475 ;
        RECT 159.920 301.025 189.690 302.525 ;
        RECT 14.635 299.835 189.690 301.025 ;
        RECT 159.920 298.335 189.690 299.835 ;
        RECT 14.635 296.385 189.690 298.335 ;
        RECT 159.920 294.885 189.690 296.385 ;
        RECT 14.635 293.695 189.690 294.885 ;
        RECT 159.920 292.195 189.690 293.695 ;
        RECT 14.635 290.245 189.690 292.195 ;
        RECT 159.920 288.745 189.690 290.245 ;
        RECT 14.635 287.555 189.690 288.745 ;
        RECT 159.920 286.055 189.690 287.555 ;
        RECT 14.635 284.105 189.690 286.055 ;
        RECT 159.920 282.605 189.690 284.105 ;
        RECT 14.635 281.415 189.690 282.605 ;
        RECT 159.920 279.915 189.690 281.415 ;
        RECT 14.635 277.965 189.690 279.915 ;
        RECT 159.920 276.465 189.690 277.965 ;
        RECT 14.635 275.275 189.690 276.465 ;
        RECT 159.920 273.775 189.690 275.275 ;
        RECT 14.635 271.825 189.690 273.775 ;
        RECT 159.920 270.325 189.690 271.825 ;
        RECT 14.635 269.135 189.690 270.325 ;
        RECT 159.920 267.635 189.690 269.135 ;
        RECT 14.635 265.685 189.690 267.635 ;
        RECT 159.920 264.185 189.690 265.685 ;
        RECT 14.635 262.995 189.690 264.185 ;
        RECT 159.920 261.495 189.690 262.995 ;
        RECT 14.635 259.545 189.690 261.495 ;
        RECT 159.920 258.045 189.690 259.545 ;
        RECT 14.635 256.855 189.690 258.045 ;
        RECT 159.920 255.355 189.690 256.855 ;
        RECT 14.635 253.405 189.690 255.355 ;
        RECT 159.920 251.905 189.690 253.405 ;
        RECT 14.635 250.715 189.690 251.905 ;
        RECT 159.920 249.215 189.690 250.715 ;
        RECT 14.635 247.265 189.690 249.215 ;
        RECT 159.920 245.765 189.690 247.265 ;
        RECT 14.635 244.575 189.690 245.765 ;
        RECT 159.920 243.075 189.690 244.575 ;
        RECT 14.635 241.125 189.690 243.075 ;
        RECT 159.920 239.625 189.690 241.125 ;
        RECT 14.635 238.435 189.690 239.625 ;
        RECT 159.920 236.935 189.690 238.435 ;
        RECT 14.635 234.985 189.690 236.935 ;
        RECT 159.920 233.485 189.690 234.985 ;
        RECT 14.635 232.295 189.690 233.485 ;
        RECT 159.920 230.795 189.690 232.295 ;
        RECT 14.635 228.845 189.690 230.795 ;
        RECT 159.920 227.345 189.690 228.845 ;
        RECT 14.635 226.155 189.690 227.345 ;
        RECT 159.920 224.655 189.690 226.155 ;
        RECT 14.635 222.705 189.690 224.655 ;
        RECT 159.920 221.205 189.690 222.705 ;
        RECT 14.635 220.015 189.690 221.205 ;
        RECT 159.920 218.515 189.690 220.015 ;
        RECT 14.635 216.565 189.690 218.515 ;
        RECT 159.920 215.065 189.690 216.565 ;
        RECT 14.635 213.875 189.690 215.065 ;
        RECT 159.920 212.375 189.690 213.875 ;
        RECT 14.635 210.425 189.690 212.375 ;
        RECT 159.920 208.925 189.690 210.425 ;
        RECT 14.635 207.735 189.690 208.925 ;
        RECT 159.920 206.235 189.690 207.735 ;
        RECT 14.635 204.285 189.690 206.235 ;
        RECT 159.920 202.785 189.690 204.285 ;
        RECT 14.635 201.595 189.690 202.785 ;
        RECT 159.920 200.095 189.690 201.595 ;
        RECT 14.635 198.145 189.690 200.095 ;
        RECT 159.920 196.645 189.690 198.145 ;
        RECT 14.635 195.455 189.690 196.645 ;
        RECT 159.920 193.955 189.690 195.455 ;
        RECT 14.635 192.005 189.690 193.955 ;
        RECT 159.920 190.505 189.690 192.005 ;
        RECT 14.635 189.315 189.690 190.505 ;
        RECT 159.920 187.815 189.690 189.315 ;
        RECT 14.635 185.865 189.690 187.815 ;
        RECT 159.920 184.365 189.690 185.865 ;
        RECT 14.635 183.175 189.690 184.365 ;
        RECT 159.920 181.675 189.690 183.175 ;
        RECT 14.635 179.725 189.690 181.675 ;
        RECT 159.920 178.225 189.690 179.725 ;
        RECT 14.635 177.035 189.690 178.225 ;
        RECT 159.920 175.535 189.690 177.035 ;
        RECT 14.635 173.585 189.690 175.535 ;
        RECT 159.920 172.085 189.690 173.585 ;
        RECT 14.635 170.895 189.690 172.085 ;
        RECT 159.920 169.395 189.690 170.895 ;
        RECT 14.635 167.445 189.690 169.395 ;
        RECT 159.920 165.945 189.690 167.445 ;
        RECT 14.635 164.755 189.690 165.945 ;
        RECT 159.920 163.255 189.690 164.755 ;
        RECT 14.635 161.305 189.690 163.255 ;
        RECT 159.920 159.805 189.690 161.305 ;
        RECT 14.635 158.615 189.690 159.805 ;
        RECT 159.920 157.115 189.690 158.615 ;
        RECT 14.635 155.165 189.690 157.115 ;
        RECT 159.920 153.665 189.690 155.165 ;
        RECT 14.635 152.475 189.690 153.665 ;
        RECT 159.920 150.975 189.690 152.475 ;
        RECT 14.635 149.025 189.690 150.975 ;
        RECT 159.920 147.525 189.690 149.025 ;
        RECT 14.635 146.335 189.690 147.525 ;
        RECT 159.920 144.835 189.690 146.335 ;
        RECT 14.635 142.885 189.690 144.835 ;
        RECT 159.920 141.385 189.690 142.885 ;
        RECT 14.635 140.195 189.690 141.385 ;
        RECT 159.920 138.695 189.690 140.195 ;
        RECT 14.635 136.745 189.690 138.695 ;
        RECT 159.920 135.245 189.690 136.745 ;
        RECT 14.635 134.055 189.690 135.245 ;
        RECT 159.920 132.555 189.690 134.055 ;
        RECT 14.635 130.605 189.690 132.555 ;
        RECT 159.920 129.105 189.690 130.605 ;
        RECT 14.635 127.915 189.690 129.105 ;
        RECT 159.920 126.415 189.690 127.915 ;
        RECT 14.635 124.465 189.690 126.415 ;
        RECT 159.920 122.965 189.690 124.465 ;
        RECT 14.635 121.775 189.690 122.965 ;
        RECT 159.920 120.275 189.690 121.775 ;
        RECT 14.635 118.325 189.690 120.275 ;
        RECT 159.920 116.825 189.690 118.325 ;
        RECT 14.635 115.635 189.690 116.825 ;
        RECT 159.920 114.135 189.690 115.635 ;
        RECT 14.635 112.185 189.690 114.135 ;
        RECT 159.920 110.685 189.690 112.185 ;
        RECT 14.635 109.495 189.690 110.685 ;
        RECT 159.920 107.995 189.690 109.495 ;
        RECT 14.635 106.045 189.690 107.995 ;
        RECT 159.920 104.545 189.690 106.045 ;
        RECT 14.635 103.355 189.690 104.545 ;
        RECT 159.920 101.855 189.690 103.355 ;
        RECT 14.635 99.905 189.690 101.855 ;
        RECT 159.920 98.405 189.690 99.905 ;
        RECT 14.635 97.215 189.690 98.405 ;
        RECT 159.920 95.715 189.690 97.215 ;
        RECT 14.635 93.765 189.690 95.715 ;
        RECT 159.920 92.265 189.690 93.765 ;
        RECT 14.635 91.075 189.690 92.265 ;
        RECT 159.920 89.575 189.690 91.075 ;
        RECT 14.635 87.625 189.690 89.575 ;
        RECT 159.920 86.125 189.690 87.625 ;
        RECT 14.635 84.935 189.690 86.125 ;
        RECT 159.920 83.435 189.690 84.935 ;
        RECT 14.635 81.485 189.690 83.435 ;
        RECT 159.920 79.985 189.690 81.485 ;
        RECT 14.635 78.795 189.690 79.985 ;
        RECT 159.920 77.295 189.690 78.795 ;
        RECT 14.635 75.345 189.690 77.295 ;
        RECT 159.920 73.845 189.690 75.345 ;
        RECT 14.635 72.655 189.690 73.845 ;
        RECT 159.920 71.155 189.690 72.655 ;
        RECT 14.635 69.205 189.690 71.155 ;
        RECT 159.920 67.705 189.690 69.205 ;
        RECT 14.635 66.515 189.690 67.705 ;
        RECT 159.920 65.015 189.690 66.515 ;
        RECT 14.635 63.065 189.690 65.015 ;
        RECT 159.920 61.565 189.690 63.065 ;
        RECT 14.635 60.375 189.690 61.565 ;
        RECT 159.920 58.875 189.690 60.375 ;
        RECT 14.635 56.925 189.690 58.875 ;
        RECT 159.920 55.425 189.690 56.925 ;
        RECT 14.635 54.235 189.690 55.425 ;
        RECT 159.920 52.735 189.690 54.235 ;
        RECT 14.635 50.785 189.690 52.735 ;
        RECT 159.920 49.285 189.690 50.785 ;
        RECT 14.635 48.095 189.690 49.285 ;
        RECT 159.920 46.595 189.690 48.095 ;
        RECT 14.635 44.645 189.690 46.595 ;
        RECT 159.920 43.145 189.690 44.645 ;
        RECT 14.635 41.955 189.690 43.145 ;
        RECT 159.920 40.455 189.690 41.955 ;
        RECT 14.635 38.505 189.690 40.455 ;
        RECT 159.920 37.005 189.690 38.505 ;
        RECT 14.635 35.815 189.690 37.005 ;
        RECT 159.920 34.315 189.690 35.815 ;
        RECT 14.635 32.365 189.690 34.315 ;
        RECT 159.920 30.865 189.690 32.365 ;
        RECT 14.635 29.675 189.690 30.865 ;
        RECT 159.920 28.175 189.690 29.675 ;
        RECT 14.635 26.225 189.690 28.175 ;
        RECT 159.920 24.725 189.690 26.225 ;
        RECT 14.635 23.535 189.690 24.725 ;
        RECT 159.920 22.035 189.690 23.535 ;
        RECT 14.635 20.085 189.690 22.035 ;
        RECT 159.920 18.585 189.690 20.085 ;
        RECT 14.635 17.395 189.690 18.585 ;
        RECT 159.920 15.895 189.690 17.395 ;
        RECT 14.635 13.945 189.690 15.895 ;
        RECT 159.920 12.445 189.690 13.945 ;
        RECT 14.635 11.255 189.690 12.445 ;
        RECT 159.920 9.755 189.690 11.255 ;
        RECT 14.635 7.805 189.690 9.755 ;
        RECT 159.920 7.740 189.690 7.805 ;
      LAYER met4 ;
        RECT 124.905 17.750 189.220 431.940 ;
  END
END top
END LIBRARY

