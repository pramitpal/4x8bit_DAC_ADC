magic
tech sky130A
magscale 1 2
timestamp 1688008296
<< nwell >>
rect 1280 4596 1946 4802
rect 3378 4784 4292 4792
rect 5622 4784 6250 4792
rect 3378 4596 4984 4784
rect 1280 4524 4984 4596
rect 1328 4272 4984 4524
rect 5622 4272 6942 4784
rect 1328 4264 3480 4272
rect 1328 4262 3408 4264
rect 2832 4258 3146 4262
rect 1280 3368 1946 3574
rect 3378 3556 4292 3564
rect 5622 3556 6250 3564
rect 3378 3368 4984 3556
rect 1280 3296 4984 3368
rect 1328 3044 4984 3296
rect 5622 3044 6942 3556
rect 1328 3036 3480 3044
rect 1328 3034 3408 3036
rect 2832 3030 3146 3034
rect 1280 2140 1946 2346
rect 3378 2328 4292 2336
rect 5622 2328 6250 2336
rect 3378 2140 4984 2328
rect 1280 2068 4984 2140
rect 1328 1816 4984 2068
rect 5622 1816 6942 2328
rect 1328 1808 3480 1816
rect 1328 1806 3408 1808
rect 2832 1802 3146 1806
rect 1280 912 1946 1118
rect 3378 1100 4292 1108
rect 3378 912 4984 1100
rect 1280 840 4984 912
rect 1328 588 4984 840
rect 1328 580 3480 588
rect 1328 578 3408 580
rect 2832 574 3146 578
<< pwell >>
rect 808 4650 1098 4656
rect 518 3978 1098 4650
rect 4364 4226 4940 4228
rect 6322 4226 6898 4228
rect 1372 4064 3350 4216
rect 3704 4076 4940 4226
rect 5662 4076 6898 4226
rect 3704 4074 4280 4076
rect 5662 4074 6238 4076
rect 3704 4070 4270 4074
rect 5662 4070 6228 4074
rect 1372 4058 1985 4064
rect 518 3972 800 3978
rect 1298 3878 1985 4058
rect 3678 3878 4270 4070
rect 5636 3878 6228 4070
rect 808 3422 1098 3428
rect 518 2750 1098 3422
rect 4364 2998 4940 3000
rect 6322 2998 6898 3000
rect 1372 2836 3350 2988
rect 3704 2848 4940 2998
rect 5662 2848 6898 2998
rect 3704 2846 4280 2848
rect 5662 2846 6238 2848
rect 3704 2842 4270 2846
rect 5662 2842 6228 2846
rect 1372 2830 1985 2836
rect 518 2744 800 2750
rect 1298 2650 1985 2830
rect 3678 2650 4270 2842
rect 5636 2650 6228 2842
rect 808 2194 1098 2200
rect 518 1522 1098 2194
rect 4364 1770 4940 1772
rect 6322 1770 6898 1772
rect 1372 1608 3350 1760
rect 3704 1620 4940 1770
rect 5662 1620 6898 1770
rect 3704 1618 4280 1620
rect 5662 1618 6238 1620
rect 3704 1614 4270 1618
rect 5662 1614 6228 1618
rect 1372 1602 1985 1608
rect 518 1516 800 1522
rect 1298 1422 1985 1602
rect 3678 1422 4270 1614
rect 5636 1422 6228 1614
rect 808 966 1098 972
rect 518 294 1098 966
rect 4364 542 4940 544
rect 1372 380 3350 532
rect 3704 392 4940 542
rect 3704 390 4280 392
rect 3704 386 4270 390
rect 1372 374 1985 380
rect 518 288 800 294
rect 1298 194 1985 374
rect 3678 194 4270 386
<< mvnmos >>
rect 1456 4090 1556 4190
rect 1744 4090 1844 4190
rect 2076 4090 2176 4190
rect 2418 4090 2518 4190
rect 2822 4090 2922 4190
rect 3166 4090 3266 4190
rect 3788 4100 3888 4200
rect 4096 4100 4196 4200
rect 4448 4102 4548 4202
rect 4756 4102 4856 4202
rect 5746 4100 5846 4200
rect 6054 4100 6154 4200
rect 6406 4102 6506 4202
rect 6714 4102 6814 4202
rect 1456 2862 1556 2962
rect 1744 2862 1844 2962
rect 2076 2862 2176 2962
rect 2418 2862 2518 2962
rect 2822 2862 2922 2962
rect 3166 2862 3266 2962
rect 3788 2872 3888 2972
rect 4096 2872 4196 2972
rect 4448 2874 4548 2974
rect 4756 2874 4856 2974
rect 5746 2872 5846 2972
rect 6054 2872 6154 2972
rect 6406 2874 6506 2974
rect 6714 2874 6814 2974
rect 1456 1634 1556 1734
rect 1744 1634 1844 1734
rect 2076 1634 2176 1734
rect 2418 1634 2518 1734
rect 2822 1634 2922 1734
rect 3166 1634 3266 1734
rect 3788 1644 3888 1744
rect 4096 1644 4196 1744
rect 4448 1646 4548 1746
rect 4756 1646 4856 1746
rect 5746 1644 5846 1744
rect 6054 1644 6154 1744
rect 6406 1646 6506 1746
rect 6714 1646 6814 1746
rect 1456 406 1556 506
rect 1744 406 1844 506
rect 2076 406 2176 506
rect 2418 406 2518 506
rect 2822 406 2922 506
rect 3166 406 3266 506
rect 3788 416 3888 516
rect 4096 416 4196 516
rect 4448 418 4548 518
rect 4756 418 4856 518
<< mvpmos >>
rect 1456 4328 1556 4528
rect 1744 4328 1844 4528
rect 2076 4328 2176 4528
rect 2418 4328 2518 4528
rect 2822 4328 2922 4528
rect 3166 4328 3266 4528
rect 3788 4338 3888 4538
rect 4096 4338 4196 4538
rect 4448 4338 4548 4538
rect 4756 4338 4856 4538
rect 5746 4338 5846 4538
rect 6054 4338 6154 4538
rect 6406 4338 6506 4538
rect 6714 4338 6814 4538
rect 1456 3100 1556 3300
rect 1744 3100 1844 3300
rect 2076 3100 2176 3300
rect 2418 3100 2518 3300
rect 2822 3100 2922 3300
rect 3166 3100 3266 3300
rect 3788 3110 3888 3310
rect 4096 3110 4196 3310
rect 4448 3110 4548 3310
rect 4756 3110 4856 3310
rect 5746 3110 5846 3310
rect 6054 3110 6154 3310
rect 6406 3110 6506 3310
rect 6714 3110 6814 3310
rect 1456 1872 1556 2072
rect 1744 1872 1844 2072
rect 2076 1872 2176 2072
rect 2418 1872 2518 2072
rect 2822 1872 2922 2072
rect 3166 1872 3266 2072
rect 3788 1882 3888 2082
rect 4096 1882 4196 2082
rect 4448 1882 4548 2082
rect 4756 1882 4856 2082
rect 5746 1882 5846 2082
rect 6054 1882 6154 2082
rect 6406 1882 6506 2082
rect 6714 1882 6814 2082
rect 1456 644 1556 844
rect 1744 644 1844 844
rect 2076 644 2176 844
rect 2418 644 2518 844
rect 2822 644 2922 844
rect 3166 644 3266 844
rect 3788 654 3888 854
rect 4096 654 4196 854
rect 4448 654 4548 854
rect 4756 654 4856 854
<< mvndiff >>
rect 544 4612 628 4624
rect 544 4578 569 4612
rect 603 4578 628 4612
rect 544 4521 628 4578
rect 544 4044 628 4101
rect 544 4010 569 4044
rect 603 4010 628 4044
rect 544 3998 628 4010
rect 690 4612 774 4624
rect 690 4578 715 4612
rect 749 4578 774 4612
rect 690 4521 774 4578
rect 690 4044 774 4101
rect 690 4010 715 4044
rect 749 4010 774 4044
rect 690 3998 774 4010
rect 834 4618 918 4630
rect 834 4584 859 4618
rect 893 4584 918 4618
rect 834 4527 918 4584
rect 834 4050 918 4107
rect 834 4016 859 4050
rect 893 4016 918 4050
rect 834 4004 918 4016
rect 988 4618 1072 4630
rect 988 4584 1013 4618
rect 1047 4584 1072 4618
rect 988 4527 1072 4584
rect 988 4050 1072 4107
rect 1398 4157 1456 4190
rect 1398 4123 1410 4157
rect 1444 4123 1456 4157
rect 1398 4090 1456 4123
rect 1556 4157 1614 4190
rect 1556 4123 1568 4157
rect 1602 4123 1614 4157
rect 1556 4090 1614 4123
rect 1686 4157 1744 4190
rect 1686 4123 1698 4157
rect 1732 4123 1744 4157
rect 1686 4090 1744 4123
rect 1844 4157 1902 4190
rect 1844 4123 1856 4157
rect 1890 4123 1902 4157
rect 1844 4090 1902 4123
rect 2018 4157 2076 4190
rect 2018 4123 2030 4157
rect 2064 4123 2076 4157
rect 2018 4090 2076 4123
rect 2176 4157 2234 4190
rect 2176 4123 2188 4157
rect 2222 4123 2234 4157
rect 2176 4090 2234 4123
rect 2360 4157 2418 4190
rect 2360 4123 2372 4157
rect 2406 4123 2418 4157
rect 2360 4090 2418 4123
rect 2518 4157 2576 4190
rect 2518 4123 2530 4157
rect 2564 4123 2576 4157
rect 2518 4090 2576 4123
rect 2764 4157 2822 4190
rect 2764 4123 2776 4157
rect 2810 4123 2822 4157
rect 2764 4090 2822 4123
rect 2922 4157 2980 4190
rect 2922 4123 2934 4157
rect 2968 4123 2980 4157
rect 2922 4090 2980 4123
rect 3108 4157 3166 4190
rect 3108 4123 3120 4157
rect 3154 4123 3166 4157
rect 3108 4090 3166 4123
rect 3266 4157 3324 4190
rect 3266 4123 3278 4157
rect 3312 4123 3324 4157
rect 3266 4090 3324 4123
rect 3730 4167 3788 4200
rect 3730 4133 3742 4167
rect 3776 4133 3788 4167
rect 3730 4100 3788 4133
rect 3888 4167 3946 4200
rect 3888 4133 3900 4167
rect 3934 4133 3946 4167
rect 3888 4100 3946 4133
rect 4038 4167 4096 4200
rect 4038 4133 4050 4167
rect 4084 4133 4096 4167
rect 4038 4100 4096 4133
rect 4196 4167 4254 4200
rect 4196 4133 4208 4167
rect 4242 4133 4254 4167
rect 4196 4100 4254 4133
rect 4390 4169 4448 4202
rect 4390 4135 4402 4169
rect 4436 4135 4448 4169
rect 4390 4102 4448 4135
rect 4548 4169 4606 4202
rect 4548 4135 4560 4169
rect 4594 4135 4606 4169
rect 4548 4102 4606 4135
rect 4698 4169 4756 4202
rect 4698 4135 4710 4169
rect 4744 4135 4756 4169
rect 4698 4102 4756 4135
rect 4856 4169 4914 4202
rect 4856 4135 4868 4169
rect 4902 4135 4914 4169
rect 4856 4102 4914 4135
rect 5688 4168 5746 4200
rect 5688 4134 5700 4168
rect 5734 4134 5746 4168
rect 5688 4100 5746 4134
rect 5846 4168 5904 4200
rect 5846 4134 5858 4168
rect 5892 4134 5904 4168
rect 5846 4100 5904 4134
rect 5996 4168 6054 4200
rect 5996 4134 6008 4168
rect 6042 4134 6054 4168
rect 5996 4100 6054 4134
rect 6154 4168 6212 4200
rect 6154 4134 6166 4168
rect 6200 4134 6212 4168
rect 6154 4100 6212 4134
rect 6348 4170 6406 4202
rect 6348 4136 6360 4170
rect 6394 4136 6406 4170
rect 6348 4102 6406 4136
rect 6506 4170 6564 4202
rect 6506 4136 6518 4170
rect 6552 4136 6564 4170
rect 6506 4102 6564 4136
rect 6656 4170 6714 4202
rect 6656 4136 6668 4170
rect 6702 4136 6714 4170
rect 6656 4102 6714 4136
rect 6814 4170 6872 4202
rect 6814 4136 6826 4170
rect 6860 4136 6872 4170
rect 6814 4102 6872 4136
rect 988 4016 1013 4050
rect 1047 4016 1072 4050
rect 988 4004 1072 4016
rect 544 3384 628 3396
rect 544 3350 569 3384
rect 603 3350 628 3384
rect 544 3293 628 3350
rect 544 2816 628 2873
rect 544 2782 569 2816
rect 603 2782 628 2816
rect 544 2770 628 2782
rect 690 3384 774 3396
rect 690 3350 715 3384
rect 749 3350 774 3384
rect 690 3293 774 3350
rect 690 2816 774 2873
rect 690 2782 715 2816
rect 749 2782 774 2816
rect 690 2770 774 2782
rect 834 3390 918 3402
rect 834 3356 859 3390
rect 893 3356 918 3390
rect 834 3299 918 3356
rect 834 2822 918 2879
rect 834 2788 859 2822
rect 893 2788 918 2822
rect 834 2776 918 2788
rect 988 3390 1072 3402
rect 988 3356 1013 3390
rect 1047 3356 1072 3390
rect 988 3299 1072 3356
rect 988 2822 1072 2879
rect 1398 2929 1456 2962
rect 1398 2895 1410 2929
rect 1444 2895 1456 2929
rect 1398 2862 1456 2895
rect 1556 2929 1614 2962
rect 1556 2895 1568 2929
rect 1602 2895 1614 2929
rect 1556 2862 1614 2895
rect 1686 2929 1744 2962
rect 1686 2895 1698 2929
rect 1732 2895 1744 2929
rect 1686 2862 1744 2895
rect 1844 2929 1902 2962
rect 1844 2895 1856 2929
rect 1890 2895 1902 2929
rect 1844 2862 1902 2895
rect 2018 2929 2076 2962
rect 2018 2895 2030 2929
rect 2064 2895 2076 2929
rect 2018 2862 2076 2895
rect 2176 2929 2234 2962
rect 2176 2895 2188 2929
rect 2222 2895 2234 2929
rect 2176 2862 2234 2895
rect 2360 2929 2418 2962
rect 2360 2895 2372 2929
rect 2406 2895 2418 2929
rect 2360 2862 2418 2895
rect 2518 2929 2576 2962
rect 2518 2895 2530 2929
rect 2564 2895 2576 2929
rect 2518 2862 2576 2895
rect 2764 2929 2822 2962
rect 2764 2895 2776 2929
rect 2810 2895 2822 2929
rect 2764 2862 2822 2895
rect 2922 2929 2980 2962
rect 2922 2895 2934 2929
rect 2968 2895 2980 2929
rect 2922 2862 2980 2895
rect 3108 2929 3166 2962
rect 3108 2895 3120 2929
rect 3154 2895 3166 2929
rect 3108 2862 3166 2895
rect 3266 2929 3324 2962
rect 3266 2895 3278 2929
rect 3312 2895 3324 2929
rect 3266 2862 3324 2895
rect 3730 2939 3788 2972
rect 3730 2905 3742 2939
rect 3776 2905 3788 2939
rect 3730 2872 3788 2905
rect 3888 2939 3946 2972
rect 3888 2905 3900 2939
rect 3934 2905 3946 2939
rect 3888 2872 3946 2905
rect 4038 2939 4096 2972
rect 4038 2905 4050 2939
rect 4084 2905 4096 2939
rect 4038 2872 4096 2905
rect 4196 2939 4254 2972
rect 4196 2905 4208 2939
rect 4242 2905 4254 2939
rect 4196 2872 4254 2905
rect 4390 2941 4448 2974
rect 4390 2907 4402 2941
rect 4436 2907 4448 2941
rect 4390 2874 4448 2907
rect 4548 2941 4606 2974
rect 4548 2907 4560 2941
rect 4594 2907 4606 2941
rect 4548 2874 4606 2907
rect 4698 2941 4756 2974
rect 4698 2907 4710 2941
rect 4744 2907 4756 2941
rect 4698 2874 4756 2907
rect 4856 2941 4914 2974
rect 4856 2907 4868 2941
rect 4902 2907 4914 2941
rect 4856 2874 4914 2907
rect 5688 2940 5746 2972
rect 5688 2906 5700 2940
rect 5734 2906 5746 2940
rect 5688 2872 5746 2906
rect 5846 2940 5904 2972
rect 5846 2906 5858 2940
rect 5892 2906 5904 2940
rect 5846 2872 5904 2906
rect 5996 2940 6054 2972
rect 5996 2906 6008 2940
rect 6042 2906 6054 2940
rect 5996 2872 6054 2906
rect 6154 2940 6212 2972
rect 6154 2906 6166 2940
rect 6200 2906 6212 2940
rect 6154 2872 6212 2906
rect 6348 2942 6406 2974
rect 6348 2908 6360 2942
rect 6394 2908 6406 2942
rect 6348 2874 6406 2908
rect 6506 2942 6564 2974
rect 6506 2908 6518 2942
rect 6552 2908 6564 2942
rect 6506 2874 6564 2908
rect 6656 2942 6714 2974
rect 6656 2908 6668 2942
rect 6702 2908 6714 2942
rect 6656 2874 6714 2908
rect 6814 2942 6872 2974
rect 6814 2908 6826 2942
rect 6860 2908 6872 2942
rect 6814 2874 6872 2908
rect 988 2788 1013 2822
rect 1047 2788 1072 2822
rect 988 2776 1072 2788
rect 544 2156 628 2168
rect 544 2122 569 2156
rect 603 2122 628 2156
rect 544 2065 628 2122
rect 544 1588 628 1645
rect 544 1554 569 1588
rect 603 1554 628 1588
rect 544 1542 628 1554
rect 690 2156 774 2168
rect 690 2122 715 2156
rect 749 2122 774 2156
rect 690 2065 774 2122
rect 690 1588 774 1645
rect 690 1554 715 1588
rect 749 1554 774 1588
rect 690 1542 774 1554
rect 834 2162 918 2174
rect 834 2128 859 2162
rect 893 2128 918 2162
rect 834 2071 918 2128
rect 834 1594 918 1651
rect 834 1560 859 1594
rect 893 1560 918 1594
rect 834 1548 918 1560
rect 988 2162 1072 2174
rect 988 2128 1013 2162
rect 1047 2128 1072 2162
rect 988 2071 1072 2128
rect 988 1594 1072 1651
rect 1398 1701 1456 1734
rect 1398 1667 1410 1701
rect 1444 1667 1456 1701
rect 1398 1634 1456 1667
rect 1556 1701 1614 1734
rect 1556 1667 1568 1701
rect 1602 1667 1614 1701
rect 1556 1634 1614 1667
rect 1686 1701 1744 1734
rect 1686 1667 1698 1701
rect 1732 1667 1744 1701
rect 1686 1634 1744 1667
rect 1844 1701 1902 1734
rect 1844 1667 1856 1701
rect 1890 1667 1902 1701
rect 1844 1634 1902 1667
rect 2018 1701 2076 1734
rect 2018 1667 2030 1701
rect 2064 1667 2076 1701
rect 2018 1634 2076 1667
rect 2176 1701 2234 1734
rect 2176 1667 2188 1701
rect 2222 1667 2234 1701
rect 2176 1634 2234 1667
rect 2360 1701 2418 1734
rect 2360 1667 2372 1701
rect 2406 1667 2418 1701
rect 2360 1634 2418 1667
rect 2518 1701 2576 1734
rect 2518 1667 2530 1701
rect 2564 1667 2576 1701
rect 2518 1634 2576 1667
rect 2764 1701 2822 1734
rect 2764 1667 2776 1701
rect 2810 1667 2822 1701
rect 2764 1634 2822 1667
rect 2922 1701 2980 1734
rect 2922 1667 2934 1701
rect 2968 1667 2980 1701
rect 2922 1634 2980 1667
rect 3108 1701 3166 1734
rect 3108 1667 3120 1701
rect 3154 1667 3166 1701
rect 3108 1634 3166 1667
rect 3266 1701 3324 1734
rect 3266 1667 3278 1701
rect 3312 1667 3324 1701
rect 3266 1634 3324 1667
rect 3730 1711 3788 1744
rect 3730 1677 3742 1711
rect 3776 1677 3788 1711
rect 3730 1644 3788 1677
rect 3888 1711 3946 1744
rect 3888 1677 3900 1711
rect 3934 1677 3946 1711
rect 3888 1644 3946 1677
rect 4038 1711 4096 1744
rect 4038 1677 4050 1711
rect 4084 1677 4096 1711
rect 4038 1644 4096 1677
rect 4196 1711 4254 1744
rect 4196 1677 4208 1711
rect 4242 1677 4254 1711
rect 4196 1644 4254 1677
rect 4390 1713 4448 1746
rect 4390 1679 4402 1713
rect 4436 1679 4448 1713
rect 4390 1646 4448 1679
rect 4548 1713 4606 1746
rect 4548 1679 4560 1713
rect 4594 1679 4606 1713
rect 4548 1646 4606 1679
rect 4698 1713 4756 1746
rect 4698 1679 4710 1713
rect 4744 1679 4756 1713
rect 4698 1646 4756 1679
rect 4856 1713 4914 1746
rect 4856 1679 4868 1713
rect 4902 1679 4914 1713
rect 4856 1646 4914 1679
rect 5688 1712 5746 1744
rect 5688 1678 5700 1712
rect 5734 1678 5746 1712
rect 5688 1644 5746 1678
rect 5846 1712 5904 1744
rect 5846 1678 5858 1712
rect 5892 1678 5904 1712
rect 5846 1644 5904 1678
rect 5996 1712 6054 1744
rect 5996 1678 6008 1712
rect 6042 1678 6054 1712
rect 5996 1644 6054 1678
rect 6154 1712 6212 1744
rect 6154 1678 6166 1712
rect 6200 1678 6212 1712
rect 6154 1644 6212 1678
rect 6348 1714 6406 1746
rect 6348 1680 6360 1714
rect 6394 1680 6406 1714
rect 6348 1646 6406 1680
rect 6506 1714 6564 1746
rect 6506 1680 6518 1714
rect 6552 1680 6564 1714
rect 6506 1646 6564 1680
rect 6656 1714 6714 1746
rect 6656 1680 6668 1714
rect 6702 1680 6714 1714
rect 6656 1646 6714 1680
rect 6814 1714 6872 1746
rect 6814 1680 6826 1714
rect 6860 1680 6872 1714
rect 6814 1646 6872 1680
rect 988 1560 1013 1594
rect 1047 1560 1072 1594
rect 988 1548 1072 1560
rect 544 928 628 940
rect 544 894 569 928
rect 603 894 628 928
rect 544 837 628 894
rect 544 360 628 417
rect 544 326 569 360
rect 603 326 628 360
rect 544 314 628 326
rect 690 928 774 940
rect 690 894 715 928
rect 749 894 774 928
rect 690 837 774 894
rect 690 360 774 417
rect 690 326 715 360
rect 749 326 774 360
rect 690 314 774 326
rect 834 934 918 946
rect 834 900 859 934
rect 893 900 918 934
rect 834 843 918 900
rect 834 366 918 423
rect 834 332 859 366
rect 893 332 918 366
rect 834 320 918 332
rect 988 934 1072 946
rect 988 900 1013 934
rect 1047 900 1072 934
rect 988 843 1072 900
rect 988 366 1072 423
rect 1398 473 1456 506
rect 1398 439 1410 473
rect 1444 439 1456 473
rect 1398 406 1456 439
rect 1556 473 1614 506
rect 1556 439 1568 473
rect 1602 439 1614 473
rect 1556 406 1614 439
rect 1686 473 1744 506
rect 1686 439 1698 473
rect 1732 439 1744 473
rect 1686 406 1744 439
rect 1844 473 1902 506
rect 1844 439 1856 473
rect 1890 439 1902 473
rect 1844 406 1902 439
rect 2018 473 2076 506
rect 2018 439 2030 473
rect 2064 439 2076 473
rect 2018 406 2076 439
rect 2176 473 2234 506
rect 2176 439 2188 473
rect 2222 439 2234 473
rect 2176 406 2234 439
rect 2360 473 2418 506
rect 2360 439 2372 473
rect 2406 439 2418 473
rect 2360 406 2418 439
rect 2518 473 2576 506
rect 2518 439 2530 473
rect 2564 439 2576 473
rect 2518 406 2576 439
rect 2764 473 2822 506
rect 2764 439 2776 473
rect 2810 439 2822 473
rect 2764 406 2822 439
rect 2922 473 2980 506
rect 2922 439 2934 473
rect 2968 439 2980 473
rect 2922 406 2980 439
rect 3108 473 3166 506
rect 3108 439 3120 473
rect 3154 439 3166 473
rect 3108 406 3166 439
rect 3266 473 3324 506
rect 3266 439 3278 473
rect 3312 439 3324 473
rect 3266 406 3324 439
rect 3730 483 3788 516
rect 3730 449 3742 483
rect 3776 449 3788 483
rect 3730 416 3788 449
rect 3888 483 3946 516
rect 3888 449 3900 483
rect 3934 449 3946 483
rect 3888 416 3946 449
rect 4038 483 4096 516
rect 4038 449 4050 483
rect 4084 449 4096 483
rect 4038 416 4096 449
rect 4196 483 4254 516
rect 4196 449 4208 483
rect 4242 449 4254 483
rect 4196 416 4254 449
rect 4390 485 4448 518
rect 4390 451 4402 485
rect 4436 451 4448 485
rect 4390 418 4448 451
rect 4548 485 4606 518
rect 4548 451 4560 485
rect 4594 451 4606 485
rect 4548 418 4606 451
rect 4698 485 4756 518
rect 4698 451 4710 485
rect 4744 451 4756 485
rect 4698 418 4756 451
rect 4856 485 4914 518
rect 4856 451 4868 485
rect 4902 451 4914 485
rect 4856 418 4914 451
rect 988 332 1013 366
rect 1047 332 1072 366
rect 988 320 1072 332
<< mvpdiff >>
rect 1398 4513 1456 4528
rect 1398 4479 1410 4513
rect 1444 4479 1456 4513
rect 1398 4445 1456 4479
rect 1398 4411 1410 4445
rect 1444 4411 1456 4445
rect 1398 4377 1456 4411
rect 1398 4343 1410 4377
rect 1444 4343 1456 4377
rect 1398 4328 1456 4343
rect 1556 4513 1614 4528
rect 1556 4479 1568 4513
rect 1602 4479 1614 4513
rect 1556 4445 1614 4479
rect 1556 4411 1568 4445
rect 1602 4411 1614 4445
rect 1556 4377 1614 4411
rect 1556 4343 1568 4377
rect 1602 4343 1614 4377
rect 1556 4328 1614 4343
rect 1686 4513 1744 4528
rect 1686 4479 1698 4513
rect 1732 4479 1744 4513
rect 1686 4445 1744 4479
rect 1686 4411 1698 4445
rect 1732 4411 1744 4445
rect 1686 4377 1744 4411
rect 1686 4343 1698 4377
rect 1732 4343 1744 4377
rect 1686 4328 1744 4343
rect 1844 4513 1902 4528
rect 1844 4479 1856 4513
rect 1890 4479 1902 4513
rect 1844 4445 1902 4479
rect 1844 4411 1856 4445
rect 1890 4411 1902 4445
rect 1844 4377 1902 4411
rect 1844 4343 1856 4377
rect 1890 4343 1902 4377
rect 1844 4328 1902 4343
rect 2018 4513 2076 4528
rect 2018 4479 2030 4513
rect 2064 4479 2076 4513
rect 2018 4445 2076 4479
rect 2018 4411 2030 4445
rect 2064 4411 2076 4445
rect 2018 4377 2076 4411
rect 2018 4343 2030 4377
rect 2064 4343 2076 4377
rect 2018 4328 2076 4343
rect 2176 4513 2234 4528
rect 2176 4479 2188 4513
rect 2222 4479 2234 4513
rect 2176 4445 2234 4479
rect 2176 4411 2188 4445
rect 2222 4411 2234 4445
rect 2176 4377 2234 4411
rect 2176 4343 2188 4377
rect 2222 4343 2234 4377
rect 2176 4328 2234 4343
rect 2360 4513 2418 4528
rect 2360 4479 2372 4513
rect 2406 4479 2418 4513
rect 2360 4445 2418 4479
rect 2360 4411 2372 4445
rect 2406 4411 2418 4445
rect 2360 4377 2418 4411
rect 2360 4343 2372 4377
rect 2406 4343 2418 4377
rect 2360 4328 2418 4343
rect 2518 4513 2576 4528
rect 2518 4479 2530 4513
rect 2564 4479 2576 4513
rect 2518 4445 2576 4479
rect 2518 4411 2530 4445
rect 2564 4411 2576 4445
rect 2518 4377 2576 4411
rect 2518 4343 2530 4377
rect 2564 4343 2576 4377
rect 2518 4328 2576 4343
rect 2764 4513 2822 4528
rect 2764 4479 2776 4513
rect 2810 4479 2822 4513
rect 2764 4445 2822 4479
rect 2764 4411 2776 4445
rect 2810 4411 2822 4445
rect 2764 4377 2822 4411
rect 2764 4343 2776 4377
rect 2810 4343 2822 4377
rect 2764 4328 2822 4343
rect 2922 4513 2980 4528
rect 2922 4479 2934 4513
rect 2968 4479 2980 4513
rect 2922 4445 2980 4479
rect 2922 4411 2934 4445
rect 2968 4411 2980 4445
rect 2922 4377 2980 4411
rect 2922 4343 2934 4377
rect 2968 4343 2980 4377
rect 2922 4328 2980 4343
rect 3108 4513 3166 4528
rect 3108 4479 3120 4513
rect 3154 4479 3166 4513
rect 3108 4445 3166 4479
rect 3108 4411 3120 4445
rect 3154 4411 3166 4445
rect 3108 4377 3166 4411
rect 3108 4343 3120 4377
rect 3154 4343 3166 4377
rect 3108 4328 3166 4343
rect 3266 4513 3324 4528
rect 3266 4479 3278 4513
rect 3312 4479 3324 4513
rect 3266 4445 3324 4479
rect 3266 4411 3278 4445
rect 3312 4411 3324 4445
rect 3266 4377 3324 4411
rect 3266 4343 3278 4377
rect 3312 4343 3324 4377
rect 3266 4328 3324 4343
rect 3730 4523 3788 4538
rect 3730 4489 3742 4523
rect 3776 4489 3788 4523
rect 3730 4455 3788 4489
rect 3730 4421 3742 4455
rect 3776 4421 3788 4455
rect 3730 4387 3788 4421
rect 3730 4353 3742 4387
rect 3776 4353 3788 4387
rect 3730 4338 3788 4353
rect 3888 4523 3946 4538
rect 3888 4489 3900 4523
rect 3934 4489 3946 4523
rect 3888 4455 3946 4489
rect 3888 4421 3900 4455
rect 3934 4421 3946 4455
rect 3888 4387 3946 4421
rect 3888 4353 3900 4387
rect 3934 4353 3946 4387
rect 3888 4338 3946 4353
rect 4038 4523 4096 4538
rect 4038 4489 4050 4523
rect 4084 4489 4096 4523
rect 4038 4455 4096 4489
rect 4038 4421 4050 4455
rect 4084 4421 4096 4455
rect 4038 4387 4096 4421
rect 4038 4353 4050 4387
rect 4084 4353 4096 4387
rect 4038 4338 4096 4353
rect 4196 4523 4254 4538
rect 4196 4489 4208 4523
rect 4242 4489 4254 4523
rect 4196 4455 4254 4489
rect 4196 4421 4208 4455
rect 4242 4421 4254 4455
rect 4196 4387 4254 4421
rect 4196 4353 4208 4387
rect 4242 4353 4254 4387
rect 4196 4338 4254 4353
rect 4390 4523 4448 4538
rect 4390 4489 4402 4523
rect 4436 4489 4448 4523
rect 4390 4455 4448 4489
rect 4390 4421 4402 4455
rect 4436 4421 4448 4455
rect 4390 4387 4448 4421
rect 4390 4353 4402 4387
rect 4436 4353 4448 4387
rect 4390 4338 4448 4353
rect 4548 4523 4606 4538
rect 4548 4489 4560 4523
rect 4594 4489 4606 4523
rect 4548 4455 4606 4489
rect 4548 4421 4560 4455
rect 4594 4421 4606 4455
rect 4548 4387 4606 4421
rect 4548 4353 4560 4387
rect 4594 4353 4606 4387
rect 4548 4338 4606 4353
rect 4698 4523 4756 4538
rect 4698 4489 4710 4523
rect 4744 4489 4756 4523
rect 4698 4455 4756 4489
rect 4698 4421 4710 4455
rect 4744 4421 4756 4455
rect 4698 4387 4756 4421
rect 4698 4353 4710 4387
rect 4744 4353 4756 4387
rect 4698 4338 4756 4353
rect 4856 4523 4914 4538
rect 4856 4489 4868 4523
rect 4902 4489 4914 4523
rect 4856 4455 4914 4489
rect 4856 4421 4868 4455
rect 4902 4421 4914 4455
rect 4856 4387 4914 4421
rect 4856 4353 4868 4387
rect 4902 4353 4914 4387
rect 4856 4338 4914 4353
rect 5688 4524 5746 4538
rect 5688 4490 5700 4524
rect 5734 4490 5746 4524
rect 5688 4456 5746 4490
rect 5688 4422 5700 4456
rect 5734 4422 5746 4456
rect 5688 4388 5746 4422
rect 5688 4354 5700 4388
rect 5734 4354 5746 4388
rect 5688 4338 5746 4354
rect 5846 4524 5904 4538
rect 5846 4490 5858 4524
rect 5892 4490 5904 4524
rect 5846 4456 5904 4490
rect 5846 4422 5858 4456
rect 5892 4422 5904 4456
rect 5846 4388 5904 4422
rect 5846 4354 5858 4388
rect 5892 4354 5904 4388
rect 5846 4338 5904 4354
rect 5996 4524 6054 4538
rect 5996 4490 6008 4524
rect 6042 4490 6054 4524
rect 5996 4456 6054 4490
rect 5996 4422 6008 4456
rect 6042 4422 6054 4456
rect 5996 4388 6054 4422
rect 5996 4354 6008 4388
rect 6042 4354 6054 4388
rect 5996 4338 6054 4354
rect 6154 4524 6212 4538
rect 6154 4490 6166 4524
rect 6200 4490 6212 4524
rect 6154 4456 6212 4490
rect 6154 4422 6166 4456
rect 6200 4422 6212 4456
rect 6154 4388 6212 4422
rect 6154 4354 6166 4388
rect 6200 4354 6212 4388
rect 6154 4338 6212 4354
rect 6348 4524 6406 4538
rect 6348 4490 6360 4524
rect 6394 4490 6406 4524
rect 6348 4456 6406 4490
rect 6348 4422 6360 4456
rect 6394 4422 6406 4456
rect 6348 4388 6406 4422
rect 6348 4354 6360 4388
rect 6394 4354 6406 4388
rect 6348 4338 6406 4354
rect 6506 4524 6564 4538
rect 6506 4490 6518 4524
rect 6552 4490 6564 4524
rect 6506 4456 6564 4490
rect 6506 4422 6518 4456
rect 6552 4422 6564 4456
rect 6506 4388 6564 4422
rect 6506 4354 6518 4388
rect 6552 4354 6564 4388
rect 6506 4338 6564 4354
rect 6656 4524 6714 4538
rect 6656 4490 6668 4524
rect 6702 4490 6714 4524
rect 6656 4456 6714 4490
rect 6656 4422 6668 4456
rect 6702 4422 6714 4456
rect 6656 4388 6714 4422
rect 6656 4354 6668 4388
rect 6702 4354 6714 4388
rect 6656 4338 6714 4354
rect 6814 4524 6872 4538
rect 6814 4490 6826 4524
rect 6860 4490 6872 4524
rect 6814 4456 6872 4490
rect 6814 4422 6826 4456
rect 6860 4422 6872 4456
rect 6814 4388 6872 4422
rect 6814 4354 6826 4388
rect 6860 4354 6872 4388
rect 6814 4338 6872 4354
rect 1398 3285 1456 3300
rect 1398 3251 1410 3285
rect 1444 3251 1456 3285
rect 1398 3217 1456 3251
rect 1398 3183 1410 3217
rect 1444 3183 1456 3217
rect 1398 3149 1456 3183
rect 1398 3115 1410 3149
rect 1444 3115 1456 3149
rect 1398 3100 1456 3115
rect 1556 3285 1614 3300
rect 1556 3251 1568 3285
rect 1602 3251 1614 3285
rect 1556 3217 1614 3251
rect 1556 3183 1568 3217
rect 1602 3183 1614 3217
rect 1556 3149 1614 3183
rect 1556 3115 1568 3149
rect 1602 3115 1614 3149
rect 1556 3100 1614 3115
rect 1686 3285 1744 3300
rect 1686 3251 1698 3285
rect 1732 3251 1744 3285
rect 1686 3217 1744 3251
rect 1686 3183 1698 3217
rect 1732 3183 1744 3217
rect 1686 3149 1744 3183
rect 1686 3115 1698 3149
rect 1732 3115 1744 3149
rect 1686 3100 1744 3115
rect 1844 3285 1902 3300
rect 1844 3251 1856 3285
rect 1890 3251 1902 3285
rect 1844 3217 1902 3251
rect 1844 3183 1856 3217
rect 1890 3183 1902 3217
rect 1844 3149 1902 3183
rect 1844 3115 1856 3149
rect 1890 3115 1902 3149
rect 1844 3100 1902 3115
rect 2018 3285 2076 3300
rect 2018 3251 2030 3285
rect 2064 3251 2076 3285
rect 2018 3217 2076 3251
rect 2018 3183 2030 3217
rect 2064 3183 2076 3217
rect 2018 3149 2076 3183
rect 2018 3115 2030 3149
rect 2064 3115 2076 3149
rect 2018 3100 2076 3115
rect 2176 3285 2234 3300
rect 2176 3251 2188 3285
rect 2222 3251 2234 3285
rect 2176 3217 2234 3251
rect 2176 3183 2188 3217
rect 2222 3183 2234 3217
rect 2176 3149 2234 3183
rect 2176 3115 2188 3149
rect 2222 3115 2234 3149
rect 2176 3100 2234 3115
rect 2360 3285 2418 3300
rect 2360 3251 2372 3285
rect 2406 3251 2418 3285
rect 2360 3217 2418 3251
rect 2360 3183 2372 3217
rect 2406 3183 2418 3217
rect 2360 3149 2418 3183
rect 2360 3115 2372 3149
rect 2406 3115 2418 3149
rect 2360 3100 2418 3115
rect 2518 3285 2576 3300
rect 2518 3251 2530 3285
rect 2564 3251 2576 3285
rect 2518 3217 2576 3251
rect 2518 3183 2530 3217
rect 2564 3183 2576 3217
rect 2518 3149 2576 3183
rect 2518 3115 2530 3149
rect 2564 3115 2576 3149
rect 2518 3100 2576 3115
rect 2764 3285 2822 3300
rect 2764 3251 2776 3285
rect 2810 3251 2822 3285
rect 2764 3217 2822 3251
rect 2764 3183 2776 3217
rect 2810 3183 2822 3217
rect 2764 3149 2822 3183
rect 2764 3115 2776 3149
rect 2810 3115 2822 3149
rect 2764 3100 2822 3115
rect 2922 3285 2980 3300
rect 2922 3251 2934 3285
rect 2968 3251 2980 3285
rect 2922 3217 2980 3251
rect 2922 3183 2934 3217
rect 2968 3183 2980 3217
rect 2922 3149 2980 3183
rect 2922 3115 2934 3149
rect 2968 3115 2980 3149
rect 2922 3100 2980 3115
rect 3108 3285 3166 3300
rect 3108 3251 3120 3285
rect 3154 3251 3166 3285
rect 3108 3217 3166 3251
rect 3108 3183 3120 3217
rect 3154 3183 3166 3217
rect 3108 3149 3166 3183
rect 3108 3115 3120 3149
rect 3154 3115 3166 3149
rect 3108 3100 3166 3115
rect 3266 3285 3324 3300
rect 3266 3251 3278 3285
rect 3312 3251 3324 3285
rect 3266 3217 3324 3251
rect 3266 3183 3278 3217
rect 3312 3183 3324 3217
rect 3266 3149 3324 3183
rect 3266 3115 3278 3149
rect 3312 3115 3324 3149
rect 3266 3100 3324 3115
rect 3730 3295 3788 3310
rect 3730 3261 3742 3295
rect 3776 3261 3788 3295
rect 3730 3227 3788 3261
rect 3730 3193 3742 3227
rect 3776 3193 3788 3227
rect 3730 3159 3788 3193
rect 3730 3125 3742 3159
rect 3776 3125 3788 3159
rect 3730 3110 3788 3125
rect 3888 3295 3946 3310
rect 3888 3261 3900 3295
rect 3934 3261 3946 3295
rect 3888 3227 3946 3261
rect 3888 3193 3900 3227
rect 3934 3193 3946 3227
rect 3888 3159 3946 3193
rect 3888 3125 3900 3159
rect 3934 3125 3946 3159
rect 3888 3110 3946 3125
rect 4038 3295 4096 3310
rect 4038 3261 4050 3295
rect 4084 3261 4096 3295
rect 4038 3227 4096 3261
rect 4038 3193 4050 3227
rect 4084 3193 4096 3227
rect 4038 3159 4096 3193
rect 4038 3125 4050 3159
rect 4084 3125 4096 3159
rect 4038 3110 4096 3125
rect 4196 3295 4254 3310
rect 4196 3261 4208 3295
rect 4242 3261 4254 3295
rect 4196 3227 4254 3261
rect 4196 3193 4208 3227
rect 4242 3193 4254 3227
rect 4196 3159 4254 3193
rect 4196 3125 4208 3159
rect 4242 3125 4254 3159
rect 4196 3110 4254 3125
rect 4390 3295 4448 3310
rect 4390 3261 4402 3295
rect 4436 3261 4448 3295
rect 4390 3227 4448 3261
rect 4390 3193 4402 3227
rect 4436 3193 4448 3227
rect 4390 3159 4448 3193
rect 4390 3125 4402 3159
rect 4436 3125 4448 3159
rect 4390 3110 4448 3125
rect 4548 3295 4606 3310
rect 4548 3261 4560 3295
rect 4594 3261 4606 3295
rect 4548 3227 4606 3261
rect 4548 3193 4560 3227
rect 4594 3193 4606 3227
rect 4548 3159 4606 3193
rect 4548 3125 4560 3159
rect 4594 3125 4606 3159
rect 4548 3110 4606 3125
rect 4698 3295 4756 3310
rect 4698 3261 4710 3295
rect 4744 3261 4756 3295
rect 4698 3227 4756 3261
rect 4698 3193 4710 3227
rect 4744 3193 4756 3227
rect 4698 3159 4756 3193
rect 4698 3125 4710 3159
rect 4744 3125 4756 3159
rect 4698 3110 4756 3125
rect 4856 3295 4914 3310
rect 4856 3261 4868 3295
rect 4902 3261 4914 3295
rect 4856 3227 4914 3261
rect 4856 3193 4868 3227
rect 4902 3193 4914 3227
rect 4856 3159 4914 3193
rect 4856 3125 4868 3159
rect 4902 3125 4914 3159
rect 4856 3110 4914 3125
rect 5688 3296 5746 3310
rect 5688 3262 5700 3296
rect 5734 3262 5746 3296
rect 5688 3228 5746 3262
rect 5688 3194 5700 3228
rect 5734 3194 5746 3228
rect 5688 3160 5746 3194
rect 5688 3126 5700 3160
rect 5734 3126 5746 3160
rect 5688 3110 5746 3126
rect 5846 3296 5904 3310
rect 5846 3262 5858 3296
rect 5892 3262 5904 3296
rect 5846 3228 5904 3262
rect 5846 3194 5858 3228
rect 5892 3194 5904 3228
rect 5846 3160 5904 3194
rect 5846 3126 5858 3160
rect 5892 3126 5904 3160
rect 5846 3110 5904 3126
rect 5996 3296 6054 3310
rect 5996 3262 6008 3296
rect 6042 3262 6054 3296
rect 5996 3228 6054 3262
rect 5996 3194 6008 3228
rect 6042 3194 6054 3228
rect 5996 3160 6054 3194
rect 5996 3126 6008 3160
rect 6042 3126 6054 3160
rect 5996 3110 6054 3126
rect 6154 3296 6212 3310
rect 6154 3262 6166 3296
rect 6200 3262 6212 3296
rect 6154 3228 6212 3262
rect 6154 3194 6166 3228
rect 6200 3194 6212 3228
rect 6154 3160 6212 3194
rect 6154 3126 6166 3160
rect 6200 3126 6212 3160
rect 6154 3110 6212 3126
rect 6348 3296 6406 3310
rect 6348 3262 6360 3296
rect 6394 3262 6406 3296
rect 6348 3228 6406 3262
rect 6348 3194 6360 3228
rect 6394 3194 6406 3228
rect 6348 3160 6406 3194
rect 6348 3126 6360 3160
rect 6394 3126 6406 3160
rect 6348 3110 6406 3126
rect 6506 3296 6564 3310
rect 6506 3262 6518 3296
rect 6552 3262 6564 3296
rect 6506 3228 6564 3262
rect 6506 3194 6518 3228
rect 6552 3194 6564 3228
rect 6506 3160 6564 3194
rect 6506 3126 6518 3160
rect 6552 3126 6564 3160
rect 6506 3110 6564 3126
rect 6656 3296 6714 3310
rect 6656 3262 6668 3296
rect 6702 3262 6714 3296
rect 6656 3228 6714 3262
rect 6656 3194 6668 3228
rect 6702 3194 6714 3228
rect 6656 3160 6714 3194
rect 6656 3126 6668 3160
rect 6702 3126 6714 3160
rect 6656 3110 6714 3126
rect 6814 3296 6872 3310
rect 6814 3262 6826 3296
rect 6860 3262 6872 3296
rect 6814 3228 6872 3262
rect 6814 3194 6826 3228
rect 6860 3194 6872 3228
rect 6814 3160 6872 3194
rect 6814 3126 6826 3160
rect 6860 3126 6872 3160
rect 6814 3110 6872 3126
rect 1398 2057 1456 2072
rect 1398 2023 1410 2057
rect 1444 2023 1456 2057
rect 1398 1989 1456 2023
rect 1398 1955 1410 1989
rect 1444 1955 1456 1989
rect 1398 1921 1456 1955
rect 1398 1887 1410 1921
rect 1444 1887 1456 1921
rect 1398 1872 1456 1887
rect 1556 2057 1614 2072
rect 1556 2023 1568 2057
rect 1602 2023 1614 2057
rect 1556 1989 1614 2023
rect 1556 1955 1568 1989
rect 1602 1955 1614 1989
rect 1556 1921 1614 1955
rect 1556 1887 1568 1921
rect 1602 1887 1614 1921
rect 1556 1872 1614 1887
rect 1686 2057 1744 2072
rect 1686 2023 1698 2057
rect 1732 2023 1744 2057
rect 1686 1989 1744 2023
rect 1686 1955 1698 1989
rect 1732 1955 1744 1989
rect 1686 1921 1744 1955
rect 1686 1887 1698 1921
rect 1732 1887 1744 1921
rect 1686 1872 1744 1887
rect 1844 2057 1902 2072
rect 1844 2023 1856 2057
rect 1890 2023 1902 2057
rect 1844 1989 1902 2023
rect 1844 1955 1856 1989
rect 1890 1955 1902 1989
rect 1844 1921 1902 1955
rect 1844 1887 1856 1921
rect 1890 1887 1902 1921
rect 1844 1872 1902 1887
rect 2018 2057 2076 2072
rect 2018 2023 2030 2057
rect 2064 2023 2076 2057
rect 2018 1989 2076 2023
rect 2018 1955 2030 1989
rect 2064 1955 2076 1989
rect 2018 1921 2076 1955
rect 2018 1887 2030 1921
rect 2064 1887 2076 1921
rect 2018 1872 2076 1887
rect 2176 2057 2234 2072
rect 2176 2023 2188 2057
rect 2222 2023 2234 2057
rect 2176 1989 2234 2023
rect 2176 1955 2188 1989
rect 2222 1955 2234 1989
rect 2176 1921 2234 1955
rect 2176 1887 2188 1921
rect 2222 1887 2234 1921
rect 2176 1872 2234 1887
rect 2360 2057 2418 2072
rect 2360 2023 2372 2057
rect 2406 2023 2418 2057
rect 2360 1989 2418 2023
rect 2360 1955 2372 1989
rect 2406 1955 2418 1989
rect 2360 1921 2418 1955
rect 2360 1887 2372 1921
rect 2406 1887 2418 1921
rect 2360 1872 2418 1887
rect 2518 2057 2576 2072
rect 2518 2023 2530 2057
rect 2564 2023 2576 2057
rect 2518 1989 2576 2023
rect 2518 1955 2530 1989
rect 2564 1955 2576 1989
rect 2518 1921 2576 1955
rect 2518 1887 2530 1921
rect 2564 1887 2576 1921
rect 2518 1872 2576 1887
rect 2764 2057 2822 2072
rect 2764 2023 2776 2057
rect 2810 2023 2822 2057
rect 2764 1989 2822 2023
rect 2764 1955 2776 1989
rect 2810 1955 2822 1989
rect 2764 1921 2822 1955
rect 2764 1887 2776 1921
rect 2810 1887 2822 1921
rect 2764 1872 2822 1887
rect 2922 2057 2980 2072
rect 2922 2023 2934 2057
rect 2968 2023 2980 2057
rect 2922 1989 2980 2023
rect 2922 1955 2934 1989
rect 2968 1955 2980 1989
rect 2922 1921 2980 1955
rect 2922 1887 2934 1921
rect 2968 1887 2980 1921
rect 2922 1872 2980 1887
rect 3108 2057 3166 2072
rect 3108 2023 3120 2057
rect 3154 2023 3166 2057
rect 3108 1989 3166 2023
rect 3108 1955 3120 1989
rect 3154 1955 3166 1989
rect 3108 1921 3166 1955
rect 3108 1887 3120 1921
rect 3154 1887 3166 1921
rect 3108 1872 3166 1887
rect 3266 2057 3324 2072
rect 3266 2023 3278 2057
rect 3312 2023 3324 2057
rect 3266 1989 3324 2023
rect 3266 1955 3278 1989
rect 3312 1955 3324 1989
rect 3266 1921 3324 1955
rect 3266 1887 3278 1921
rect 3312 1887 3324 1921
rect 3266 1872 3324 1887
rect 3730 2067 3788 2082
rect 3730 2033 3742 2067
rect 3776 2033 3788 2067
rect 3730 1999 3788 2033
rect 3730 1965 3742 1999
rect 3776 1965 3788 1999
rect 3730 1931 3788 1965
rect 3730 1897 3742 1931
rect 3776 1897 3788 1931
rect 3730 1882 3788 1897
rect 3888 2067 3946 2082
rect 3888 2033 3900 2067
rect 3934 2033 3946 2067
rect 3888 1999 3946 2033
rect 3888 1965 3900 1999
rect 3934 1965 3946 1999
rect 3888 1931 3946 1965
rect 3888 1897 3900 1931
rect 3934 1897 3946 1931
rect 3888 1882 3946 1897
rect 4038 2067 4096 2082
rect 4038 2033 4050 2067
rect 4084 2033 4096 2067
rect 4038 1999 4096 2033
rect 4038 1965 4050 1999
rect 4084 1965 4096 1999
rect 4038 1931 4096 1965
rect 4038 1897 4050 1931
rect 4084 1897 4096 1931
rect 4038 1882 4096 1897
rect 4196 2067 4254 2082
rect 4196 2033 4208 2067
rect 4242 2033 4254 2067
rect 4196 1999 4254 2033
rect 4196 1965 4208 1999
rect 4242 1965 4254 1999
rect 4196 1931 4254 1965
rect 4196 1897 4208 1931
rect 4242 1897 4254 1931
rect 4196 1882 4254 1897
rect 4390 2067 4448 2082
rect 4390 2033 4402 2067
rect 4436 2033 4448 2067
rect 4390 1999 4448 2033
rect 4390 1965 4402 1999
rect 4436 1965 4448 1999
rect 4390 1931 4448 1965
rect 4390 1897 4402 1931
rect 4436 1897 4448 1931
rect 4390 1882 4448 1897
rect 4548 2067 4606 2082
rect 4548 2033 4560 2067
rect 4594 2033 4606 2067
rect 4548 1999 4606 2033
rect 4548 1965 4560 1999
rect 4594 1965 4606 1999
rect 4548 1931 4606 1965
rect 4548 1897 4560 1931
rect 4594 1897 4606 1931
rect 4548 1882 4606 1897
rect 4698 2067 4756 2082
rect 4698 2033 4710 2067
rect 4744 2033 4756 2067
rect 4698 1999 4756 2033
rect 4698 1965 4710 1999
rect 4744 1965 4756 1999
rect 4698 1931 4756 1965
rect 4698 1897 4710 1931
rect 4744 1897 4756 1931
rect 4698 1882 4756 1897
rect 4856 2067 4914 2082
rect 4856 2033 4868 2067
rect 4902 2033 4914 2067
rect 4856 1999 4914 2033
rect 4856 1965 4868 1999
rect 4902 1965 4914 1999
rect 4856 1931 4914 1965
rect 4856 1897 4868 1931
rect 4902 1897 4914 1931
rect 4856 1882 4914 1897
rect 5688 2068 5746 2082
rect 5688 2034 5700 2068
rect 5734 2034 5746 2068
rect 5688 2000 5746 2034
rect 5688 1966 5700 2000
rect 5734 1966 5746 2000
rect 5688 1932 5746 1966
rect 5688 1898 5700 1932
rect 5734 1898 5746 1932
rect 5688 1882 5746 1898
rect 5846 2068 5904 2082
rect 5846 2034 5858 2068
rect 5892 2034 5904 2068
rect 5846 2000 5904 2034
rect 5846 1966 5858 2000
rect 5892 1966 5904 2000
rect 5846 1932 5904 1966
rect 5846 1898 5858 1932
rect 5892 1898 5904 1932
rect 5846 1882 5904 1898
rect 5996 2068 6054 2082
rect 5996 2034 6008 2068
rect 6042 2034 6054 2068
rect 5996 2000 6054 2034
rect 5996 1966 6008 2000
rect 6042 1966 6054 2000
rect 5996 1932 6054 1966
rect 5996 1898 6008 1932
rect 6042 1898 6054 1932
rect 5996 1882 6054 1898
rect 6154 2068 6212 2082
rect 6154 2034 6166 2068
rect 6200 2034 6212 2068
rect 6154 2000 6212 2034
rect 6154 1966 6166 2000
rect 6200 1966 6212 2000
rect 6154 1932 6212 1966
rect 6154 1898 6166 1932
rect 6200 1898 6212 1932
rect 6154 1882 6212 1898
rect 6348 2068 6406 2082
rect 6348 2034 6360 2068
rect 6394 2034 6406 2068
rect 6348 2000 6406 2034
rect 6348 1966 6360 2000
rect 6394 1966 6406 2000
rect 6348 1932 6406 1966
rect 6348 1898 6360 1932
rect 6394 1898 6406 1932
rect 6348 1882 6406 1898
rect 6506 2068 6564 2082
rect 6506 2034 6518 2068
rect 6552 2034 6564 2068
rect 6506 2000 6564 2034
rect 6506 1966 6518 2000
rect 6552 1966 6564 2000
rect 6506 1932 6564 1966
rect 6506 1898 6518 1932
rect 6552 1898 6564 1932
rect 6506 1882 6564 1898
rect 6656 2068 6714 2082
rect 6656 2034 6668 2068
rect 6702 2034 6714 2068
rect 6656 2000 6714 2034
rect 6656 1966 6668 2000
rect 6702 1966 6714 2000
rect 6656 1932 6714 1966
rect 6656 1898 6668 1932
rect 6702 1898 6714 1932
rect 6656 1882 6714 1898
rect 6814 2068 6872 2082
rect 6814 2034 6826 2068
rect 6860 2034 6872 2068
rect 6814 2000 6872 2034
rect 6814 1966 6826 2000
rect 6860 1966 6872 2000
rect 6814 1932 6872 1966
rect 6814 1898 6826 1932
rect 6860 1898 6872 1932
rect 6814 1882 6872 1898
rect 1398 829 1456 844
rect 1398 795 1410 829
rect 1444 795 1456 829
rect 1398 761 1456 795
rect 1398 727 1410 761
rect 1444 727 1456 761
rect 1398 693 1456 727
rect 1398 659 1410 693
rect 1444 659 1456 693
rect 1398 644 1456 659
rect 1556 829 1614 844
rect 1556 795 1568 829
rect 1602 795 1614 829
rect 1556 761 1614 795
rect 1556 727 1568 761
rect 1602 727 1614 761
rect 1556 693 1614 727
rect 1556 659 1568 693
rect 1602 659 1614 693
rect 1556 644 1614 659
rect 1686 829 1744 844
rect 1686 795 1698 829
rect 1732 795 1744 829
rect 1686 761 1744 795
rect 1686 727 1698 761
rect 1732 727 1744 761
rect 1686 693 1744 727
rect 1686 659 1698 693
rect 1732 659 1744 693
rect 1686 644 1744 659
rect 1844 829 1902 844
rect 1844 795 1856 829
rect 1890 795 1902 829
rect 1844 761 1902 795
rect 1844 727 1856 761
rect 1890 727 1902 761
rect 1844 693 1902 727
rect 1844 659 1856 693
rect 1890 659 1902 693
rect 1844 644 1902 659
rect 2018 829 2076 844
rect 2018 795 2030 829
rect 2064 795 2076 829
rect 2018 761 2076 795
rect 2018 727 2030 761
rect 2064 727 2076 761
rect 2018 693 2076 727
rect 2018 659 2030 693
rect 2064 659 2076 693
rect 2018 644 2076 659
rect 2176 829 2234 844
rect 2176 795 2188 829
rect 2222 795 2234 829
rect 2176 761 2234 795
rect 2176 727 2188 761
rect 2222 727 2234 761
rect 2176 693 2234 727
rect 2176 659 2188 693
rect 2222 659 2234 693
rect 2176 644 2234 659
rect 2360 829 2418 844
rect 2360 795 2372 829
rect 2406 795 2418 829
rect 2360 761 2418 795
rect 2360 727 2372 761
rect 2406 727 2418 761
rect 2360 693 2418 727
rect 2360 659 2372 693
rect 2406 659 2418 693
rect 2360 644 2418 659
rect 2518 829 2576 844
rect 2518 795 2530 829
rect 2564 795 2576 829
rect 2518 761 2576 795
rect 2518 727 2530 761
rect 2564 727 2576 761
rect 2518 693 2576 727
rect 2518 659 2530 693
rect 2564 659 2576 693
rect 2518 644 2576 659
rect 2764 829 2822 844
rect 2764 795 2776 829
rect 2810 795 2822 829
rect 2764 761 2822 795
rect 2764 727 2776 761
rect 2810 727 2822 761
rect 2764 693 2822 727
rect 2764 659 2776 693
rect 2810 659 2822 693
rect 2764 644 2822 659
rect 2922 829 2980 844
rect 2922 795 2934 829
rect 2968 795 2980 829
rect 2922 761 2980 795
rect 2922 727 2934 761
rect 2968 727 2980 761
rect 2922 693 2980 727
rect 2922 659 2934 693
rect 2968 659 2980 693
rect 2922 644 2980 659
rect 3108 829 3166 844
rect 3108 795 3120 829
rect 3154 795 3166 829
rect 3108 761 3166 795
rect 3108 727 3120 761
rect 3154 727 3166 761
rect 3108 693 3166 727
rect 3108 659 3120 693
rect 3154 659 3166 693
rect 3108 644 3166 659
rect 3266 829 3324 844
rect 3266 795 3278 829
rect 3312 795 3324 829
rect 3266 761 3324 795
rect 3266 727 3278 761
rect 3312 727 3324 761
rect 3266 693 3324 727
rect 3266 659 3278 693
rect 3312 659 3324 693
rect 3266 644 3324 659
rect 3730 839 3788 854
rect 3730 805 3742 839
rect 3776 805 3788 839
rect 3730 771 3788 805
rect 3730 737 3742 771
rect 3776 737 3788 771
rect 3730 703 3788 737
rect 3730 669 3742 703
rect 3776 669 3788 703
rect 3730 654 3788 669
rect 3888 839 3946 854
rect 3888 805 3900 839
rect 3934 805 3946 839
rect 3888 771 3946 805
rect 3888 737 3900 771
rect 3934 737 3946 771
rect 3888 703 3946 737
rect 3888 669 3900 703
rect 3934 669 3946 703
rect 3888 654 3946 669
rect 4038 839 4096 854
rect 4038 805 4050 839
rect 4084 805 4096 839
rect 4038 771 4096 805
rect 4038 737 4050 771
rect 4084 737 4096 771
rect 4038 703 4096 737
rect 4038 669 4050 703
rect 4084 669 4096 703
rect 4038 654 4096 669
rect 4196 839 4254 854
rect 4196 805 4208 839
rect 4242 805 4254 839
rect 4196 771 4254 805
rect 4196 737 4208 771
rect 4242 737 4254 771
rect 4196 703 4254 737
rect 4196 669 4208 703
rect 4242 669 4254 703
rect 4196 654 4254 669
rect 4390 839 4448 854
rect 4390 805 4402 839
rect 4436 805 4448 839
rect 4390 771 4448 805
rect 4390 737 4402 771
rect 4436 737 4448 771
rect 4390 703 4448 737
rect 4390 669 4402 703
rect 4436 669 4448 703
rect 4390 654 4448 669
rect 4548 839 4606 854
rect 4548 805 4560 839
rect 4594 805 4606 839
rect 4548 771 4606 805
rect 4548 737 4560 771
rect 4594 737 4606 771
rect 4548 703 4606 737
rect 4548 669 4560 703
rect 4594 669 4606 703
rect 4548 654 4606 669
rect 4698 839 4756 854
rect 4698 805 4710 839
rect 4744 805 4756 839
rect 4698 771 4756 805
rect 4698 737 4710 771
rect 4744 737 4756 771
rect 4698 703 4756 737
rect 4698 669 4710 703
rect 4744 669 4756 703
rect 4698 654 4756 669
rect 4856 839 4914 854
rect 4856 805 4868 839
rect 4902 805 4914 839
rect 4856 771 4914 805
rect 4856 737 4868 771
rect 4902 737 4914 771
rect 4856 703 4914 737
rect 4856 669 4868 703
rect 4902 669 4914 703
rect 4856 654 4914 669
<< mvndiffc >>
rect 569 4578 603 4612
rect 569 4010 603 4044
rect 715 4578 749 4612
rect 715 4010 749 4044
rect 859 4584 893 4618
rect 859 4016 893 4050
rect 1013 4584 1047 4618
rect 1410 4123 1444 4157
rect 1568 4123 1602 4157
rect 1698 4123 1732 4157
rect 1856 4123 1890 4157
rect 2030 4123 2064 4157
rect 2188 4123 2222 4157
rect 2372 4123 2406 4157
rect 2530 4123 2564 4157
rect 2776 4123 2810 4157
rect 2934 4123 2968 4157
rect 3120 4123 3154 4157
rect 3278 4123 3312 4157
rect 3742 4133 3776 4167
rect 3900 4133 3934 4167
rect 4050 4133 4084 4167
rect 4208 4133 4242 4167
rect 4402 4135 4436 4169
rect 4560 4135 4594 4169
rect 4710 4135 4744 4169
rect 4868 4135 4902 4169
rect 5700 4134 5734 4168
rect 5858 4134 5892 4168
rect 6008 4134 6042 4168
rect 6166 4134 6200 4168
rect 6360 4136 6394 4170
rect 6518 4136 6552 4170
rect 6668 4136 6702 4170
rect 6826 4136 6860 4170
rect 1013 4016 1047 4050
rect 569 3350 603 3384
rect 569 2782 603 2816
rect 715 3350 749 3384
rect 715 2782 749 2816
rect 859 3356 893 3390
rect 859 2788 893 2822
rect 1013 3356 1047 3390
rect 1410 2895 1444 2929
rect 1568 2895 1602 2929
rect 1698 2895 1732 2929
rect 1856 2895 1890 2929
rect 2030 2895 2064 2929
rect 2188 2895 2222 2929
rect 2372 2895 2406 2929
rect 2530 2895 2564 2929
rect 2776 2895 2810 2929
rect 2934 2895 2968 2929
rect 3120 2895 3154 2929
rect 3278 2895 3312 2929
rect 3742 2905 3776 2939
rect 3900 2905 3934 2939
rect 4050 2905 4084 2939
rect 4208 2905 4242 2939
rect 4402 2907 4436 2941
rect 4560 2907 4594 2941
rect 4710 2907 4744 2941
rect 4868 2907 4902 2941
rect 5700 2906 5734 2940
rect 5858 2906 5892 2940
rect 6008 2906 6042 2940
rect 6166 2906 6200 2940
rect 6360 2908 6394 2942
rect 6518 2908 6552 2942
rect 6668 2908 6702 2942
rect 6826 2908 6860 2942
rect 1013 2788 1047 2822
rect 569 2122 603 2156
rect 569 1554 603 1588
rect 715 2122 749 2156
rect 715 1554 749 1588
rect 859 2128 893 2162
rect 859 1560 893 1594
rect 1013 2128 1047 2162
rect 1410 1667 1444 1701
rect 1568 1667 1602 1701
rect 1698 1667 1732 1701
rect 1856 1667 1890 1701
rect 2030 1667 2064 1701
rect 2188 1667 2222 1701
rect 2372 1667 2406 1701
rect 2530 1667 2564 1701
rect 2776 1667 2810 1701
rect 2934 1667 2968 1701
rect 3120 1667 3154 1701
rect 3278 1667 3312 1701
rect 3742 1677 3776 1711
rect 3900 1677 3934 1711
rect 4050 1677 4084 1711
rect 4208 1677 4242 1711
rect 4402 1679 4436 1713
rect 4560 1679 4594 1713
rect 4710 1679 4744 1713
rect 4868 1679 4902 1713
rect 5700 1678 5734 1712
rect 5858 1678 5892 1712
rect 6008 1678 6042 1712
rect 6166 1678 6200 1712
rect 6360 1680 6394 1714
rect 6518 1680 6552 1714
rect 6668 1680 6702 1714
rect 6826 1680 6860 1714
rect 1013 1560 1047 1594
rect 569 894 603 928
rect 569 326 603 360
rect 715 894 749 928
rect 715 326 749 360
rect 859 900 893 934
rect 859 332 893 366
rect 1013 900 1047 934
rect 1410 439 1444 473
rect 1568 439 1602 473
rect 1698 439 1732 473
rect 1856 439 1890 473
rect 2030 439 2064 473
rect 2188 439 2222 473
rect 2372 439 2406 473
rect 2530 439 2564 473
rect 2776 439 2810 473
rect 2934 439 2968 473
rect 3120 439 3154 473
rect 3278 439 3312 473
rect 3742 449 3776 483
rect 3900 449 3934 483
rect 4050 449 4084 483
rect 4208 449 4242 483
rect 4402 451 4436 485
rect 4560 451 4594 485
rect 4710 451 4744 485
rect 4868 451 4902 485
rect 1013 332 1047 366
<< mvpdiffc >>
rect 1410 4479 1444 4513
rect 1410 4411 1444 4445
rect 1410 4343 1444 4377
rect 1568 4479 1602 4513
rect 1568 4411 1602 4445
rect 1568 4343 1602 4377
rect 1698 4479 1732 4513
rect 1698 4411 1732 4445
rect 1698 4343 1732 4377
rect 1856 4479 1890 4513
rect 1856 4411 1890 4445
rect 1856 4343 1890 4377
rect 2030 4479 2064 4513
rect 2030 4411 2064 4445
rect 2030 4343 2064 4377
rect 2188 4479 2222 4513
rect 2188 4411 2222 4445
rect 2188 4343 2222 4377
rect 2372 4479 2406 4513
rect 2372 4411 2406 4445
rect 2372 4343 2406 4377
rect 2530 4479 2564 4513
rect 2530 4411 2564 4445
rect 2530 4343 2564 4377
rect 2776 4479 2810 4513
rect 2776 4411 2810 4445
rect 2776 4343 2810 4377
rect 2934 4479 2968 4513
rect 2934 4411 2968 4445
rect 2934 4343 2968 4377
rect 3120 4479 3154 4513
rect 3120 4411 3154 4445
rect 3120 4343 3154 4377
rect 3278 4479 3312 4513
rect 3278 4411 3312 4445
rect 3278 4343 3312 4377
rect 3742 4489 3776 4523
rect 3742 4421 3776 4455
rect 3742 4353 3776 4387
rect 3900 4489 3934 4523
rect 3900 4421 3934 4455
rect 3900 4353 3934 4387
rect 4050 4489 4084 4523
rect 4050 4421 4084 4455
rect 4050 4353 4084 4387
rect 4208 4489 4242 4523
rect 4208 4421 4242 4455
rect 4208 4353 4242 4387
rect 4402 4489 4436 4523
rect 4402 4421 4436 4455
rect 4402 4353 4436 4387
rect 4560 4489 4594 4523
rect 4560 4421 4594 4455
rect 4560 4353 4594 4387
rect 4710 4489 4744 4523
rect 4710 4421 4744 4455
rect 4710 4353 4744 4387
rect 4868 4489 4902 4523
rect 4868 4421 4902 4455
rect 4868 4353 4902 4387
rect 5700 4490 5734 4524
rect 5700 4422 5734 4456
rect 5700 4354 5734 4388
rect 5858 4490 5892 4524
rect 5858 4422 5892 4456
rect 5858 4354 5892 4388
rect 6008 4490 6042 4524
rect 6008 4422 6042 4456
rect 6008 4354 6042 4388
rect 6166 4490 6200 4524
rect 6166 4422 6200 4456
rect 6166 4354 6200 4388
rect 6360 4490 6394 4524
rect 6360 4422 6394 4456
rect 6360 4354 6394 4388
rect 6518 4490 6552 4524
rect 6518 4422 6552 4456
rect 6518 4354 6552 4388
rect 6668 4490 6702 4524
rect 6668 4422 6702 4456
rect 6668 4354 6702 4388
rect 6826 4490 6860 4524
rect 6826 4422 6860 4456
rect 6826 4354 6860 4388
rect 1410 3251 1444 3285
rect 1410 3183 1444 3217
rect 1410 3115 1444 3149
rect 1568 3251 1602 3285
rect 1568 3183 1602 3217
rect 1568 3115 1602 3149
rect 1698 3251 1732 3285
rect 1698 3183 1732 3217
rect 1698 3115 1732 3149
rect 1856 3251 1890 3285
rect 1856 3183 1890 3217
rect 1856 3115 1890 3149
rect 2030 3251 2064 3285
rect 2030 3183 2064 3217
rect 2030 3115 2064 3149
rect 2188 3251 2222 3285
rect 2188 3183 2222 3217
rect 2188 3115 2222 3149
rect 2372 3251 2406 3285
rect 2372 3183 2406 3217
rect 2372 3115 2406 3149
rect 2530 3251 2564 3285
rect 2530 3183 2564 3217
rect 2530 3115 2564 3149
rect 2776 3251 2810 3285
rect 2776 3183 2810 3217
rect 2776 3115 2810 3149
rect 2934 3251 2968 3285
rect 2934 3183 2968 3217
rect 2934 3115 2968 3149
rect 3120 3251 3154 3285
rect 3120 3183 3154 3217
rect 3120 3115 3154 3149
rect 3278 3251 3312 3285
rect 3278 3183 3312 3217
rect 3278 3115 3312 3149
rect 3742 3261 3776 3295
rect 3742 3193 3776 3227
rect 3742 3125 3776 3159
rect 3900 3261 3934 3295
rect 3900 3193 3934 3227
rect 3900 3125 3934 3159
rect 4050 3261 4084 3295
rect 4050 3193 4084 3227
rect 4050 3125 4084 3159
rect 4208 3261 4242 3295
rect 4208 3193 4242 3227
rect 4208 3125 4242 3159
rect 4402 3261 4436 3295
rect 4402 3193 4436 3227
rect 4402 3125 4436 3159
rect 4560 3261 4594 3295
rect 4560 3193 4594 3227
rect 4560 3125 4594 3159
rect 4710 3261 4744 3295
rect 4710 3193 4744 3227
rect 4710 3125 4744 3159
rect 4868 3261 4902 3295
rect 4868 3193 4902 3227
rect 4868 3125 4902 3159
rect 5700 3262 5734 3296
rect 5700 3194 5734 3228
rect 5700 3126 5734 3160
rect 5858 3262 5892 3296
rect 5858 3194 5892 3228
rect 5858 3126 5892 3160
rect 6008 3262 6042 3296
rect 6008 3194 6042 3228
rect 6008 3126 6042 3160
rect 6166 3262 6200 3296
rect 6166 3194 6200 3228
rect 6166 3126 6200 3160
rect 6360 3262 6394 3296
rect 6360 3194 6394 3228
rect 6360 3126 6394 3160
rect 6518 3262 6552 3296
rect 6518 3194 6552 3228
rect 6518 3126 6552 3160
rect 6668 3262 6702 3296
rect 6668 3194 6702 3228
rect 6668 3126 6702 3160
rect 6826 3262 6860 3296
rect 6826 3194 6860 3228
rect 6826 3126 6860 3160
rect 1410 2023 1444 2057
rect 1410 1955 1444 1989
rect 1410 1887 1444 1921
rect 1568 2023 1602 2057
rect 1568 1955 1602 1989
rect 1568 1887 1602 1921
rect 1698 2023 1732 2057
rect 1698 1955 1732 1989
rect 1698 1887 1732 1921
rect 1856 2023 1890 2057
rect 1856 1955 1890 1989
rect 1856 1887 1890 1921
rect 2030 2023 2064 2057
rect 2030 1955 2064 1989
rect 2030 1887 2064 1921
rect 2188 2023 2222 2057
rect 2188 1955 2222 1989
rect 2188 1887 2222 1921
rect 2372 2023 2406 2057
rect 2372 1955 2406 1989
rect 2372 1887 2406 1921
rect 2530 2023 2564 2057
rect 2530 1955 2564 1989
rect 2530 1887 2564 1921
rect 2776 2023 2810 2057
rect 2776 1955 2810 1989
rect 2776 1887 2810 1921
rect 2934 2023 2968 2057
rect 2934 1955 2968 1989
rect 2934 1887 2968 1921
rect 3120 2023 3154 2057
rect 3120 1955 3154 1989
rect 3120 1887 3154 1921
rect 3278 2023 3312 2057
rect 3278 1955 3312 1989
rect 3278 1887 3312 1921
rect 3742 2033 3776 2067
rect 3742 1965 3776 1999
rect 3742 1897 3776 1931
rect 3900 2033 3934 2067
rect 3900 1965 3934 1999
rect 3900 1897 3934 1931
rect 4050 2033 4084 2067
rect 4050 1965 4084 1999
rect 4050 1897 4084 1931
rect 4208 2033 4242 2067
rect 4208 1965 4242 1999
rect 4208 1897 4242 1931
rect 4402 2033 4436 2067
rect 4402 1965 4436 1999
rect 4402 1897 4436 1931
rect 4560 2033 4594 2067
rect 4560 1965 4594 1999
rect 4560 1897 4594 1931
rect 4710 2033 4744 2067
rect 4710 1965 4744 1999
rect 4710 1897 4744 1931
rect 4868 2033 4902 2067
rect 4868 1965 4902 1999
rect 4868 1897 4902 1931
rect 5700 2034 5734 2068
rect 5700 1966 5734 2000
rect 5700 1898 5734 1932
rect 5858 2034 5892 2068
rect 5858 1966 5892 2000
rect 5858 1898 5892 1932
rect 6008 2034 6042 2068
rect 6008 1966 6042 2000
rect 6008 1898 6042 1932
rect 6166 2034 6200 2068
rect 6166 1966 6200 2000
rect 6166 1898 6200 1932
rect 6360 2034 6394 2068
rect 6360 1966 6394 2000
rect 6360 1898 6394 1932
rect 6518 2034 6552 2068
rect 6518 1966 6552 2000
rect 6518 1898 6552 1932
rect 6668 2034 6702 2068
rect 6668 1966 6702 2000
rect 6668 1898 6702 1932
rect 6826 2034 6860 2068
rect 6826 1966 6860 2000
rect 6826 1898 6860 1932
rect 1410 795 1444 829
rect 1410 727 1444 761
rect 1410 659 1444 693
rect 1568 795 1602 829
rect 1568 727 1602 761
rect 1568 659 1602 693
rect 1698 795 1732 829
rect 1698 727 1732 761
rect 1698 659 1732 693
rect 1856 795 1890 829
rect 1856 727 1890 761
rect 1856 659 1890 693
rect 2030 795 2064 829
rect 2030 727 2064 761
rect 2030 659 2064 693
rect 2188 795 2222 829
rect 2188 727 2222 761
rect 2188 659 2222 693
rect 2372 795 2406 829
rect 2372 727 2406 761
rect 2372 659 2406 693
rect 2530 795 2564 829
rect 2530 727 2564 761
rect 2530 659 2564 693
rect 2776 795 2810 829
rect 2776 727 2810 761
rect 2776 659 2810 693
rect 2934 795 2968 829
rect 2934 727 2968 761
rect 2934 659 2968 693
rect 3120 795 3154 829
rect 3120 727 3154 761
rect 3120 659 3154 693
rect 3278 795 3312 829
rect 3278 727 3312 761
rect 3278 659 3312 693
rect 3742 805 3776 839
rect 3742 737 3776 771
rect 3742 669 3776 703
rect 3900 805 3934 839
rect 3900 737 3934 771
rect 3900 669 3934 703
rect 4050 805 4084 839
rect 4050 737 4084 771
rect 4050 669 4084 703
rect 4208 805 4242 839
rect 4208 737 4242 771
rect 4208 669 4242 703
rect 4402 805 4436 839
rect 4402 737 4436 771
rect 4402 669 4436 703
rect 4560 805 4594 839
rect 4560 737 4594 771
rect 4560 669 4594 703
rect 4710 805 4744 839
rect 4710 737 4744 771
rect 4710 669 4744 703
rect 4868 805 4902 839
rect 4868 737 4902 771
rect 4868 669 4902 703
<< psubdiff >>
rect 1324 3980 1959 4032
rect 1324 3946 1353 3980
rect 1387 3946 1421 3980
rect 1455 3946 1489 3980
rect 1523 3946 1557 3980
rect 1591 3946 1625 3980
rect 1659 3946 1693 3980
rect 1727 3946 1761 3980
rect 1795 3946 1829 3980
rect 1863 3946 1897 3980
rect 1931 3946 1959 3980
rect 1324 3904 1959 3946
rect 3704 3991 4244 4044
rect 3704 3957 3753 3991
rect 3787 3957 3821 3991
rect 3855 3957 3889 3991
rect 3923 3957 3957 3991
rect 3991 3957 4025 3991
rect 4059 3957 4093 3991
rect 4127 3957 4161 3991
rect 4195 3957 4244 3991
rect 3704 3904 4244 3957
rect 5662 3992 6202 4044
rect 5662 3958 5712 3992
rect 5746 3958 5780 3992
rect 5814 3958 5848 3992
rect 5882 3958 5916 3992
rect 5950 3958 5984 3992
rect 6018 3958 6052 3992
rect 6086 3958 6120 3992
rect 6154 3958 6202 3992
rect 5662 3904 6202 3958
rect 1324 2752 1959 2804
rect 1324 2718 1353 2752
rect 1387 2718 1421 2752
rect 1455 2718 1489 2752
rect 1523 2718 1557 2752
rect 1591 2718 1625 2752
rect 1659 2718 1693 2752
rect 1727 2718 1761 2752
rect 1795 2718 1829 2752
rect 1863 2718 1897 2752
rect 1931 2718 1959 2752
rect 1324 2676 1959 2718
rect 3704 2763 4244 2816
rect 3704 2729 3753 2763
rect 3787 2729 3821 2763
rect 3855 2729 3889 2763
rect 3923 2729 3957 2763
rect 3991 2729 4025 2763
rect 4059 2729 4093 2763
rect 4127 2729 4161 2763
rect 4195 2729 4244 2763
rect 3704 2676 4244 2729
rect 5662 2764 6202 2816
rect 5662 2730 5712 2764
rect 5746 2730 5780 2764
rect 5814 2730 5848 2764
rect 5882 2730 5916 2764
rect 5950 2730 5984 2764
rect 6018 2730 6052 2764
rect 6086 2730 6120 2764
rect 6154 2730 6202 2764
rect 5662 2676 6202 2730
rect 1324 1524 1959 1576
rect 1324 1490 1353 1524
rect 1387 1490 1421 1524
rect 1455 1490 1489 1524
rect 1523 1490 1557 1524
rect 1591 1490 1625 1524
rect 1659 1490 1693 1524
rect 1727 1490 1761 1524
rect 1795 1490 1829 1524
rect 1863 1490 1897 1524
rect 1931 1490 1959 1524
rect 1324 1448 1959 1490
rect 3704 1535 4244 1588
rect 3704 1501 3753 1535
rect 3787 1501 3821 1535
rect 3855 1501 3889 1535
rect 3923 1501 3957 1535
rect 3991 1501 4025 1535
rect 4059 1501 4093 1535
rect 4127 1501 4161 1535
rect 4195 1501 4244 1535
rect 3704 1448 4244 1501
rect 5662 1536 6202 1588
rect 5662 1502 5712 1536
rect 5746 1502 5780 1536
rect 5814 1502 5848 1536
rect 5882 1502 5916 1536
rect 5950 1502 5984 1536
rect 6018 1502 6052 1536
rect 6086 1502 6120 1536
rect 6154 1502 6202 1536
rect 5662 1448 6202 1502
rect 1324 296 1959 348
rect 1324 262 1353 296
rect 1387 262 1421 296
rect 1455 262 1489 296
rect 1523 262 1557 296
rect 1591 262 1625 296
rect 1659 262 1693 296
rect 1727 262 1761 296
rect 1795 262 1829 296
rect 1863 262 1897 296
rect 1931 262 1959 296
rect 1324 220 1959 262
rect 3704 307 4244 360
rect 3704 273 3753 307
rect 3787 273 3821 307
rect 3855 273 3889 307
rect 3923 273 3957 307
rect 3991 273 4025 307
rect 4059 273 4093 307
rect 4127 273 4161 307
rect 4195 273 4244 307
rect 3704 220 4244 273
<< mvnsubdiff >>
rect 1348 4682 1880 4734
rect 1348 4648 1395 4682
rect 1429 4648 1463 4682
rect 1497 4648 1531 4682
rect 1565 4648 1599 4682
rect 1633 4648 1667 4682
rect 1701 4648 1735 4682
rect 1769 4648 1803 4682
rect 1837 4648 1880 4682
rect 1348 4594 1880 4648
rect 3734 4681 4254 4724
rect 3734 4647 3773 4681
rect 3807 4647 3841 4681
rect 3875 4647 3909 4681
rect 3943 4647 3977 4681
rect 4011 4647 4045 4681
rect 4079 4647 4113 4681
rect 4147 4647 4181 4681
rect 4215 4647 4254 4681
rect 3734 4604 4254 4647
rect 5692 4680 6212 4724
rect 5692 4646 5732 4680
rect 5766 4646 5800 4680
rect 5834 4646 5868 4680
rect 5902 4646 5936 4680
rect 5970 4646 6004 4680
rect 6038 4646 6072 4680
rect 6106 4646 6140 4680
rect 6174 4646 6212 4680
rect 5692 4604 6212 4646
rect 1348 3454 1880 3506
rect 1348 3420 1395 3454
rect 1429 3420 1463 3454
rect 1497 3420 1531 3454
rect 1565 3420 1599 3454
rect 1633 3420 1667 3454
rect 1701 3420 1735 3454
rect 1769 3420 1803 3454
rect 1837 3420 1880 3454
rect 1348 3366 1880 3420
rect 3734 3453 4254 3496
rect 3734 3419 3773 3453
rect 3807 3419 3841 3453
rect 3875 3419 3909 3453
rect 3943 3419 3977 3453
rect 4011 3419 4045 3453
rect 4079 3419 4113 3453
rect 4147 3419 4181 3453
rect 4215 3419 4254 3453
rect 3734 3376 4254 3419
rect 5692 3452 6212 3496
rect 5692 3418 5732 3452
rect 5766 3418 5800 3452
rect 5834 3418 5868 3452
rect 5902 3418 5936 3452
rect 5970 3418 6004 3452
rect 6038 3418 6072 3452
rect 6106 3418 6140 3452
rect 6174 3418 6212 3452
rect 5692 3376 6212 3418
rect 1348 2226 1880 2278
rect 1348 2192 1395 2226
rect 1429 2192 1463 2226
rect 1497 2192 1531 2226
rect 1565 2192 1599 2226
rect 1633 2192 1667 2226
rect 1701 2192 1735 2226
rect 1769 2192 1803 2226
rect 1837 2192 1880 2226
rect 1348 2138 1880 2192
rect 3734 2225 4254 2268
rect 3734 2191 3773 2225
rect 3807 2191 3841 2225
rect 3875 2191 3909 2225
rect 3943 2191 3977 2225
rect 4011 2191 4045 2225
rect 4079 2191 4113 2225
rect 4147 2191 4181 2225
rect 4215 2191 4254 2225
rect 3734 2148 4254 2191
rect 5692 2224 6212 2268
rect 5692 2190 5732 2224
rect 5766 2190 5800 2224
rect 5834 2190 5868 2224
rect 5902 2190 5936 2224
rect 5970 2190 6004 2224
rect 6038 2190 6072 2224
rect 6106 2190 6140 2224
rect 6174 2190 6212 2224
rect 5692 2148 6212 2190
rect 1348 998 1880 1050
rect 1348 964 1395 998
rect 1429 964 1463 998
rect 1497 964 1531 998
rect 1565 964 1599 998
rect 1633 964 1667 998
rect 1701 964 1735 998
rect 1769 964 1803 998
rect 1837 964 1880 998
rect 1348 910 1880 964
rect 3734 997 4254 1040
rect 3734 963 3773 997
rect 3807 963 3841 997
rect 3875 963 3909 997
rect 3943 963 3977 997
rect 4011 963 4045 997
rect 4079 963 4113 997
rect 4147 963 4181 997
rect 4215 963 4254 997
rect 3734 920 4254 963
<< psubdiffcont >>
rect 1353 3946 1387 3980
rect 1421 3946 1455 3980
rect 1489 3946 1523 3980
rect 1557 3946 1591 3980
rect 1625 3946 1659 3980
rect 1693 3946 1727 3980
rect 1761 3946 1795 3980
rect 1829 3946 1863 3980
rect 1897 3946 1931 3980
rect 3753 3957 3787 3991
rect 3821 3957 3855 3991
rect 3889 3957 3923 3991
rect 3957 3957 3991 3991
rect 4025 3957 4059 3991
rect 4093 3957 4127 3991
rect 4161 3957 4195 3991
rect 5712 3958 5746 3992
rect 5780 3958 5814 3992
rect 5848 3958 5882 3992
rect 5916 3958 5950 3992
rect 5984 3958 6018 3992
rect 6052 3958 6086 3992
rect 6120 3958 6154 3992
rect 1353 2718 1387 2752
rect 1421 2718 1455 2752
rect 1489 2718 1523 2752
rect 1557 2718 1591 2752
rect 1625 2718 1659 2752
rect 1693 2718 1727 2752
rect 1761 2718 1795 2752
rect 1829 2718 1863 2752
rect 1897 2718 1931 2752
rect 3753 2729 3787 2763
rect 3821 2729 3855 2763
rect 3889 2729 3923 2763
rect 3957 2729 3991 2763
rect 4025 2729 4059 2763
rect 4093 2729 4127 2763
rect 4161 2729 4195 2763
rect 5712 2730 5746 2764
rect 5780 2730 5814 2764
rect 5848 2730 5882 2764
rect 5916 2730 5950 2764
rect 5984 2730 6018 2764
rect 6052 2730 6086 2764
rect 6120 2730 6154 2764
rect 1353 1490 1387 1524
rect 1421 1490 1455 1524
rect 1489 1490 1523 1524
rect 1557 1490 1591 1524
rect 1625 1490 1659 1524
rect 1693 1490 1727 1524
rect 1761 1490 1795 1524
rect 1829 1490 1863 1524
rect 1897 1490 1931 1524
rect 3753 1501 3787 1535
rect 3821 1501 3855 1535
rect 3889 1501 3923 1535
rect 3957 1501 3991 1535
rect 4025 1501 4059 1535
rect 4093 1501 4127 1535
rect 4161 1501 4195 1535
rect 5712 1502 5746 1536
rect 5780 1502 5814 1536
rect 5848 1502 5882 1536
rect 5916 1502 5950 1536
rect 5984 1502 6018 1536
rect 6052 1502 6086 1536
rect 6120 1502 6154 1536
rect 1353 262 1387 296
rect 1421 262 1455 296
rect 1489 262 1523 296
rect 1557 262 1591 296
rect 1625 262 1659 296
rect 1693 262 1727 296
rect 1761 262 1795 296
rect 1829 262 1863 296
rect 1897 262 1931 296
rect 3753 273 3787 307
rect 3821 273 3855 307
rect 3889 273 3923 307
rect 3957 273 3991 307
rect 4025 273 4059 307
rect 4093 273 4127 307
rect 4161 273 4195 307
<< mvnsubdiffcont >>
rect 1395 4648 1429 4682
rect 1463 4648 1497 4682
rect 1531 4648 1565 4682
rect 1599 4648 1633 4682
rect 1667 4648 1701 4682
rect 1735 4648 1769 4682
rect 1803 4648 1837 4682
rect 3773 4647 3807 4681
rect 3841 4647 3875 4681
rect 3909 4647 3943 4681
rect 3977 4647 4011 4681
rect 4045 4647 4079 4681
rect 4113 4647 4147 4681
rect 4181 4647 4215 4681
rect 5732 4646 5766 4680
rect 5800 4646 5834 4680
rect 5868 4646 5902 4680
rect 5936 4646 5970 4680
rect 6004 4646 6038 4680
rect 6072 4646 6106 4680
rect 6140 4646 6174 4680
rect 1395 3420 1429 3454
rect 1463 3420 1497 3454
rect 1531 3420 1565 3454
rect 1599 3420 1633 3454
rect 1667 3420 1701 3454
rect 1735 3420 1769 3454
rect 1803 3420 1837 3454
rect 3773 3419 3807 3453
rect 3841 3419 3875 3453
rect 3909 3419 3943 3453
rect 3977 3419 4011 3453
rect 4045 3419 4079 3453
rect 4113 3419 4147 3453
rect 4181 3419 4215 3453
rect 5732 3418 5766 3452
rect 5800 3418 5834 3452
rect 5868 3418 5902 3452
rect 5936 3418 5970 3452
rect 6004 3418 6038 3452
rect 6072 3418 6106 3452
rect 6140 3418 6174 3452
rect 1395 2192 1429 2226
rect 1463 2192 1497 2226
rect 1531 2192 1565 2226
rect 1599 2192 1633 2226
rect 1667 2192 1701 2226
rect 1735 2192 1769 2226
rect 1803 2192 1837 2226
rect 3773 2191 3807 2225
rect 3841 2191 3875 2225
rect 3909 2191 3943 2225
rect 3977 2191 4011 2225
rect 4045 2191 4079 2225
rect 4113 2191 4147 2225
rect 4181 2191 4215 2225
rect 5732 2190 5766 2224
rect 5800 2190 5834 2224
rect 5868 2190 5902 2224
rect 5936 2190 5970 2224
rect 6004 2190 6038 2224
rect 6072 2190 6106 2224
rect 6140 2190 6174 2224
rect 1395 964 1429 998
rect 1463 964 1497 998
rect 1531 964 1565 998
rect 1599 964 1633 998
rect 1667 964 1701 998
rect 1735 964 1769 998
rect 1803 964 1837 998
rect 3773 963 3807 997
rect 3841 963 3875 997
rect 3909 963 3943 997
rect 3977 963 4011 997
rect 4045 963 4079 997
rect 4113 963 4147 997
rect 4181 963 4215 997
<< poly >>
rect 1456 4528 1556 4554
rect 1744 4528 1844 4554
rect 2076 4528 2176 4554
rect 2418 4528 2518 4554
rect 2822 4528 2922 4554
rect 3166 4528 3266 4554
rect 3788 4538 3888 4564
rect 4096 4538 4196 4564
rect 4448 4538 4548 4564
rect 4756 4538 4856 4564
rect 5746 4538 5846 4564
rect 6054 4538 6154 4564
rect 6406 4538 6506 4564
rect 6714 4538 6814 4564
rect 1456 4300 1556 4328
rect 1239 4275 1556 4300
rect 1239 4241 1269 4275
rect 1303 4241 1556 4275
rect 1239 4217 1556 4241
rect 1456 4190 1556 4217
rect 1744 4275 1844 4328
rect 1744 4241 1773 4275
rect 1807 4241 1844 4275
rect 1744 4190 1844 4241
rect 2076 4285 2176 4328
rect 2418 4306 2518 4328
rect 2621 4306 2707 4307
rect 2076 4273 2325 4285
rect 2076 4239 2273 4273
rect 2307 4239 2325 4273
rect 2076 4227 2325 4239
rect 2418 4283 2712 4306
rect 2418 4249 2647 4283
rect 2681 4249 2712 4283
rect 2076 4190 2176 4227
rect 2418 4215 2712 4249
rect 2822 4271 2922 4328
rect 2822 4237 2857 4271
rect 2891 4237 2922 4271
rect 2418 4190 2518 4215
rect 2822 4190 2922 4237
rect 3019 4281 3073 4287
rect 3166 4281 3266 4328
rect 3019 4271 3266 4281
rect 3019 4237 3029 4271
rect 3063 4237 3266 4271
rect 3654 4297 3720 4305
rect 3788 4297 3888 4338
rect 3654 4295 3888 4297
rect 3654 4261 3670 4295
rect 3704 4261 3888 4295
rect 3654 4258 3888 4261
rect 3654 4251 3720 4258
rect 3019 4227 3266 4237
rect 3019 4221 3073 4227
rect 3166 4190 3266 4227
rect 3788 4200 3888 4258
rect 3968 4288 4034 4296
rect 4096 4288 4196 4338
rect 3968 4286 4196 4288
rect 3968 4252 3984 4286
rect 4018 4252 4196 4286
rect 3968 4249 4196 4252
rect 3968 4242 4034 4249
rect 4096 4200 4196 4249
rect 4290 4280 4356 4290
rect 4448 4280 4548 4338
rect 4290 4246 4306 4280
rect 4340 4246 4548 4280
rect 4627 4298 4681 4314
rect 4627 4264 4637 4298
rect 4671 4296 4681 4298
rect 4756 4296 4856 4338
rect 4671 4265 4856 4296
rect 4671 4264 4681 4265
rect 4627 4248 4681 4264
rect 4290 4245 4548 4246
rect 4290 4236 4356 4245
rect 4448 4202 4548 4245
rect 4756 4202 4856 4265
rect 5612 4298 5678 4306
rect 5746 4298 5846 4338
rect 5612 4296 5846 4298
rect 5612 4262 5628 4296
rect 5662 4262 5846 4296
rect 5612 4258 5846 4262
rect 5612 4252 5678 4258
rect 5746 4200 5846 4258
rect 5926 4288 5992 4296
rect 6054 4288 6154 4338
rect 5926 4286 6154 4288
rect 5926 4252 5942 4286
rect 5976 4252 6154 4286
rect 5926 4250 6154 4252
rect 5926 4242 5992 4250
rect 6054 4200 6154 4250
rect 6248 4280 6314 4290
rect 6406 4280 6506 4338
rect 6248 4246 6264 4280
rect 6298 4246 6506 4280
rect 6586 4298 6640 4314
rect 6586 4264 6596 4298
rect 6630 4296 6640 4298
rect 6714 4296 6814 4338
rect 6630 4266 6814 4296
rect 6630 4264 6640 4266
rect 6586 4248 6640 4264
rect 6248 4236 6314 4246
rect 6406 4202 6506 4246
rect 6714 4202 6814 4266
rect 1456 4064 1556 4090
rect 1744 4064 1844 4090
rect 2076 4064 2176 4090
rect 2418 4064 2518 4090
rect 2822 4064 2922 4090
rect 3166 4064 3266 4090
rect 3788 4074 3888 4100
rect 4096 4074 4196 4100
rect 4448 4076 4548 4102
rect 4756 4076 4856 4102
rect 5746 4074 5846 4100
rect 6054 4074 6154 4100
rect 6406 4076 6506 4102
rect 6714 4076 6814 4102
rect 1456 3300 1556 3326
rect 1744 3300 1844 3326
rect 2076 3300 2176 3326
rect 2418 3300 2518 3326
rect 2822 3300 2922 3326
rect 3166 3300 3266 3326
rect 3788 3310 3888 3336
rect 4096 3310 4196 3336
rect 4448 3310 4548 3336
rect 4756 3310 4856 3336
rect 5746 3310 5846 3336
rect 6054 3310 6154 3336
rect 6406 3310 6506 3336
rect 6714 3310 6814 3336
rect 1456 3072 1556 3100
rect 1239 3047 1556 3072
rect 1239 3013 1269 3047
rect 1303 3013 1556 3047
rect 1239 2989 1556 3013
rect 1456 2962 1556 2989
rect 1744 3047 1844 3100
rect 1744 3013 1773 3047
rect 1807 3013 1844 3047
rect 1744 2962 1844 3013
rect 2076 3057 2176 3100
rect 2418 3078 2518 3100
rect 2621 3078 2707 3079
rect 2076 3045 2325 3057
rect 2076 3011 2273 3045
rect 2307 3011 2325 3045
rect 2076 2999 2325 3011
rect 2418 3055 2712 3078
rect 2418 3021 2647 3055
rect 2681 3021 2712 3055
rect 2076 2962 2176 2999
rect 2418 2987 2712 3021
rect 2822 3043 2922 3100
rect 2822 3009 2857 3043
rect 2891 3009 2922 3043
rect 2418 2962 2518 2987
rect 2822 2962 2922 3009
rect 3019 3053 3073 3059
rect 3166 3053 3266 3100
rect 3019 3043 3266 3053
rect 3019 3009 3029 3043
rect 3063 3009 3266 3043
rect 3654 3069 3720 3077
rect 3788 3069 3888 3110
rect 3654 3067 3888 3069
rect 3654 3033 3670 3067
rect 3704 3033 3888 3067
rect 3654 3030 3888 3033
rect 3654 3023 3720 3030
rect 3019 2999 3266 3009
rect 3019 2993 3073 2999
rect 3166 2962 3266 2999
rect 3788 2972 3888 3030
rect 3968 3060 4034 3068
rect 4096 3060 4196 3110
rect 3968 3058 4196 3060
rect 3968 3024 3984 3058
rect 4018 3024 4196 3058
rect 3968 3021 4196 3024
rect 3968 3014 4034 3021
rect 4096 2972 4196 3021
rect 4290 3052 4356 3062
rect 4448 3052 4548 3110
rect 4290 3018 4306 3052
rect 4340 3018 4548 3052
rect 4627 3070 4681 3086
rect 4627 3036 4637 3070
rect 4671 3068 4681 3070
rect 4756 3068 4856 3110
rect 4671 3037 4856 3068
rect 4671 3036 4681 3037
rect 4627 3020 4681 3036
rect 4290 3017 4548 3018
rect 4290 3008 4356 3017
rect 4448 2974 4548 3017
rect 4756 2974 4856 3037
rect 5612 3070 5678 3078
rect 5746 3070 5846 3110
rect 5612 3068 5846 3070
rect 5612 3034 5628 3068
rect 5662 3034 5846 3068
rect 5612 3030 5846 3034
rect 5612 3024 5678 3030
rect 5746 2972 5846 3030
rect 5926 3060 5992 3068
rect 6054 3060 6154 3110
rect 5926 3058 6154 3060
rect 5926 3024 5942 3058
rect 5976 3024 6154 3058
rect 5926 3022 6154 3024
rect 5926 3014 5992 3022
rect 6054 2972 6154 3022
rect 6248 3052 6314 3062
rect 6406 3052 6506 3110
rect 6248 3018 6264 3052
rect 6298 3018 6506 3052
rect 6586 3070 6640 3086
rect 6586 3036 6596 3070
rect 6630 3068 6640 3070
rect 6714 3068 6814 3110
rect 6630 3038 6814 3068
rect 6630 3036 6640 3038
rect 6586 3020 6640 3036
rect 6248 3008 6314 3018
rect 6406 2974 6506 3018
rect 6714 2974 6814 3038
rect 1456 2836 1556 2862
rect 1744 2836 1844 2862
rect 2076 2836 2176 2862
rect 2418 2836 2518 2862
rect 2822 2836 2922 2862
rect 3166 2836 3266 2862
rect 3788 2846 3888 2872
rect 4096 2846 4196 2872
rect 4448 2848 4548 2874
rect 4756 2848 4856 2874
rect 5746 2846 5846 2872
rect 6054 2846 6154 2872
rect 6406 2848 6506 2874
rect 6714 2848 6814 2874
rect 1456 2072 1556 2098
rect 1744 2072 1844 2098
rect 2076 2072 2176 2098
rect 2418 2072 2518 2098
rect 2822 2072 2922 2098
rect 3166 2072 3266 2098
rect 3788 2082 3888 2108
rect 4096 2082 4196 2108
rect 4448 2082 4548 2108
rect 4756 2082 4856 2108
rect 5746 2082 5846 2108
rect 6054 2082 6154 2108
rect 6406 2082 6506 2108
rect 6714 2082 6814 2108
rect 1456 1844 1556 1872
rect 1239 1819 1556 1844
rect 1239 1785 1269 1819
rect 1303 1785 1556 1819
rect 1239 1761 1556 1785
rect 1456 1734 1556 1761
rect 1744 1819 1844 1872
rect 1744 1785 1773 1819
rect 1807 1785 1844 1819
rect 1744 1734 1844 1785
rect 2076 1829 2176 1872
rect 2418 1850 2518 1872
rect 2621 1850 2707 1851
rect 2076 1817 2325 1829
rect 2076 1783 2273 1817
rect 2307 1783 2325 1817
rect 2076 1771 2325 1783
rect 2418 1827 2712 1850
rect 2418 1793 2647 1827
rect 2681 1793 2712 1827
rect 2076 1734 2176 1771
rect 2418 1759 2712 1793
rect 2822 1815 2922 1872
rect 2822 1781 2857 1815
rect 2891 1781 2922 1815
rect 2418 1734 2518 1759
rect 2822 1734 2922 1781
rect 3019 1825 3073 1831
rect 3166 1825 3266 1872
rect 3019 1815 3266 1825
rect 3019 1781 3029 1815
rect 3063 1781 3266 1815
rect 3654 1841 3720 1849
rect 3788 1841 3888 1882
rect 3654 1839 3888 1841
rect 3654 1805 3670 1839
rect 3704 1805 3888 1839
rect 3654 1802 3888 1805
rect 3654 1795 3720 1802
rect 3019 1771 3266 1781
rect 3019 1765 3073 1771
rect 3166 1734 3266 1771
rect 3788 1744 3888 1802
rect 3968 1832 4034 1840
rect 4096 1832 4196 1882
rect 3968 1830 4196 1832
rect 3968 1796 3984 1830
rect 4018 1796 4196 1830
rect 3968 1793 4196 1796
rect 3968 1786 4034 1793
rect 4096 1744 4196 1793
rect 4290 1824 4356 1834
rect 4448 1824 4548 1882
rect 4290 1790 4306 1824
rect 4340 1790 4548 1824
rect 4627 1842 4681 1858
rect 4627 1808 4637 1842
rect 4671 1840 4681 1842
rect 4756 1840 4856 1882
rect 4671 1809 4856 1840
rect 4671 1808 4681 1809
rect 4627 1792 4681 1808
rect 4290 1789 4548 1790
rect 4290 1780 4356 1789
rect 4448 1746 4548 1789
rect 4756 1746 4856 1809
rect 5612 1842 5678 1850
rect 5746 1842 5846 1882
rect 5612 1840 5846 1842
rect 5612 1806 5628 1840
rect 5662 1806 5846 1840
rect 5612 1802 5846 1806
rect 5612 1796 5678 1802
rect 5746 1744 5846 1802
rect 5926 1832 5992 1840
rect 6054 1832 6154 1882
rect 5926 1830 6154 1832
rect 5926 1796 5942 1830
rect 5976 1796 6154 1830
rect 5926 1794 6154 1796
rect 5926 1786 5992 1794
rect 6054 1744 6154 1794
rect 6248 1824 6314 1834
rect 6406 1824 6506 1882
rect 6248 1790 6264 1824
rect 6298 1790 6506 1824
rect 6586 1842 6640 1858
rect 6586 1808 6596 1842
rect 6630 1840 6640 1842
rect 6714 1840 6814 1882
rect 6630 1810 6814 1840
rect 6630 1808 6640 1810
rect 6586 1792 6640 1808
rect 6248 1780 6314 1790
rect 6406 1746 6506 1790
rect 6714 1746 6814 1810
rect 1456 1608 1556 1634
rect 1744 1608 1844 1634
rect 2076 1608 2176 1634
rect 2418 1608 2518 1634
rect 2822 1608 2922 1634
rect 3166 1608 3266 1634
rect 3788 1618 3888 1644
rect 4096 1618 4196 1644
rect 4448 1620 4548 1646
rect 4756 1620 4856 1646
rect 5746 1618 5846 1644
rect 6054 1618 6154 1644
rect 6406 1620 6506 1646
rect 6714 1620 6814 1646
rect 1456 844 1556 870
rect 1744 844 1844 870
rect 2076 844 2176 870
rect 2418 844 2518 870
rect 2822 844 2922 870
rect 3166 844 3266 870
rect 3788 854 3888 880
rect 4096 854 4196 880
rect 4448 854 4548 880
rect 4756 854 4856 880
rect 1456 616 1556 644
rect 1239 591 1556 616
rect 1239 557 1269 591
rect 1303 557 1556 591
rect 1239 533 1556 557
rect 1456 506 1556 533
rect 1744 591 1844 644
rect 1744 557 1773 591
rect 1807 557 1844 591
rect 1744 506 1844 557
rect 2076 601 2176 644
rect 2418 622 2518 644
rect 2621 622 2707 623
rect 2076 589 2325 601
rect 2076 555 2273 589
rect 2307 555 2325 589
rect 2076 543 2325 555
rect 2418 599 2712 622
rect 2418 565 2647 599
rect 2681 565 2712 599
rect 2076 506 2176 543
rect 2418 531 2712 565
rect 2822 587 2922 644
rect 2822 553 2857 587
rect 2891 553 2922 587
rect 2418 506 2518 531
rect 2822 506 2922 553
rect 3019 597 3073 603
rect 3166 597 3266 644
rect 3019 587 3266 597
rect 3019 553 3029 587
rect 3063 553 3266 587
rect 3654 613 3720 621
rect 3788 613 3888 654
rect 3654 611 3888 613
rect 3654 577 3670 611
rect 3704 577 3888 611
rect 3654 574 3888 577
rect 3654 567 3720 574
rect 3019 543 3266 553
rect 3019 537 3073 543
rect 3166 506 3266 543
rect 3788 516 3888 574
rect 3968 604 4034 612
rect 4096 604 4196 654
rect 3968 602 4196 604
rect 3968 568 3984 602
rect 4018 568 4196 602
rect 3968 565 4196 568
rect 3968 558 4034 565
rect 4096 516 4196 565
rect 4290 596 4356 606
rect 4448 596 4548 654
rect 4290 562 4306 596
rect 4340 562 4548 596
rect 4627 614 4681 630
rect 4627 580 4637 614
rect 4671 612 4681 614
rect 4756 612 4856 654
rect 4671 581 4856 612
rect 4671 580 4681 581
rect 4627 564 4681 580
rect 4290 561 4548 562
rect 4290 552 4356 561
rect 4448 518 4548 561
rect 4756 518 4856 581
rect 1456 380 1556 406
rect 1744 380 1844 406
rect 2076 380 2176 406
rect 2418 380 2518 406
rect 2822 380 2922 406
rect 3166 380 3266 406
rect 3788 390 3888 416
rect 4096 390 4196 416
rect 4448 392 4548 418
rect 4756 392 4856 418
<< polycont >>
rect 1269 4241 1303 4275
rect 1773 4241 1807 4275
rect 2273 4239 2307 4273
rect 2647 4249 2681 4283
rect 2857 4237 2891 4271
rect 3029 4237 3063 4271
rect 3670 4261 3704 4295
rect 3984 4252 4018 4286
rect 4306 4246 4340 4280
rect 4637 4264 4671 4298
rect 5628 4262 5662 4296
rect 5942 4252 5976 4286
rect 6264 4246 6298 4280
rect 6596 4264 6630 4298
rect 1269 3013 1303 3047
rect 1773 3013 1807 3047
rect 2273 3011 2307 3045
rect 2647 3021 2681 3055
rect 2857 3009 2891 3043
rect 3029 3009 3063 3043
rect 3670 3033 3704 3067
rect 3984 3024 4018 3058
rect 4306 3018 4340 3052
rect 4637 3036 4671 3070
rect 5628 3034 5662 3068
rect 5942 3024 5976 3058
rect 6264 3018 6298 3052
rect 6596 3036 6630 3070
rect 1269 1785 1303 1819
rect 1773 1785 1807 1819
rect 2273 1783 2307 1817
rect 2647 1793 2681 1827
rect 2857 1781 2891 1815
rect 3029 1781 3063 1815
rect 3670 1805 3704 1839
rect 3984 1796 4018 1830
rect 4306 1790 4340 1824
rect 4637 1808 4671 1842
rect 5628 1806 5662 1840
rect 5942 1796 5976 1830
rect 6264 1790 6298 1824
rect 6596 1808 6630 1842
rect 1269 557 1303 591
rect 1773 557 1807 591
rect 2273 555 2307 589
rect 2647 565 2681 599
rect 2857 553 2891 587
rect 3029 553 3063 587
rect 3670 577 3704 611
rect 3984 568 4018 602
rect 4306 562 4340 596
rect 4637 580 4671 614
<< mvndiffres >>
rect 544 4101 628 4521
rect 690 4101 774 4521
rect 834 4107 918 4527
rect 988 4107 1072 4527
rect 544 2873 628 3293
rect 690 2873 774 3293
rect 834 2879 918 3299
rect 988 2879 1072 3299
rect 544 1645 628 2065
rect 690 1645 774 2065
rect 834 1651 918 2071
rect 988 1651 1072 2071
rect 544 417 628 837
rect 690 417 774 837
rect 834 423 918 843
rect 988 423 1072 843
<< locali >>
rect 1348 4682 1880 4734
rect 1348 4648 1383 4682
rect 1429 4648 1455 4682
rect 1497 4648 1527 4682
rect 1565 4648 1599 4682
rect 1633 4648 1667 4682
rect 1705 4648 1735 4682
rect 1777 4648 1803 4682
rect 1849 4648 1880 4682
rect 3724 4681 4264 4734
rect 540 4596 569 4612
rect 603 4596 632 4612
rect 540 4578 566 4596
rect 607 4578 632 4596
rect 686 4596 715 4612
rect 749 4596 778 4612
rect 686 4578 710 4596
rect 751 4578 778 4596
rect 830 4601 859 4618
rect 893 4601 922 4618
rect 830 4584 856 4601
rect 897 4584 922 4601
rect 984 4601 1013 4618
rect 1047 4601 1076 4618
rect 984 4584 1009 4601
rect 1050 4584 1076 4601
rect 1348 4594 1880 4648
rect 2627 4601 3073 4655
rect 556 4556 566 4578
rect 607 4556 616 4578
rect 556 4538 616 4556
rect 702 4556 710 4578
rect 751 4556 762 4578
rect 702 4538 762 4556
rect 846 4561 856 4584
rect 897 4561 906 4584
rect 846 4544 906 4561
rect 1000 4561 1009 4584
rect 1050 4561 1060 4584
rect 1000 4544 1060 4561
rect 1410 4513 1444 4532
rect 1410 4445 1444 4447
rect 1410 4409 1444 4411
rect 1410 4324 1444 4343
rect 1568 4513 1602 4532
rect 1568 4445 1602 4447
rect 1568 4409 1602 4411
rect 1568 4324 1602 4343
rect 1698 4513 1732 4532
rect 1698 4445 1732 4447
rect 1698 4409 1732 4411
rect 1698 4324 1732 4343
rect 1856 4513 1890 4532
rect 1856 4445 1890 4447
rect 1856 4409 1890 4411
rect 1856 4324 1890 4343
rect 2030 4513 2064 4532
rect 2030 4445 2064 4447
rect 2030 4409 2064 4411
rect 2030 4324 2064 4343
rect 2188 4513 2222 4532
rect 2188 4445 2222 4447
rect 2188 4409 2222 4411
rect 2188 4324 2222 4343
rect 2372 4513 2406 4532
rect 2372 4445 2406 4447
rect 2372 4409 2406 4411
rect 2372 4324 2406 4343
rect 2530 4513 2564 4532
rect 2627 4451 2681 4601
rect 2776 4513 2810 4532
rect 2530 4445 2564 4447
rect 2530 4409 2564 4411
rect 2530 4324 2564 4343
rect 2625 4429 2703 4451
rect 2625 4395 2647 4429
rect 2681 4395 2703 4429
rect 1255 4294 1318 4306
rect 1251 4275 1322 4294
rect 2625 4291 2703 4395
rect 2776 4445 2810 4447
rect 2776 4409 2810 4411
rect 2776 4324 2810 4343
rect 2934 4513 2968 4532
rect 2934 4445 2968 4447
rect 2934 4409 2968 4411
rect 2934 4324 2968 4343
rect 1773 4282 1807 4291
rect 2271 4285 2309 4291
rect 1251 4241 1269 4275
rect 1303 4241 1322 4275
rect 1251 4223 1322 4241
rect 1766 4275 1814 4282
rect 1766 4241 1773 4275
rect 1807 4241 1814 4275
rect 1766 4234 1814 4241
rect 2261 4273 2319 4285
rect 2261 4239 2273 4273
rect 2307 4239 2319 4273
rect 2615 4283 2713 4291
rect 2615 4249 2647 4283
rect 2681 4249 2713 4283
rect 2857 4278 2891 4287
rect 2615 4242 2713 4249
rect 2850 4271 2898 4278
rect 3019 4271 3073 4601
rect 3724 4647 3773 4681
rect 3831 4647 3841 4681
rect 3903 4647 3909 4681
rect 3975 4647 3977 4681
rect 4011 4647 4013 4681
rect 4079 4647 4085 4681
rect 4147 4647 4157 4681
rect 4215 4647 4264 4681
rect 3724 4594 4264 4647
rect 5682 4680 6222 4734
rect 5682 4646 5732 4680
rect 5790 4646 5800 4680
rect 5862 4646 5868 4680
rect 5934 4646 5936 4680
rect 5970 4646 5972 4680
rect 6038 4646 6044 4680
rect 6106 4646 6116 4680
rect 6174 4646 6222 4680
rect 5682 4594 6222 4646
rect 3120 4513 3154 4532
rect 3120 4445 3154 4447
rect 3120 4409 3154 4411
rect 3120 4324 3154 4343
rect 3278 4513 3312 4532
rect 3278 4445 3312 4447
rect 3278 4409 3312 4411
rect 3278 4324 3312 4343
rect 3742 4523 3776 4542
rect 3742 4455 3776 4457
rect 3742 4419 3776 4421
rect 3742 4334 3776 4353
rect 3900 4523 3934 4542
rect 3900 4455 3934 4457
rect 3900 4419 3934 4421
rect 3900 4334 3934 4353
rect 4050 4523 4084 4542
rect 4050 4455 4084 4457
rect 4050 4419 4084 4421
rect 4050 4334 4084 4353
rect 4208 4523 4242 4542
rect 4208 4455 4242 4457
rect 4208 4419 4242 4421
rect 4208 4334 4242 4353
rect 4402 4523 4436 4542
rect 4402 4455 4436 4457
rect 4402 4419 4436 4421
rect 4402 4334 4436 4353
rect 4560 4523 4594 4542
rect 4560 4455 4594 4457
rect 4560 4419 4594 4421
rect 4560 4334 4594 4353
rect 4710 4523 4744 4542
rect 4710 4455 4744 4457
rect 4710 4419 4744 4421
rect 4710 4334 4744 4353
rect 4868 4523 4902 4542
rect 4868 4455 4902 4457
rect 4868 4419 4902 4421
rect 4868 4334 4902 4353
rect 5700 4524 5734 4542
rect 5700 4456 5734 4458
rect 5700 4420 5734 4422
rect 5700 4334 5734 4354
rect 5858 4524 5892 4542
rect 5858 4456 5892 4458
rect 5858 4420 5892 4422
rect 5858 4334 5892 4354
rect 6008 4524 6042 4542
rect 6008 4456 6042 4458
rect 6008 4420 6042 4422
rect 6008 4334 6042 4354
rect 6166 4524 6200 4542
rect 6166 4456 6200 4458
rect 6166 4420 6200 4422
rect 6166 4334 6200 4354
rect 6360 4524 6394 4542
rect 6360 4456 6394 4458
rect 6360 4420 6394 4422
rect 6360 4334 6394 4354
rect 6518 4524 6552 4542
rect 6518 4456 6552 4458
rect 6518 4420 6552 4422
rect 6518 4334 6552 4354
rect 6668 4524 6702 4542
rect 6668 4456 6702 4458
rect 6668 4420 6702 4422
rect 6668 4334 6702 4354
rect 6826 4524 6860 4542
rect 6826 4456 6860 4458
rect 6826 4420 6860 4422
rect 6826 4334 6860 4354
rect 3670 4298 3704 4311
rect 3668 4295 3707 4298
rect 1773 4225 1807 4234
rect 2261 4227 2319 4239
rect 2625 4228 2703 4242
rect 2850 4237 2857 4271
rect 2891 4237 2898 4271
rect 3013 4237 3029 4271
rect 3063 4237 3079 4271
rect 3668 4261 3670 4295
rect 3704 4261 3707 4295
rect 3984 4289 4018 4302
rect 5628 4298 5662 4312
rect 3668 4259 3707 4261
rect 3982 4286 4021 4289
rect 3670 4245 3704 4259
rect 3982 4252 3984 4286
rect 4018 4252 4021 4286
rect 3982 4250 4021 4252
rect 4306 4281 4340 4296
rect 4306 4280 4341 4281
rect 2850 4230 2898 4237
rect 1255 4211 1318 4223
rect 2271 4221 2309 4227
rect 1410 4157 1444 4194
rect 556 4068 616 4084
rect 556 4044 565 4068
rect 606 4044 616 4068
rect 702 4068 762 4084
rect 702 4044 712 4068
rect 753 4044 762 4068
rect 846 4073 906 4090
rect 846 4050 856 4073
rect 897 4050 906 4073
rect 1000 4074 1060 4090
rect 1410 4086 1444 4123
rect 1568 4157 1602 4194
rect 1568 4086 1602 4123
rect 1698 4157 1732 4194
rect 1698 4086 1732 4123
rect 1856 4157 1890 4194
rect 1856 4086 1890 4123
rect 2030 4157 2064 4194
rect 2030 4086 2064 4123
rect 2188 4157 2222 4194
rect 2188 4086 2222 4123
rect 2352 4157 2420 4200
rect 2352 4123 2372 4157
rect 2406 4123 2420 4157
rect 1000 4050 1010 4074
rect 1051 4050 1060 4074
rect 540 4028 565 4044
rect 606 4028 632 4044
rect 540 4010 569 4028
rect 603 4010 632 4028
rect 686 4028 712 4044
rect 753 4028 778 4044
rect 686 4010 715 4028
rect 749 4010 778 4028
rect 830 4033 856 4050
rect 897 4033 922 4050
rect 830 4016 859 4033
rect 893 4016 922 4033
rect 984 4034 1010 4050
rect 1051 4034 1076 4050
rect 984 4016 1013 4034
rect 1047 4016 1076 4034
rect 1324 3980 1960 4044
rect 1324 3946 1353 3980
rect 1407 3946 1421 3980
rect 1479 3946 1489 3980
rect 1551 3946 1557 3980
rect 1623 3946 1625 3980
rect 1659 3946 1661 3980
rect 1727 3946 1733 3980
rect 1795 3946 1805 3980
rect 1863 3946 1877 3980
rect 1931 3946 1960 3980
rect 1324 3904 1960 3946
rect 2352 3955 2420 4123
rect 2530 4157 2564 4194
rect 2530 4086 2564 4123
rect 2352 3921 2369 3955
rect 2403 3921 2420 3955
rect 2352 3904 2420 3921
rect 2642 3859 2696 4228
rect 2857 4221 2891 4230
rect 3019 4227 3073 4237
rect 3984 4236 4018 4250
rect 4340 4246 4341 4280
rect 4621 4264 4637 4298
rect 4671 4264 4687 4298
rect 5626 4296 5666 4298
rect 5626 4262 5628 4296
rect 5662 4262 5666 4296
rect 5942 4290 5976 4302
rect 5626 4260 5666 4262
rect 5940 4286 5980 4290
rect 5628 4246 5662 4260
rect 5940 4252 5942 4286
rect 5976 4252 5980 4286
rect 5940 4250 5980 4252
rect 6264 4282 6298 4296
rect 6264 4280 6300 4282
rect 4306 4230 4340 4246
rect 5942 4236 5976 4250
rect 6298 4246 6300 4280
rect 6580 4264 6596 4298
rect 6630 4264 6646 4298
rect 6264 4230 6298 4246
rect 2776 4157 2810 4194
rect 2776 4086 2810 4123
rect 2934 4157 2968 4194
rect 2934 4086 2968 4123
rect 3120 4157 3154 4194
rect 3120 4086 3154 4123
rect 3278 4157 3312 4194
rect 3278 4086 3312 4123
rect 3742 4167 3776 4204
rect 3742 4096 3776 4133
rect 3900 4167 3934 4204
rect 3900 4096 3934 4133
rect 4050 4167 4084 4204
rect 4050 4096 4084 4133
rect 4208 4167 4242 4204
rect 4208 4096 4242 4133
rect 4402 4169 4436 4206
rect 4402 4098 4436 4135
rect 4560 4169 4594 4206
rect 4560 4098 4594 4135
rect 4710 4169 4744 4206
rect 4710 4098 4744 4135
rect 4868 4169 4902 4206
rect 4868 4098 4902 4135
rect 5700 4168 5734 4204
rect 5700 4096 5734 4134
rect 5858 4168 5892 4204
rect 5858 4096 5892 4134
rect 6008 4168 6042 4204
rect 6008 4096 6042 4134
rect 6166 4168 6200 4204
rect 6166 4096 6200 4134
rect 6360 4170 6394 4206
rect 6360 4098 6394 4136
rect 6518 4170 6552 4206
rect 6518 4098 6552 4136
rect 6668 4170 6702 4206
rect 6668 4098 6702 4136
rect 6826 4170 6860 4206
rect 6826 4098 6860 4136
rect 3704 3991 4244 4044
rect 3704 3957 3741 3991
rect 3787 3957 3813 3991
rect 3855 3957 3885 3991
rect 3923 3957 3957 3991
rect 3991 3957 4025 3991
rect 4063 3957 4093 3991
rect 4135 3957 4161 3991
rect 4207 3957 4244 3991
rect 3704 3904 4244 3957
rect 5662 3992 6202 4044
rect 5662 3958 5700 3992
rect 5746 3958 5772 3992
rect 5814 3958 5844 3992
rect 5882 3958 5916 3992
rect 5950 3958 5984 3992
rect 6022 3958 6052 3992
rect 6094 3958 6120 3992
rect 6166 3958 6202 3992
rect 5662 3904 6202 3958
rect 1348 3454 1880 3506
rect 1348 3420 1383 3454
rect 1429 3420 1455 3454
rect 1497 3420 1527 3454
rect 1565 3420 1599 3454
rect 1633 3420 1667 3454
rect 1705 3420 1735 3454
rect 1777 3420 1803 3454
rect 1849 3420 1880 3454
rect 3724 3453 4264 3506
rect 540 3368 569 3384
rect 603 3368 632 3384
rect 540 3350 566 3368
rect 607 3350 632 3368
rect 686 3368 715 3384
rect 749 3368 778 3384
rect 686 3350 710 3368
rect 751 3350 778 3368
rect 830 3373 859 3390
rect 893 3373 922 3390
rect 830 3356 856 3373
rect 897 3356 922 3373
rect 984 3373 1013 3390
rect 1047 3373 1076 3390
rect 984 3356 1009 3373
rect 1050 3356 1076 3373
rect 1348 3366 1880 3420
rect 2627 3373 3073 3427
rect 556 3328 566 3350
rect 607 3328 616 3350
rect 556 3310 616 3328
rect 702 3328 710 3350
rect 751 3328 762 3350
rect 702 3310 762 3328
rect 846 3333 856 3356
rect 897 3333 906 3356
rect 846 3316 906 3333
rect 1000 3333 1009 3356
rect 1050 3333 1060 3356
rect 1000 3316 1060 3333
rect 1410 3285 1444 3304
rect 1410 3217 1444 3219
rect 1410 3181 1444 3183
rect 1410 3096 1444 3115
rect 1568 3285 1602 3304
rect 1568 3217 1602 3219
rect 1568 3181 1602 3183
rect 1568 3096 1602 3115
rect 1698 3285 1732 3304
rect 1698 3217 1732 3219
rect 1698 3181 1732 3183
rect 1698 3096 1732 3115
rect 1856 3285 1890 3304
rect 1856 3217 1890 3219
rect 1856 3181 1890 3183
rect 1856 3096 1890 3115
rect 2030 3285 2064 3304
rect 2030 3217 2064 3219
rect 2030 3181 2064 3183
rect 2030 3096 2064 3115
rect 2188 3285 2222 3304
rect 2188 3217 2222 3219
rect 2188 3181 2222 3183
rect 2188 3096 2222 3115
rect 2372 3285 2406 3304
rect 2372 3217 2406 3219
rect 2372 3181 2406 3183
rect 2372 3096 2406 3115
rect 2530 3285 2564 3304
rect 2627 3223 2681 3373
rect 2776 3285 2810 3304
rect 2530 3217 2564 3219
rect 2530 3181 2564 3183
rect 2530 3096 2564 3115
rect 2625 3201 2703 3223
rect 2625 3167 2647 3201
rect 2681 3167 2703 3201
rect 1255 3066 1318 3078
rect 1251 3047 1322 3066
rect 2625 3063 2703 3167
rect 2776 3217 2810 3219
rect 2776 3181 2810 3183
rect 2776 3096 2810 3115
rect 2934 3285 2968 3304
rect 2934 3217 2968 3219
rect 2934 3181 2968 3183
rect 2934 3096 2968 3115
rect 1773 3054 1807 3063
rect 2271 3057 2309 3063
rect 1251 3013 1269 3047
rect 1303 3013 1322 3047
rect 1251 2995 1322 3013
rect 1766 3047 1814 3054
rect 1766 3013 1773 3047
rect 1807 3013 1814 3047
rect 1766 3006 1814 3013
rect 2261 3045 2319 3057
rect 2261 3011 2273 3045
rect 2307 3011 2319 3045
rect 2615 3055 2713 3063
rect 2615 3021 2647 3055
rect 2681 3021 2713 3055
rect 2857 3050 2891 3059
rect 2615 3014 2713 3021
rect 2850 3043 2898 3050
rect 3019 3043 3073 3373
rect 3724 3419 3773 3453
rect 3831 3419 3841 3453
rect 3903 3419 3909 3453
rect 3975 3419 3977 3453
rect 4011 3419 4013 3453
rect 4079 3419 4085 3453
rect 4147 3419 4157 3453
rect 4215 3419 4264 3453
rect 3724 3366 4264 3419
rect 5682 3452 6222 3506
rect 5682 3418 5732 3452
rect 5790 3418 5800 3452
rect 5862 3418 5868 3452
rect 5934 3418 5936 3452
rect 5970 3418 5972 3452
rect 6038 3418 6044 3452
rect 6106 3418 6116 3452
rect 6174 3418 6222 3452
rect 5682 3366 6222 3418
rect 3120 3285 3154 3304
rect 3120 3217 3154 3219
rect 3120 3181 3154 3183
rect 3120 3096 3154 3115
rect 3278 3285 3312 3304
rect 3278 3217 3312 3219
rect 3278 3181 3312 3183
rect 3278 3096 3312 3115
rect 3742 3295 3776 3314
rect 3742 3227 3776 3229
rect 3742 3191 3776 3193
rect 3742 3106 3776 3125
rect 3900 3295 3934 3314
rect 3900 3227 3934 3229
rect 3900 3191 3934 3193
rect 3900 3106 3934 3125
rect 4050 3295 4084 3314
rect 4050 3227 4084 3229
rect 4050 3191 4084 3193
rect 4050 3106 4084 3125
rect 4208 3295 4242 3314
rect 4208 3227 4242 3229
rect 4208 3191 4242 3193
rect 4208 3106 4242 3125
rect 4402 3295 4436 3314
rect 4402 3227 4436 3229
rect 4402 3191 4436 3193
rect 4402 3106 4436 3125
rect 4560 3295 4594 3314
rect 4560 3227 4594 3229
rect 4560 3191 4594 3193
rect 4560 3106 4594 3125
rect 4710 3295 4744 3314
rect 4710 3227 4744 3229
rect 4710 3191 4744 3193
rect 4710 3106 4744 3125
rect 4868 3295 4902 3314
rect 4868 3227 4902 3229
rect 4868 3191 4902 3193
rect 4868 3106 4902 3125
rect 5700 3296 5734 3314
rect 5700 3228 5734 3230
rect 5700 3192 5734 3194
rect 5700 3106 5734 3126
rect 5858 3296 5892 3314
rect 5858 3228 5892 3230
rect 5858 3192 5892 3194
rect 5858 3106 5892 3126
rect 6008 3296 6042 3314
rect 6008 3228 6042 3230
rect 6008 3192 6042 3194
rect 6008 3106 6042 3126
rect 6166 3296 6200 3314
rect 6166 3228 6200 3230
rect 6166 3192 6200 3194
rect 6166 3106 6200 3126
rect 6360 3296 6394 3314
rect 6360 3228 6394 3230
rect 6360 3192 6394 3194
rect 6360 3106 6394 3126
rect 6518 3296 6552 3314
rect 6518 3228 6552 3230
rect 6518 3192 6552 3194
rect 6518 3106 6552 3126
rect 6668 3296 6702 3314
rect 6668 3228 6702 3230
rect 6668 3192 6702 3194
rect 6668 3106 6702 3126
rect 6826 3296 6860 3314
rect 6826 3228 6860 3230
rect 6826 3192 6860 3194
rect 6826 3106 6860 3126
rect 3670 3070 3704 3083
rect 3668 3067 3707 3070
rect 1773 2997 1807 3006
rect 2261 2999 2319 3011
rect 2625 3000 2703 3014
rect 2850 3009 2857 3043
rect 2891 3009 2898 3043
rect 3013 3009 3029 3043
rect 3063 3009 3079 3043
rect 3668 3033 3670 3067
rect 3704 3033 3707 3067
rect 3984 3061 4018 3074
rect 5628 3070 5662 3084
rect 3668 3031 3707 3033
rect 3982 3058 4021 3061
rect 3670 3017 3704 3031
rect 3982 3024 3984 3058
rect 4018 3024 4021 3058
rect 3982 3022 4021 3024
rect 4306 3053 4340 3068
rect 4306 3052 4341 3053
rect 2850 3002 2898 3009
rect 1255 2983 1318 2995
rect 2271 2993 2309 2999
rect 1410 2929 1444 2966
rect 556 2840 616 2856
rect 556 2816 565 2840
rect 606 2816 616 2840
rect 702 2840 762 2856
rect 702 2816 712 2840
rect 753 2816 762 2840
rect 846 2845 906 2862
rect 846 2822 856 2845
rect 897 2822 906 2845
rect 1000 2846 1060 2862
rect 1410 2858 1444 2895
rect 1568 2929 1602 2966
rect 1568 2858 1602 2895
rect 1698 2929 1732 2966
rect 1698 2858 1732 2895
rect 1856 2929 1890 2966
rect 1856 2858 1890 2895
rect 2030 2929 2064 2966
rect 2030 2858 2064 2895
rect 2188 2929 2222 2966
rect 2188 2858 2222 2895
rect 2352 2929 2420 2972
rect 2352 2895 2372 2929
rect 2406 2895 2420 2929
rect 1000 2822 1010 2846
rect 1051 2822 1060 2846
rect 540 2800 565 2816
rect 606 2800 632 2816
rect 540 2782 569 2800
rect 603 2782 632 2800
rect 686 2800 712 2816
rect 753 2800 778 2816
rect 686 2782 715 2800
rect 749 2782 778 2800
rect 830 2805 856 2822
rect 897 2805 922 2822
rect 830 2788 859 2805
rect 893 2788 922 2805
rect 984 2806 1010 2822
rect 1051 2806 1076 2822
rect 984 2788 1013 2806
rect 1047 2788 1076 2806
rect 1324 2752 1960 2816
rect 1324 2718 1353 2752
rect 1407 2718 1421 2752
rect 1479 2718 1489 2752
rect 1551 2718 1557 2752
rect 1623 2718 1625 2752
rect 1659 2718 1661 2752
rect 1727 2718 1733 2752
rect 1795 2718 1805 2752
rect 1863 2718 1877 2752
rect 1931 2718 1960 2752
rect 1324 2676 1960 2718
rect 2352 2727 2420 2895
rect 2530 2929 2564 2966
rect 2530 2858 2564 2895
rect 2352 2693 2369 2727
rect 2403 2693 2420 2727
rect 2352 2676 2420 2693
rect 2642 2631 2696 3000
rect 2857 2993 2891 3002
rect 3019 2999 3073 3009
rect 3984 3008 4018 3022
rect 4340 3018 4341 3052
rect 4621 3036 4637 3070
rect 4671 3036 4687 3070
rect 5626 3068 5666 3070
rect 5626 3034 5628 3068
rect 5662 3034 5666 3068
rect 5942 3062 5976 3074
rect 5626 3032 5666 3034
rect 5940 3058 5980 3062
rect 5628 3018 5662 3032
rect 5940 3024 5942 3058
rect 5976 3024 5980 3058
rect 5940 3022 5980 3024
rect 6264 3054 6298 3068
rect 6264 3052 6300 3054
rect 4306 3002 4340 3018
rect 5942 3008 5976 3022
rect 6298 3018 6300 3052
rect 6580 3036 6596 3070
rect 6630 3036 6646 3070
rect 6264 3002 6298 3018
rect 2776 2929 2810 2966
rect 2776 2858 2810 2895
rect 2934 2929 2968 2966
rect 2934 2858 2968 2895
rect 3120 2929 3154 2966
rect 3120 2858 3154 2895
rect 3278 2929 3312 2966
rect 3278 2858 3312 2895
rect 3742 2939 3776 2976
rect 3742 2868 3776 2905
rect 3900 2939 3934 2976
rect 3900 2868 3934 2905
rect 4050 2939 4084 2976
rect 4050 2868 4084 2905
rect 4208 2939 4242 2976
rect 4208 2868 4242 2905
rect 4402 2941 4436 2978
rect 4402 2870 4436 2907
rect 4560 2941 4594 2978
rect 4560 2870 4594 2907
rect 4710 2941 4744 2978
rect 4710 2870 4744 2907
rect 4868 2941 4902 2978
rect 4868 2870 4902 2907
rect 5700 2940 5734 2976
rect 5700 2868 5734 2906
rect 5858 2940 5892 2976
rect 5858 2868 5892 2906
rect 6008 2940 6042 2976
rect 6008 2868 6042 2906
rect 6166 2940 6200 2976
rect 6166 2868 6200 2906
rect 6360 2942 6394 2978
rect 6360 2870 6394 2908
rect 6518 2942 6552 2978
rect 6518 2870 6552 2908
rect 6668 2942 6702 2978
rect 6668 2870 6702 2908
rect 6826 2942 6860 2978
rect 6826 2870 6860 2908
rect 3704 2763 4244 2816
rect 3704 2729 3741 2763
rect 3787 2729 3813 2763
rect 3855 2729 3885 2763
rect 3923 2729 3957 2763
rect 3991 2729 4025 2763
rect 4063 2729 4093 2763
rect 4135 2729 4161 2763
rect 4207 2729 4244 2763
rect 3704 2676 4244 2729
rect 5662 2764 6202 2816
rect 5662 2730 5700 2764
rect 5746 2730 5772 2764
rect 5814 2730 5844 2764
rect 5882 2730 5916 2764
rect 5950 2730 5984 2764
rect 6022 2730 6052 2764
rect 6094 2730 6120 2764
rect 6166 2730 6202 2764
rect 5662 2676 6202 2730
rect 1348 2226 1880 2278
rect 1348 2192 1383 2226
rect 1429 2192 1455 2226
rect 1497 2192 1527 2226
rect 1565 2192 1599 2226
rect 1633 2192 1667 2226
rect 1705 2192 1735 2226
rect 1777 2192 1803 2226
rect 1849 2192 1880 2226
rect 3724 2225 4264 2278
rect 540 2140 569 2156
rect 603 2140 632 2156
rect 540 2122 566 2140
rect 607 2122 632 2140
rect 686 2140 715 2156
rect 749 2140 778 2156
rect 686 2122 710 2140
rect 751 2122 778 2140
rect 830 2145 859 2162
rect 893 2145 922 2162
rect 830 2128 856 2145
rect 897 2128 922 2145
rect 984 2145 1013 2162
rect 1047 2145 1076 2162
rect 984 2128 1009 2145
rect 1050 2128 1076 2145
rect 1348 2138 1880 2192
rect 2627 2145 3073 2199
rect 556 2100 566 2122
rect 607 2100 616 2122
rect 556 2082 616 2100
rect 702 2100 710 2122
rect 751 2100 762 2122
rect 702 2082 762 2100
rect 846 2105 856 2128
rect 897 2105 906 2128
rect 846 2088 906 2105
rect 1000 2105 1009 2128
rect 1050 2105 1060 2128
rect 1000 2088 1060 2105
rect 1410 2057 1444 2076
rect 1410 1989 1444 1991
rect 1410 1953 1444 1955
rect 1410 1868 1444 1887
rect 1568 2057 1602 2076
rect 1568 1989 1602 1991
rect 1568 1953 1602 1955
rect 1568 1868 1602 1887
rect 1698 2057 1732 2076
rect 1698 1989 1732 1991
rect 1698 1953 1732 1955
rect 1698 1868 1732 1887
rect 1856 2057 1890 2076
rect 1856 1989 1890 1991
rect 1856 1953 1890 1955
rect 1856 1868 1890 1887
rect 2030 2057 2064 2076
rect 2030 1989 2064 1991
rect 2030 1953 2064 1955
rect 2030 1868 2064 1887
rect 2188 2057 2222 2076
rect 2188 1989 2222 1991
rect 2188 1953 2222 1955
rect 2188 1868 2222 1887
rect 2372 2057 2406 2076
rect 2372 1989 2406 1991
rect 2372 1953 2406 1955
rect 2372 1868 2406 1887
rect 2530 2057 2564 2076
rect 2627 1995 2681 2145
rect 2776 2057 2810 2076
rect 2530 1989 2564 1991
rect 2530 1953 2564 1955
rect 2530 1868 2564 1887
rect 2625 1973 2703 1995
rect 2625 1939 2647 1973
rect 2681 1939 2703 1973
rect 1255 1838 1318 1850
rect 1251 1819 1322 1838
rect 2625 1835 2703 1939
rect 2776 1989 2810 1991
rect 2776 1953 2810 1955
rect 2776 1868 2810 1887
rect 2934 2057 2968 2076
rect 2934 1989 2968 1991
rect 2934 1953 2968 1955
rect 2934 1868 2968 1887
rect 1773 1826 1807 1835
rect 2271 1829 2309 1835
rect 1251 1785 1269 1819
rect 1303 1785 1322 1819
rect 1251 1767 1322 1785
rect 1766 1819 1814 1826
rect 1766 1785 1773 1819
rect 1807 1785 1814 1819
rect 1766 1778 1814 1785
rect 2261 1817 2319 1829
rect 2261 1783 2273 1817
rect 2307 1783 2319 1817
rect 2615 1827 2713 1835
rect 2615 1793 2647 1827
rect 2681 1793 2713 1827
rect 2857 1822 2891 1831
rect 2615 1786 2713 1793
rect 2850 1815 2898 1822
rect 3019 1815 3073 2145
rect 3724 2191 3773 2225
rect 3831 2191 3841 2225
rect 3903 2191 3909 2225
rect 3975 2191 3977 2225
rect 4011 2191 4013 2225
rect 4079 2191 4085 2225
rect 4147 2191 4157 2225
rect 4215 2191 4264 2225
rect 3724 2138 4264 2191
rect 5682 2224 6222 2278
rect 5682 2190 5732 2224
rect 5790 2190 5800 2224
rect 5862 2190 5868 2224
rect 5934 2190 5936 2224
rect 5970 2190 5972 2224
rect 6038 2190 6044 2224
rect 6106 2190 6116 2224
rect 6174 2190 6222 2224
rect 5682 2138 6222 2190
rect 3120 2057 3154 2076
rect 3120 1989 3154 1991
rect 3120 1953 3154 1955
rect 3120 1868 3154 1887
rect 3278 2057 3312 2076
rect 3278 1989 3312 1991
rect 3278 1953 3312 1955
rect 3278 1868 3312 1887
rect 3742 2067 3776 2086
rect 3742 1999 3776 2001
rect 3742 1963 3776 1965
rect 3742 1878 3776 1897
rect 3900 2067 3934 2086
rect 3900 1999 3934 2001
rect 3900 1963 3934 1965
rect 3900 1878 3934 1897
rect 4050 2067 4084 2086
rect 4050 1999 4084 2001
rect 4050 1963 4084 1965
rect 4050 1878 4084 1897
rect 4208 2067 4242 2086
rect 4208 1999 4242 2001
rect 4208 1963 4242 1965
rect 4208 1878 4242 1897
rect 4402 2067 4436 2086
rect 4402 1999 4436 2001
rect 4402 1963 4436 1965
rect 4402 1878 4436 1897
rect 4560 2067 4594 2086
rect 4560 1999 4594 2001
rect 4560 1963 4594 1965
rect 4560 1878 4594 1897
rect 4710 2067 4744 2086
rect 4710 1999 4744 2001
rect 4710 1963 4744 1965
rect 4710 1878 4744 1897
rect 4868 2067 4902 2086
rect 4868 1999 4902 2001
rect 4868 1963 4902 1965
rect 4868 1878 4902 1897
rect 5700 2068 5734 2086
rect 5700 2000 5734 2002
rect 5700 1964 5734 1966
rect 5700 1878 5734 1898
rect 5858 2068 5892 2086
rect 5858 2000 5892 2002
rect 5858 1964 5892 1966
rect 5858 1878 5892 1898
rect 6008 2068 6042 2086
rect 6008 2000 6042 2002
rect 6008 1964 6042 1966
rect 6008 1878 6042 1898
rect 6166 2068 6200 2086
rect 6166 2000 6200 2002
rect 6166 1964 6200 1966
rect 6166 1878 6200 1898
rect 6360 2068 6394 2086
rect 6360 2000 6394 2002
rect 6360 1964 6394 1966
rect 6360 1878 6394 1898
rect 6518 2068 6552 2086
rect 6518 2000 6552 2002
rect 6518 1964 6552 1966
rect 6518 1878 6552 1898
rect 6668 2068 6702 2086
rect 6668 2000 6702 2002
rect 6668 1964 6702 1966
rect 6668 1878 6702 1898
rect 6826 2068 6860 2086
rect 6826 2000 6860 2002
rect 6826 1964 6860 1966
rect 6826 1878 6860 1898
rect 3670 1842 3704 1855
rect 3668 1839 3707 1842
rect 1773 1769 1807 1778
rect 2261 1771 2319 1783
rect 2625 1772 2703 1786
rect 2850 1781 2857 1815
rect 2891 1781 2898 1815
rect 3013 1781 3029 1815
rect 3063 1781 3079 1815
rect 3668 1805 3670 1839
rect 3704 1805 3707 1839
rect 3984 1833 4018 1846
rect 5628 1842 5662 1856
rect 3668 1803 3707 1805
rect 3982 1830 4021 1833
rect 3670 1789 3704 1803
rect 3982 1796 3984 1830
rect 4018 1796 4021 1830
rect 3982 1794 4021 1796
rect 4306 1825 4340 1840
rect 4306 1824 4341 1825
rect 2850 1774 2898 1781
rect 1255 1755 1318 1767
rect 2271 1765 2309 1771
rect 1410 1701 1444 1738
rect 556 1612 616 1628
rect 556 1588 565 1612
rect 606 1588 616 1612
rect 702 1612 762 1628
rect 702 1588 712 1612
rect 753 1588 762 1612
rect 846 1617 906 1634
rect 846 1594 856 1617
rect 897 1594 906 1617
rect 1000 1618 1060 1634
rect 1410 1630 1444 1667
rect 1568 1701 1602 1738
rect 1568 1630 1602 1667
rect 1698 1701 1732 1738
rect 1698 1630 1732 1667
rect 1856 1701 1890 1738
rect 1856 1630 1890 1667
rect 2030 1701 2064 1738
rect 2030 1630 2064 1667
rect 2188 1701 2222 1738
rect 2188 1630 2222 1667
rect 2352 1701 2420 1744
rect 2352 1667 2372 1701
rect 2406 1667 2420 1701
rect 1000 1594 1010 1618
rect 1051 1594 1060 1618
rect 540 1572 565 1588
rect 606 1572 632 1588
rect 540 1554 569 1572
rect 603 1554 632 1572
rect 686 1572 712 1588
rect 753 1572 778 1588
rect 686 1554 715 1572
rect 749 1554 778 1572
rect 830 1577 856 1594
rect 897 1577 922 1594
rect 830 1560 859 1577
rect 893 1560 922 1577
rect 984 1578 1010 1594
rect 1051 1578 1076 1594
rect 984 1560 1013 1578
rect 1047 1560 1076 1578
rect 1324 1524 1960 1588
rect 1324 1490 1353 1524
rect 1407 1490 1421 1524
rect 1479 1490 1489 1524
rect 1551 1490 1557 1524
rect 1623 1490 1625 1524
rect 1659 1490 1661 1524
rect 1727 1490 1733 1524
rect 1795 1490 1805 1524
rect 1863 1490 1877 1524
rect 1931 1490 1960 1524
rect 1324 1448 1960 1490
rect 2352 1499 2420 1667
rect 2530 1701 2564 1738
rect 2530 1630 2564 1667
rect 2352 1465 2369 1499
rect 2403 1465 2420 1499
rect 2352 1448 2420 1465
rect 2642 1403 2696 1772
rect 2857 1765 2891 1774
rect 3019 1771 3073 1781
rect 3984 1780 4018 1794
rect 4340 1790 4341 1824
rect 4621 1808 4637 1842
rect 4671 1808 4687 1842
rect 5626 1840 5666 1842
rect 5626 1806 5628 1840
rect 5662 1806 5666 1840
rect 5942 1834 5976 1846
rect 5626 1804 5666 1806
rect 5940 1830 5980 1834
rect 5628 1790 5662 1804
rect 5940 1796 5942 1830
rect 5976 1796 5980 1830
rect 5940 1794 5980 1796
rect 6264 1826 6298 1840
rect 6264 1824 6300 1826
rect 4306 1774 4340 1790
rect 5942 1780 5976 1794
rect 6298 1790 6300 1824
rect 6580 1808 6596 1842
rect 6630 1808 6646 1842
rect 6264 1774 6298 1790
rect 2776 1701 2810 1738
rect 2776 1630 2810 1667
rect 2934 1701 2968 1738
rect 2934 1630 2968 1667
rect 3120 1701 3154 1738
rect 3120 1630 3154 1667
rect 3278 1701 3312 1738
rect 3278 1630 3312 1667
rect 3742 1711 3776 1748
rect 3742 1640 3776 1677
rect 3900 1711 3934 1748
rect 3900 1640 3934 1677
rect 4050 1711 4084 1748
rect 4050 1640 4084 1677
rect 4208 1711 4242 1748
rect 4208 1640 4242 1677
rect 4402 1713 4436 1750
rect 4402 1642 4436 1679
rect 4560 1713 4594 1750
rect 4560 1642 4594 1679
rect 4710 1713 4744 1750
rect 4710 1642 4744 1679
rect 4868 1713 4902 1750
rect 4868 1642 4902 1679
rect 5700 1712 5734 1748
rect 5700 1640 5734 1678
rect 5858 1712 5892 1748
rect 5858 1640 5892 1678
rect 6008 1712 6042 1748
rect 6008 1640 6042 1678
rect 6166 1712 6200 1748
rect 6166 1640 6200 1678
rect 6360 1714 6394 1750
rect 6360 1642 6394 1680
rect 6518 1714 6552 1750
rect 6518 1642 6552 1680
rect 6668 1714 6702 1750
rect 6668 1642 6702 1680
rect 6826 1714 6860 1750
rect 6826 1642 6860 1680
rect 3704 1535 4244 1588
rect 3704 1501 3741 1535
rect 3787 1501 3813 1535
rect 3855 1501 3885 1535
rect 3923 1501 3957 1535
rect 3991 1501 4025 1535
rect 4063 1501 4093 1535
rect 4135 1501 4161 1535
rect 4207 1501 4244 1535
rect 3704 1448 4244 1501
rect 5662 1536 6202 1588
rect 5662 1502 5700 1536
rect 5746 1502 5772 1536
rect 5814 1502 5844 1536
rect 5882 1502 5916 1536
rect 5950 1502 5984 1536
rect 6022 1502 6052 1536
rect 6094 1502 6120 1536
rect 6166 1502 6202 1536
rect 5662 1448 6202 1502
rect 1348 998 1880 1050
rect 1348 964 1383 998
rect 1429 964 1455 998
rect 1497 964 1527 998
rect 1565 964 1599 998
rect 1633 964 1667 998
rect 1705 964 1735 998
rect 1777 964 1803 998
rect 1849 964 1880 998
rect 3724 997 4264 1050
rect 540 912 569 928
rect 603 912 632 928
rect 540 894 566 912
rect 607 894 632 912
rect 686 912 715 928
rect 749 912 778 928
rect 686 894 710 912
rect 751 894 778 912
rect 830 917 859 934
rect 893 917 922 934
rect 830 900 856 917
rect 897 900 922 917
rect 984 917 1013 934
rect 1047 917 1076 934
rect 984 900 1009 917
rect 1050 900 1076 917
rect 1348 910 1880 964
rect 2627 917 3073 971
rect 556 872 566 894
rect 607 872 616 894
rect 556 854 616 872
rect 702 872 710 894
rect 751 872 762 894
rect 702 854 762 872
rect 846 877 856 900
rect 897 877 906 900
rect 846 860 906 877
rect 1000 877 1009 900
rect 1050 877 1060 900
rect 1000 860 1060 877
rect 1410 829 1444 848
rect 1410 761 1444 763
rect 1410 725 1444 727
rect 1410 640 1444 659
rect 1568 829 1602 848
rect 1568 761 1602 763
rect 1568 725 1602 727
rect 1568 640 1602 659
rect 1698 829 1732 848
rect 1698 761 1732 763
rect 1698 725 1732 727
rect 1698 640 1732 659
rect 1856 829 1890 848
rect 1856 761 1890 763
rect 1856 725 1890 727
rect 1856 640 1890 659
rect 2030 829 2064 848
rect 2030 761 2064 763
rect 2030 725 2064 727
rect 2030 640 2064 659
rect 2188 829 2222 848
rect 2188 761 2222 763
rect 2188 725 2222 727
rect 2188 640 2222 659
rect 2372 829 2406 848
rect 2372 761 2406 763
rect 2372 725 2406 727
rect 2372 640 2406 659
rect 2530 829 2564 848
rect 2627 767 2681 917
rect 2776 829 2810 848
rect 2530 761 2564 763
rect 2530 725 2564 727
rect 2530 640 2564 659
rect 2625 745 2703 767
rect 2625 711 2647 745
rect 2681 711 2703 745
rect 1255 610 1318 622
rect 1251 591 1322 610
rect 2625 607 2703 711
rect 2776 761 2810 763
rect 2776 725 2810 727
rect 2776 640 2810 659
rect 2934 829 2968 848
rect 2934 761 2968 763
rect 2934 725 2968 727
rect 2934 640 2968 659
rect 1773 598 1807 607
rect 2271 601 2309 607
rect 1251 557 1269 591
rect 1303 557 1322 591
rect 1251 539 1322 557
rect 1766 591 1814 598
rect 1766 557 1773 591
rect 1807 557 1814 591
rect 1766 550 1814 557
rect 2261 589 2319 601
rect 2261 555 2273 589
rect 2307 555 2319 589
rect 2615 599 2713 607
rect 2615 565 2647 599
rect 2681 565 2713 599
rect 2857 594 2891 603
rect 2615 558 2713 565
rect 2850 587 2898 594
rect 3019 587 3073 917
rect 3724 963 3773 997
rect 3831 963 3841 997
rect 3903 963 3909 997
rect 3975 963 3977 997
rect 4011 963 4013 997
rect 4079 963 4085 997
rect 4147 963 4157 997
rect 4215 963 4264 997
rect 3724 910 4264 963
rect 3120 829 3154 848
rect 3120 761 3154 763
rect 3120 725 3154 727
rect 3120 640 3154 659
rect 3278 829 3312 848
rect 3278 761 3312 763
rect 3278 725 3312 727
rect 3278 640 3312 659
rect 3742 839 3776 858
rect 3742 771 3776 773
rect 3742 735 3776 737
rect 3742 650 3776 669
rect 3900 839 3934 858
rect 3900 771 3934 773
rect 3900 735 3934 737
rect 3900 650 3934 669
rect 4050 839 4084 858
rect 4050 771 4084 773
rect 4050 735 4084 737
rect 4050 650 4084 669
rect 4208 839 4242 858
rect 4208 771 4242 773
rect 4208 735 4242 737
rect 4208 650 4242 669
rect 4402 839 4436 858
rect 4402 771 4436 773
rect 4402 735 4436 737
rect 4402 650 4436 669
rect 4560 839 4594 858
rect 4560 771 4594 773
rect 4560 735 4594 737
rect 4560 650 4594 669
rect 4710 839 4744 858
rect 4710 771 4744 773
rect 4710 735 4744 737
rect 4710 650 4744 669
rect 4868 839 4902 858
rect 4868 771 4902 773
rect 4868 735 4902 737
rect 4868 650 4902 669
rect 3670 614 3704 627
rect 3668 611 3707 614
rect 1773 541 1807 550
rect 2261 543 2319 555
rect 2625 544 2703 558
rect 2850 553 2857 587
rect 2891 553 2898 587
rect 3013 553 3029 587
rect 3063 553 3079 587
rect 3668 577 3670 611
rect 3704 577 3707 611
rect 3984 605 4018 618
rect 3668 575 3707 577
rect 3982 602 4021 605
rect 3670 561 3704 575
rect 3982 568 3984 602
rect 4018 568 4021 602
rect 3982 566 4021 568
rect 4306 597 4340 612
rect 4306 596 4341 597
rect 2850 546 2898 553
rect 1255 527 1318 539
rect 2271 537 2309 543
rect 1410 473 1444 510
rect 556 384 616 400
rect 556 360 565 384
rect 606 360 616 384
rect 702 384 762 400
rect 702 360 712 384
rect 753 360 762 384
rect 846 389 906 406
rect 846 366 856 389
rect 897 366 906 389
rect 1000 390 1060 406
rect 1410 402 1444 439
rect 1568 473 1602 510
rect 1568 402 1602 439
rect 1698 473 1732 510
rect 1698 402 1732 439
rect 1856 473 1890 510
rect 1856 402 1890 439
rect 2030 473 2064 510
rect 2030 402 2064 439
rect 2188 473 2222 510
rect 2188 402 2222 439
rect 2352 473 2420 516
rect 2352 439 2372 473
rect 2406 439 2420 473
rect 1000 366 1010 390
rect 1051 366 1060 390
rect 540 344 565 360
rect 606 344 632 360
rect 540 326 569 344
rect 603 326 632 344
rect 686 344 712 360
rect 753 344 778 360
rect 686 326 715 344
rect 749 326 778 344
rect 830 349 856 366
rect 897 349 922 366
rect 830 332 859 349
rect 893 332 922 349
rect 984 350 1010 366
rect 1051 350 1076 366
rect 984 332 1013 350
rect 1047 332 1076 350
rect 1324 296 1960 360
rect 1324 262 1353 296
rect 1407 262 1421 296
rect 1479 262 1489 296
rect 1551 262 1557 296
rect 1623 262 1625 296
rect 1659 262 1661 296
rect 1727 262 1733 296
rect 1795 262 1805 296
rect 1863 262 1877 296
rect 1931 262 1960 296
rect 1324 220 1960 262
rect 2352 271 2420 439
rect 2530 473 2564 510
rect 2530 402 2564 439
rect 2352 237 2369 271
rect 2403 237 2420 271
rect 2352 220 2420 237
rect 2642 175 2696 544
rect 2857 537 2891 546
rect 3019 543 3073 553
rect 3984 552 4018 566
rect 4340 562 4341 596
rect 4621 580 4637 614
rect 4671 580 4687 614
rect 4306 546 4340 562
rect 2776 473 2810 510
rect 2776 402 2810 439
rect 2934 473 2968 510
rect 2934 402 2968 439
rect 3120 473 3154 510
rect 3120 402 3154 439
rect 3278 473 3312 510
rect 3278 402 3312 439
rect 3742 483 3776 520
rect 3742 412 3776 449
rect 3900 483 3934 520
rect 3900 412 3934 449
rect 4050 483 4084 520
rect 4050 412 4084 449
rect 4208 483 4242 520
rect 4208 412 4242 449
rect 4402 485 4436 522
rect 4402 414 4436 451
rect 4560 485 4594 522
rect 4560 414 4594 451
rect 4710 485 4744 522
rect 4710 414 4744 451
rect 4868 485 4902 522
rect 4868 414 4902 451
rect 3704 307 4244 360
rect 3704 273 3741 307
rect 3787 273 3813 307
rect 3855 273 3885 307
rect 3923 273 3957 307
rect 3991 273 4025 307
rect 4063 273 4093 307
rect 4135 273 4161 307
rect 4207 273 4244 307
rect 3704 220 4244 273
<< viali >>
rect 1383 4648 1395 4682
rect 1395 4648 1417 4682
rect 1455 4648 1463 4682
rect 1463 4648 1489 4682
rect 1527 4648 1531 4682
rect 1531 4648 1561 4682
rect 1599 4648 1633 4682
rect 1671 4648 1701 4682
rect 1701 4648 1705 4682
rect 1743 4648 1769 4682
rect 1769 4648 1777 4682
rect 1815 4648 1837 4682
rect 1837 4648 1849 4682
rect 566 4578 569 4596
rect 569 4578 603 4596
rect 603 4578 607 4596
rect 710 4578 715 4596
rect 715 4578 749 4596
rect 749 4578 751 4596
rect 856 4584 859 4601
rect 859 4584 893 4601
rect 893 4584 897 4601
rect 1009 4584 1013 4601
rect 1013 4584 1047 4601
rect 1047 4584 1050 4601
rect 566 4556 607 4578
rect 710 4556 751 4578
rect 856 4561 897 4584
rect 1009 4561 1050 4584
rect 1410 4479 1444 4481
rect 1410 4447 1444 4479
rect 1410 4377 1444 4409
rect 1410 4375 1444 4377
rect 1568 4479 1602 4481
rect 1568 4447 1602 4479
rect 1568 4377 1602 4409
rect 1568 4375 1602 4377
rect 1698 4479 1732 4481
rect 1698 4447 1732 4479
rect 1698 4377 1732 4409
rect 1698 4375 1732 4377
rect 1856 4479 1890 4481
rect 1856 4447 1890 4479
rect 1856 4377 1890 4409
rect 1856 4375 1890 4377
rect 2030 4479 2064 4481
rect 2030 4447 2064 4479
rect 2030 4377 2064 4409
rect 2030 4375 2064 4377
rect 2188 4479 2222 4481
rect 2188 4447 2222 4479
rect 2188 4377 2222 4409
rect 2188 4375 2222 4377
rect 2372 4479 2406 4481
rect 2372 4447 2406 4479
rect 2372 4377 2406 4409
rect 2372 4375 2406 4377
rect 2530 4479 2564 4481
rect 2530 4447 2564 4479
rect 2776 4479 2810 4481
rect 2530 4377 2564 4409
rect 2530 4375 2564 4377
rect 2647 4395 2681 4429
rect 2776 4447 2810 4479
rect 2776 4377 2810 4409
rect 2776 4375 2810 4377
rect 2934 4479 2968 4481
rect 2934 4447 2968 4479
rect 2934 4377 2968 4409
rect 2934 4375 2968 4377
rect 1269 4241 1303 4275
rect 1773 4241 1807 4275
rect 2273 4239 2307 4273
rect 3797 4647 3807 4681
rect 3807 4647 3831 4681
rect 3869 4647 3875 4681
rect 3875 4647 3903 4681
rect 3941 4647 3943 4681
rect 3943 4647 3975 4681
rect 4013 4647 4045 4681
rect 4045 4647 4047 4681
rect 4085 4647 4113 4681
rect 4113 4647 4119 4681
rect 4157 4647 4181 4681
rect 4181 4647 4191 4681
rect 5756 4646 5766 4680
rect 5766 4646 5790 4680
rect 5828 4646 5834 4680
rect 5834 4646 5862 4680
rect 5900 4646 5902 4680
rect 5902 4646 5934 4680
rect 5972 4646 6004 4680
rect 6004 4646 6006 4680
rect 6044 4646 6072 4680
rect 6072 4646 6078 4680
rect 6116 4646 6140 4680
rect 6140 4646 6150 4680
rect 3120 4479 3154 4481
rect 3120 4447 3154 4479
rect 3120 4377 3154 4409
rect 3120 4375 3154 4377
rect 3278 4479 3312 4481
rect 3278 4447 3312 4479
rect 3278 4377 3312 4409
rect 3278 4375 3312 4377
rect 3742 4489 3776 4491
rect 3742 4457 3776 4489
rect 3742 4387 3776 4419
rect 3742 4385 3776 4387
rect 3900 4489 3934 4491
rect 3900 4457 3934 4489
rect 3900 4387 3934 4419
rect 3900 4385 3934 4387
rect 4050 4489 4084 4491
rect 4050 4457 4084 4489
rect 4050 4387 4084 4419
rect 4050 4385 4084 4387
rect 4208 4489 4242 4491
rect 4208 4457 4242 4489
rect 4208 4387 4242 4419
rect 4208 4385 4242 4387
rect 4402 4489 4436 4491
rect 4402 4457 4436 4489
rect 4402 4387 4436 4419
rect 4402 4385 4436 4387
rect 4560 4489 4594 4491
rect 4560 4457 4594 4489
rect 4560 4387 4594 4419
rect 4560 4385 4594 4387
rect 4710 4489 4744 4491
rect 4710 4457 4744 4489
rect 4710 4387 4744 4419
rect 4710 4385 4744 4387
rect 4868 4489 4902 4491
rect 4868 4457 4902 4489
rect 4868 4387 4902 4419
rect 4868 4385 4902 4387
rect 5700 4490 5734 4492
rect 5700 4458 5734 4490
rect 5700 4388 5734 4420
rect 5700 4386 5734 4388
rect 5858 4490 5892 4492
rect 5858 4458 5892 4490
rect 5858 4388 5892 4420
rect 5858 4386 5892 4388
rect 6008 4490 6042 4492
rect 6008 4458 6042 4490
rect 6008 4388 6042 4420
rect 6008 4386 6042 4388
rect 6166 4490 6200 4492
rect 6166 4458 6200 4490
rect 6166 4388 6200 4420
rect 6166 4386 6200 4388
rect 6360 4490 6394 4492
rect 6360 4458 6394 4490
rect 6360 4388 6394 4420
rect 6360 4386 6394 4388
rect 6518 4490 6552 4492
rect 6518 4458 6552 4490
rect 6518 4388 6552 4420
rect 6518 4386 6552 4388
rect 6668 4490 6702 4492
rect 6668 4458 6702 4490
rect 6668 4388 6702 4420
rect 6668 4386 6702 4388
rect 6826 4490 6860 4492
rect 6826 4458 6860 4490
rect 6826 4388 6860 4420
rect 6826 4386 6860 4388
rect 2857 4237 2891 4271
rect 3670 4261 3704 4295
rect 3984 4252 4018 4286
rect 1410 4123 1444 4157
rect 565 4044 606 4068
rect 712 4044 753 4068
rect 856 4050 897 4073
rect 1568 4123 1602 4157
rect 1698 4123 1732 4157
rect 1856 4123 1890 4157
rect 2030 4123 2064 4157
rect 2188 4123 2222 4157
rect 2372 4123 2406 4157
rect 1010 4050 1051 4074
rect 565 4028 569 4044
rect 569 4028 603 4044
rect 603 4028 606 4044
rect 712 4028 715 4044
rect 715 4028 749 4044
rect 749 4028 753 4044
rect 856 4033 859 4050
rect 859 4033 893 4050
rect 893 4033 897 4050
rect 1010 4034 1013 4050
rect 1013 4034 1047 4050
rect 1047 4034 1051 4050
rect 1373 3946 1387 3980
rect 1387 3946 1407 3980
rect 1445 3946 1455 3980
rect 1455 3946 1479 3980
rect 1517 3946 1523 3980
rect 1523 3946 1551 3980
rect 1589 3946 1591 3980
rect 1591 3946 1623 3980
rect 1661 3946 1693 3980
rect 1693 3946 1695 3980
rect 1733 3946 1761 3980
rect 1761 3946 1767 3980
rect 1805 3946 1829 3980
rect 1829 3946 1839 3980
rect 1877 3946 1897 3980
rect 1897 3946 1911 3980
rect 2530 4123 2564 4157
rect 2369 3921 2403 3955
rect 4306 4246 4340 4280
rect 4637 4264 4671 4298
rect 5628 4262 5662 4296
rect 5942 4252 5976 4286
rect 6264 4246 6298 4280
rect 6596 4264 6630 4298
rect 2776 4123 2810 4157
rect 2934 4123 2968 4157
rect 3120 4123 3154 4157
rect 3278 4123 3312 4157
rect 3742 4133 3776 4167
rect 3900 4133 3934 4167
rect 4050 4133 4084 4167
rect 4208 4133 4242 4167
rect 4402 4135 4436 4169
rect 4560 4135 4594 4169
rect 4710 4135 4744 4169
rect 4868 4135 4902 4169
rect 5700 4134 5734 4168
rect 5858 4134 5892 4168
rect 6008 4134 6042 4168
rect 6166 4134 6200 4168
rect 6360 4136 6394 4170
rect 6518 4136 6552 4170
rect 6668 4136 6702 4170
rect 6826 4136 6860 4170
rect 3741 3957 3753 3991
rect 3753 3957 3775 3991
rect 3813 3957 3821 3991
rect 3821 3957 3847 3991
rect 3885 3957 3889 3991
rect 3889 3957 3919 3991
rect 3957 3957 3991 3991
rect 4029 3957 4059 3991
rect 4059 3957 4063 3991
rect 4101 3957 4127 3991
rect 4127 3957 4135 3991
rect 4173 3957 4195 3991
rect 4195 3957 4207 3991
rect 5700 3958 5712 3992
rect 5712 3958 5734 3992
rect 5772 3958 5780 3992
rect 5780 3958 5806 3992
rect 5844 3958 5848 3992
rect 5848 3958 5878 3992
rect 5916 3958 5950 3992
rect 5988 3958 6018 3992
rect 6018 3958 6022 3992
rect 6060 3958 6086 3992
rect 6086 3958 6094 3992
rect 6132 3958 6154 3992
rect 6154 3958 6166 3992
rect 2642 3805 2696 3859
rect 1383 3420 1395 3454
rect 1395 3420 1417 3454
rect 1455 3420 1463 3454
rect 1463 3420 1489 3454
rect 1527 3420 1531 3454
rect 1531 3420 1561 3454
rect 1599 3420 1633 3454
rect 1671 3420 1701 3454
rect 1701 3420 1705 3454
rect 1743 3420 1769 3454
rect 1769 3420 1777 3454
rect 1815 3420 1837 3454
rect 1837 3420 1849 3454
rect 566 3350 569 3368
rect 569 3350 603 3368
rect 603 3350 607 3368
rect 710 3350 715 3368
rect 715 3350 749 3368
rect 749 3350 751 3368
rect 856 3356 859 3373
rect 859 3356 893 3373
rect 893 3356 897 3373
rect 1009 3356 1013 3373
rect 1013 3356 1047 3373
rect 1047 3356 1050 3373
rect 566 3328 607 3350
rect 710 3328 751 3350
rect 856 3333 897 3356
rect 1009 3333 1050 3356
rect 1410 3251 1444 3253
rect 1410 3219 1444 3251
rect 1410 3149 1444 3181
rect 1410 3147 1444 3149
rect 1568 3251 1602 3253
rect 1568 3219 1602 3251
rect 1568 3149 1602 3181
rect 1568 3147 1602 3149
rect 1698 3251 1732 3253
rect 1698 3219 1732 3251
rect 1698 3149 1732 3181
rect 1698 3147 1732 3149
rect 1856 3251 1890 3253
rect 1856 3219 1890 3251
rect 1856 3149 1890 3181
rect 1856 3147 1890 3149
rect 2030 3251 2064 3253
rect 2030 3219 2064 3251
rect 2030 3149 2064 3181
rect 2030 3147 2064 3149
rect 2188 3251 2222 3253
rect 2188 3219 2222 3251
rect 2188 3149 2222 3181
rect 2188 3147 2222 3149
rect 2372 3251 2406 3253
rect 2372 3219 2406 3251
rect 2372 3149 2406 3181
rect 2372 3147 2406 3149
rect 2530 3251 2564 3253
rect 2530 3219 2564 3251
rect 2776 3251 2810 3253
rect 2530 3149 2564 3181
rect 2530 3147 2564 3149
rect 2647 3167 2681 3201
rect 2776 3219 2810 3251
rect 2776 3149 2810 3181
rect 2776 3147 2810 3149
rect 2934 3251 2968 3253
rect 2934 3219 2968 3251
rect 2934 3149 2968 3181
rect 2934 3147 2968 3149
rect 1269 3013 1303 3047
rect 1773 3013 1807 3047
rect 2273 3011 2307 3045
rect 3797 3419 3807 3453
rect 3807 3419 3831 3453
rect 3869 3419 3875 3453
rect 3875 3419 3903 3453
rect 3941 3419 3943 3453
rect 3943 3419 3975 3453
rect 4013 3419 4045 3453
rect 4045 3419 4047 3453
rect 4085 3419 4113 3453
rect 4113 3419 4119 3453
rect 4157 3419 4181 3453
rect 4181 3419 4191 3453
rect 5756 3418 5766 3452
rect 5766 3418 5790 3452
rect 5828 3418 5834 3452
rect 5834 3418 5862 3452
rect 5900 3418 5902 3452
rect 5902 3418 5934 3452
rect 5972 3418 6004 3452
rect 6004 3418 6006 3452
rect 6044 3418 6072 3452
rect 6072 3418 6078 3452
rect 6116 3418 6140 3452
rect 6140 3418 6150 3452
rect 3120 3251 3154 3253
rect 3120 3219 3154 3251
rect 3120 3149 3154 3181
rect 3120 3147 3154 3149
rect 3278 3251 3312 3253
rect 3278 3219 3312 3251
rect 3278 3149 3312 3181
rect 3278 3147 3312 3149
rect 3742 3261 3776 3263
rect 3742 3229 3776 3261
rect 3742 3159 3776 3191
rect 3742 3157 3776 3159
rect 3900 3261 3934 3263
rect 3900 3229 3934 3261
rect 3900 3159 3934 3191
rect 3900 3157 3934 3159
rect 4050 3261 4084 3263
rect 4050 3229 4084 3261
rect 4050 3159 4084 3191
rect 4050 3157 4084 3159
rect 4208 3261 4242 3263
rect 4208 3229 4242 3261
rect 4208 3159 4242 3191
rect 4208 3157 4242 3159
rect 4402 3261 4436 3263
rect 4402 3229 4436 3261
rect 4402 3159 4436 3191
rect 4402 3157 4436 3159
rect 4560 3261 4594 3263
rect 4560 3229 4594 3261
rect 4560 3159 4594 3191
rect 4560 3157 4594 3159
rect 4710 3261 4744 3263
rect 4710 3229 4744 3261
rect 4710 3159 4744 3191
rect 4710 3157 4744 3159
rect 4868 3261 4902 3263
rect 4868 3229 4902 3261
rect 4868 3159 4902 3191
rect 4868 3157 4902 3159
rect 5700 3262 5734 3264
rect 5700 3230 5734 3262
rect 5700 3160 5734 3192
rect 5700 3158 5734 3160
rect 5858 3262 5892 3264
rect 5858 3230 5892 3262
rect 5858 3160 5892 3192
rect 5858 3158 5892 3160
rect 6008 3262 6042 3264
rect 6008 3230 6042 3262
rect 6008 3160 6042 3192
rect 6008 3158 6042 3160
rect 6166 3262 6200 3264
rect 6166 3230 6200 3262
rect 6166 3160 6200 3192
rect 6166 3158 6200 3160
rect 6360 3262 6394 3264
rect 6360 3230 6394 3262
rect 6360 3160 6394 3192
rect 6360 3158 6394 3160
rect 6518 3262 6552 3264
rect 6518 3230 6552 3262
rect 6518 3160 6552 3192
rect 6518 3158 6552 3160
rect 6668 3262 6702 3264
rect 6668 3230 6702 3262
rect 6668 3160 6702 3192
rect 6668 3158 6702 3160
rect 6826 3262 6860 3264
rect 6826 3230 6860 3262
rect 6826 3160 6860 3192
rect 6826 3158 6860 3160
rect 2857 3009 2891 3043
rect 3670 3033 3704 3067
rect 3984 3024 4018 3058
rect 1410 2895 1444 2929
rect 565 2816 606 2840
rect 712 2816 753 2840
rect 856 2822 897 2845
rect 1568 2895 1602 2929
rect 1698 2895 1732 2929
rect 1856 2895 1890 2929
rect 2030 2895 2064 2929
rect 2188 2895 2222 2929
rect 2372 2895 2406 2929
rect 1010 2822 1051 2846
rect 565 2800 569 2816
rect 569 2800 603 2816
rect 603 2800 606 2816
rect 712 2800 715 2816
rect 715 2800 749 2816
rect 749 2800 753 2816
rect 856 2805 859 2822
rect 859 2805 893 2822
rect 893 2805 897 2822
rect 1010 2806 1013 2822
rect 1013 2806 1047 2822
rect 1047 2806 1051 2822
rect 1373 2718 1387 2752
rect 1387 2718 1407 2752
rect 1445 2718 1455 2752
rect 1455 2718 1479 2752
rect 1517 2718 1523 2752
rect 1523 2718 1551 2752
rect 1589 2718 1591 2752
rect 1591 2718 1623 2752
rect 1661 2718 1693 2752
rect 1693 2718 1695 2752
rect 1733 2718 1761 2752
rect 1761 2718 1767 2752
rect 1805 2718 1829 2752
rect 1829 2718 1839 2752
rect 1877 2718 1897 2752
rect 1897 2718 1911 2752
rect 2530 2895 2564 2929
rect 2369 2693 2403 2727
rect 4306 3018 4340 3052
rect 4637 3036 4671 3070
rect 5628 3034 5662 3068
rect 5942 3024 5976 3058
rect 6264 3018 6298 3052
rect 6596 3036 6630 3070
rect 2776 2895 2810 2929
rect 2934 2895 2968 2929
rect 3120 2895 3154 2929
rect 3278 2895 3312 2929
rect 3742 2905 3776 2939
rect 3900 2905 3934 2939
rect 4050 2905 4084 2939
rect 4208 2905 4242 2939
rect 4402 2907 4436 2941
rect 4560 2907 4594 2941
rect 4710 2907 4744 2941
rect 4868 2907 4902 2941
rect 5700 2906 5734 2940
rect 5858 2906 5892 2940
rect 6008 2906 6042 2940
rect 6166 2906 6200 2940
rect 6360 2908 6394 2942
rect 6518 2908 6552 2942
rect 6668 2908 6702 2942
rect 6826 2908 6860 2942
rect 3741 2729 3753 2763
rect 3753 2729 3775 2763
rect 3813 2729 3821 2763
rect 3821 2729 3847 2763
rect 3885 2729 3889 2763
rect 3889 2729 3919 2763
rect 3957 2729 3991 2763
rect 4029 2729 4059 2763
rect 4059 2729 4063 2763
rect 4101 2729 4127 2763
rect 4127 2729 4135 2763
rect 4173 2729 4195 2763
rect 4195 2729 4207 2763
rect 5700 2730 5712 2764
rect 5712 2730 5734 2764
rect 5772 2730 5780 2764
rect 5780 2730 5806 2764
rect 5844 2730 5848 2764
rect 5848 2730 5878 2764
rect 5916 2730 5950 2764
rect 5988 2730 6018 2764
rect 6018 2730 6022 2764
rect 6060 2730 6086 2764
rect 6086 2730 6094 2764
rect 6132 2730 6154 2764
rect 6154 2730 6166 2764
rect 2642 2577 2696 2631
rect 1383 2192 1395 2226
rect 1395 2192 1417 2226
rect 1455 2192 1463 2226
rect 1463 2192 1489 2226
rect 1527 2192 1531 2226
rect 1531 2192 1561 2226
rect 1599 2192 1633 2226
rect 1671 2192 1701 2226
rect 1701 2192 1705 2226
rect 1743 2192 1769 2226
rect 1769 2192 1777 2226
rect 1815 2192 1837 2226
rect 1837 2192 1849 2226
rect 566 2122 569 2140
rect 569 2122 603 2140
rect 603 2122 607 2140
rect 710 2122 715 2140
rect 715 2122 749 2140
rect 749 2122 751 2140
rect 856 2128 859 2145
rect 859 2128 893 2145
rect 893 2128 897 2145
rect 1009 2128 1013 2145
rect 1013 2128 1047 2145
rect 1047 2128 1050 2145
rect 566 2100 607 2122
rect 710 2100 751 2122
rect 856 2105 897 2128
rect 1009 2105 1050 2128
rect 1410 2023 1444 2025
rect 1410 1991 1444 2023
rect 1410 1921 1444 1953
rect 1410 1919 1444 1921
rect 1568 2023 1602 2025
rect 1568 1991 1602 2023
rect 1568 1921 1602 1953
rect 1568 1919 1602 1921
rect 1698 2023 1732 2025
rect 1698 1991 1732 2023
rect 1698 1921 1732 1953
rect 1698 1919 1732 1921
rect 1856 2023 1890 2025
rect 1856 1991 1890 2023
rect 1856 1921 1890 1953
rect 1856 1919 1890 1921
rect 2030 2023 2064 2025
rect 2030 1991 2064 2023
rect 2030 1921 2064 1953
rect 2030 1919 2064 1921
rect 2188 2023 2222 2025
rect 2188 1991 2222 2023
rect 2188 1921 2222 1953
rect 2188 1919 2222 1921
rect 2372 2023 2406 2025
rect 2372 1991 2406 2023
rect 2372 1921 2406 1953
rect 2372 1919 2406 1921
rect 2530 2023 2564 2025
rect 2530 1991 2564 2023
rect 2776 2023 2810 2025
rect 2530 1921 2564 1953
rect 2530 1919 2564 1921
rect 2647 1939 2681 1973
rect 2776 1991 2810 2023
rect 2776 1921 2810 1953
rect 2776 1919 2810 1921
rect 2934 2023 2968 2025
rect 2934 1991 2968 2023
rect 2934 1921 2968 1953
rect 2934 1919 2968 1921
rect 1269 1785 1303 1819
rect 1773 1785 1807 1819
rect 2273 1783 2307 1817
rect 3797 2191 3807 2225
rect 3807 2191 3831 2225
rect 3869 2191 3875 2225
rect 3875 2191 3903 2225
rect 3941 2191 3943 2225
rect 3943 2191 3975 2225
rect 4013 2191 4045 2225
rect 4045 2191 4047 2225
rect 4085 2191 4113 2225
rect 4113 2191 4119 2225
rect 4157 2191 4181 2225
rect 4181 2191 4191 2225
rect 5756 2190 5766 2224
rect 5766 2190 5790 2224
rect 5828 2190 5834 2224
rect 5834 2190 5862 2224
rect 5900 2190 5902 2224
rect 5902 2190 5934 2224
rect 5972 2190 6004 2224
rect 6004 2190 6006 2224
rect 6044 2190 6072 2224
rect 6072 2190 6078 2224
rect 6116 2190 6140 2224
rect 6140 2190 6150 2224
rect 3120 2023 3154 2025
rect 3120 1991 3154 2023
rect 3120 1921 3154 1953
rect 3120 1919 3154 1921
rect 3278 2023 3312 2025
rect 3278 1991 3312 2023
rect 3278 1921 3312 1953
rect 3278 1919 3312 1921
rect 3742 2033 3776 2035
rect 3742 2001 3776 2033
rect 3742 1931 3776 1963
rect 3742 1929 3776 1931
rect 3900 2033 3934 2035
rect 3900 2001 3934 2033
rect 3900 1931 3934 1963
rect 3900 1929 3934 1931
rect 4050 2033 4084 2035
rect 4050 2001 4084 2033
rect 4050 1931 4084 1963
rect 4050 1929 4084 1931
rect 4208 2033 4242 2035
rect 4208 2001 4242 2033
rect 4208 1931 4242 1963
rect 4208 1929 4242 1931
rect 4402 2033 4436 2035
rect 4402 2001 4436 2033
rect 4402 1931 4436 1963
rect 4402 1929 4436 1931
rect 4560 2033 4594 2035
rect 4560 2001 4594 2033
rect 4560 1931 4594 1963
rect 4560 1929 4594 1931
rect 4710 2033 4744 2035
rect 4710 2001 4744 2033
rect 4710 1931 4744 1963
rect 4710 1929 4744 1931
rect 4868 2033 4902 2035
rect 4868 2001 4902 2033
rect 4868 1931 4902 1963
rect 4868 1929 4902 1931
rect 5700 2034 5734 2036
rect 5700 2002 5734 2034
rect 5700 1932 5734 1964
rect 5700 1930 5734 1932
rect 5858 2034 5892 2036
rect 5858 2002 5892 2034
rect 5858 1932 5892 1964
rect 5858 1930 5892 1932
rect 6008 2034 6042 2036
rect 6008 2002 6042 2034
rect 6008 1932 6042 1964
rect 6008 1930 6042 1932
rect 6166 2034 6200 2036
rect 6166 2002 6200 2034
rect 6166 1932 6200 1964
rect 6166 1930 6200 1932
rect 6360 2034 6394 2036
rect 6360 2002 6394 2034
rect 6360 1932 6394 1964
rect 6360 1930 6394 1932
rect 6518 2034 6552 2036
rect 6518 2002 6552 2034
rect 6518 1932 6552 1964
rect 6518 1930 6552 1932
rect 6668 2034 6702 2036
rect 6668 2002 6702 2034
rect 6668 1932 6702 1964
rect 6668 1930 6702 1932
rect 6826 2034 6860 2036
rect 6826 2002 6860 2034
rect 6826 1932 6860 1964
rect 6826 1930 6860 1932
rect 2857 1781 2891 1815
rect 3670 1805 3704 1839
rect 3984 1796 4018 1830
rect 1410 1667 1444 1701
rect 565 1588 606 1612
rect 712 1588 753 1612
rect 856 1594 897 1617
rect 1568 1667 1602 1701
rect 1698 1667 1732 1701
rect 1856 1667 1890 1701
rect 2030 1667 2064 1701
rect 2188 1667 2222 1701
rect 2372 1667 2406 1701
rect 1010 1594 1051 1618
rect 565 1572 569 1588
rect 569 1572 603 1588
rect 603 1572 606 1588
rect 712 1572 715 1588
rect 715 1572 749 1588
rect 749 1572 753 1588
rect 856 1577 859 1594
rect 859 1577 893 1594
rect 893 1577 897 1594
rect 1010 1578 1013 1594
rect 1013 1578 1047 1594
rect 1047 1578 1051 1594
rect 1373 1490 1387 1524
rect 1387 1490 1407 1524
rect 1445 1490 1455 1524
rect 1455 1490 1479 1524
rect 1517 1490 1523 1524
rect 1523 1490 1551 1524
rect 1589 1490 1591 1524
rect 1591 1490 1623 1524
rect 1661 1490 1693 1524
rect 1693 1490 1695 1524
rect 1733 1490 1761 1524
rect 1761 1490 1767 1524
rect 1805 1490 1829 1524
rect 1829 1490 1839 1524
rect 1877 1490 1897 1524
rect 1897 1490 1911 1524
rect 2530 1667 2564 1701
rect 2369 1465 2403 1499
rect 4306 1790 4340 1824
rect 4637 1808 4671 1842
rect 5628 1806 5662 1840
rect 5942 1796 5976 1830
rect 6264 1790 6298 1824
rect 6596 1808 6630 1842
rect 2776 1667 2810 1701
rect 2934 1667 2968 1701
rect 3120 1667 3154 1701
rect 3278 1667 3312 1701
rect 3742 1677 3776 1711
rect 3900 1677 3934 1711
rect 4050 1677 4084 1711
rect 4208 1677 4242 1711
rect 4402 1679 4436 1713
rect 4560 1679 4594 1713
rect 4710 1679 4744 1713
rect 4868 1679 4902 1713
rect 5700 1678 5734 1712
rect 5858 1678 5892 1712
rect 6008 1678 6042 1712
rect 6166 1678 6200 1712
rect 6360 1680 6394 1714
rect 6518 1680 6552 1714
rect 6668 1680 6702 1714
rect 6826 1680 6860 1714
rect 3741 1501 3753 1535
rect 3753 1501 3775 1535
rect 3813 1501 3821 1535
rect 3821 1501 3847 1535
rect 3885 1501 3889 1535
rect 3889 1501 3919 1535
rect 3957 1501 3991 1535
rect 4029 1501 4059 1535
rect 4059 1501 4063 1535
rect 4101 1501 4127 1535
rect 4127 1501 4135 1535
rect 4173 1501 4195 1535
rect 4195 1501 4207 1535
rect 5700 1502 5712 1536
rect 5712 1502 5734 1536
rect 5772 1502 5780 1536
rect 5780 1502 5806 1536
rect 5844 1502 5848 1536
rect 5848 1502 5878 1536
rect 5916 1502 5950 1536
rect 5988 1502 6018 1536
rect 6018 1502 6022 1536
rect 6060 1502 6086 1536
rect 6086 1502 6094 1536
rect 6132 1502 6154 1536
rect 6154 1502 6166 1536
rect 2642 1349 2696 1403
rect 1383 964 1395 998
rect 1395 964 1417 998
rect 1455 964 1463 998
rect 1463 964 1489 998
rect 1527 964 1531 998
rect 1531 964 1561 998
rect 1599 964 1633 998
rect 1671 964 1701 998
rect 1701 964 1705 998
rect 1743 964 1769 998
rect 1769 964 1777 998
rect 1815 964 1837 998
rect 1837 964 1849 998
rect 566 894 569 912
rect 569 894 603 912
rect 603 894 607 912
rect 710 894 715 912
rect 715 894 749 912
rect 749 894 751 912
rect 856 900 859 917
rect 859 900 893 917
rect 893 900 897 917
rect 1009 900 1013 917
rect 1013 900 1047 917
rect 1047 900 1050 917
rect 566 872 607 894
rect 710 872 751 894
rect 856 877 897 900
rect 1009 877 1050 900
rect 1410 795 1444 797
rect 1410 763 1444 795
rect 1410 693 1444 725
rect 1410 691 1444 693
rect 1568 795 1602 797
rect 1568 763 1602 795
rect 1568 693 1602 725
rect 1568 691 1602 693
rect 1698 795 1732 797
rect 1698 763 1732 795
rect 1698 693 1732 725
rect 1698 691 1732 693
rect 1856 795 1890 797
rect 1856 763 1890 795
rect 1856 693 1890 725
rect 1856 691 1890 693
rect 2030 795 2064 797
rect 2030 763 2064 795
rect 2030 693 2064 725
rect 2030 691 2064 693
rect 2188 795 2222 797
rect 2188 763 2222 795
rect 2188 693 2222 725
rect 2188 691 2222 693
rect 2372 795 2406 797
rect 2372 763 2406 795
rect 2372 693 2406 725
rect 2372 691 2406 693
rect 2530 795 2564 797
rect 2530 763 2564 795
rect 2776 795 2810 797
rect 2530 693 2564 725
rect 2530 691 2564 693
rect 2647 711 2681 745
rect 2776 763 2810 795
rect 2776 693 2810 725
rect 2776 691 2810 693
rect 2934 795 2968 797
rect 2934 763 2968 795
rect 2934 693 2968 725
rect 2934 691 2968 693
rect 1269 557 1303 591
rect 1773 557 1807 591
rect 2273 555 2307 589
rect 3797 963 3807 997
rect 3807 963 3831 997
rect 3869 963 3875 997
rect 3875 963 3903 997
rect 3941 963 3943 997
rect 3943 963 3975 997
rect 4013 963 4045 997
rect 4045 963 4047 997
rect 4085 963 4113 997
rect 4113 963 4119 997
rect 4157 963 4181 997
rect 4181 963 4191 997
rect 3120 795 3154 797
rect 3120 763 3154 795
rect 3120 693 3154 725
rect 3120 691 3154 693
rect 3278 795 3312 797
rect 3278 763 3312 795
rect 3278 693 3312 725
rect 3278 691 3312 693
rect 3742 805 3776 807
rect 3742 773 3776 805
rect 3742 703 3776 735
rect 3742 701 3776 703
rect 3900 805 3934 807
rect 3900 773 3934 805
rect 3900 703 3934 735
rect 3900 701 3934 703
rect 4050 805 4084 807
rect 4050 773 4084 805
rect 4050 703 4084 735
rect 4050 701 4084 703
rect 4208 805 4242 807
rect 4208 773 4242 805
rect 4208 703 4242 735
rect 4208 701 4242 703
rect 4402 805 4436 807
rect 4402 773 4436 805
rect 4402 703 4436 735
rect 4402 701 4436 703
rect 4560 805 4594 807
rect 4560 773 4594 805
rect 4560 703 4594 735
rect 4560 701 4594 703
rect 4710 805 4744 807
rect 4710 773 4744 805
rect 4710 703 4744 735
rect 4710 701 4744 703
rect 4868 805 4902 807
rect 4868 773 4902 805
rect 4868 703 4902 735
rect 4868 701 4902 703
rect 2857 553 2891 587
rect 3670 577 3704 611
rect 3984 568 4018 602
rect 1410 439 1444 473
rect 565 360 606 384
rect 712 360 753 384
rect 856 366 897 389
rect 1568 439 1602 473
rect 1698 439 1732 473
rect 1856 439 1890 473
rect 2030 439 2064 473
rect 2188 439 2222 473
rect 2372 439 2406 473
rect 1010 366 1051 390
rect 565 344 569 360
rect 569 344 603 360
rect 603 344 606 360
rect 712 344 715 360
rect 715 344 749 360
rect 749 344 753 360
rect 856 349 859 366
rect 859 349 893 366
rect 893 349 897 366
rect 1010 350 1013 366
rect 1013 350 1047 366
rect 1047 350 1051 366
rect 1373 262 1387 296
rect 1387 262 1407 296
rect 1445 262 1455 296
rect 1455 262 1479 296
rect 1517 262 1523 296
rect 1523 262 1551 296
rect 1589 262 1591 296
rect 1591 262 1623 296
rect 1661 262 1693 296
rect 1693 262 1695 296
rect 1733 262 1761 296
rect 1761 262 1767 296
rect 1805 262 1829 296
rect 1829 262 1839 296
rect 1877 262 1897 296
rect 1897 262 1911 296
rect 2530 439 2564 473
rect 2369 237 2403 271
rect 4306 562 4340 596
rect 4637 580 4671 614
rect 2776 439 2810 473
rect 2934 439 2968 473
rect 3120 439 3154 473
rect 3278 439 3312 473
rect 3742 449 3776 483
rect 3900 449 3934 483
rect 4050 449 4084 483
rect 4208 449 4242 483
rect 4402 451 4436 485
rect 4560 451 4594 485
rect 4710 451 4744 485
rect 4868 451 4902 485
rect 3741 273 3753 307
rect 3753 273 3775 307
rect 3813 273 3821 307
rect 3821 273 3847 307
rect 3885 273 3889 307
rect 3889 273 3919 307
rect 3957 273 3991 307
rect 4029 273 4059 307
rect 4059 273 4063 307
rect 4101 273 4127 307
rect 4127 273 4135 307
rect 4173 273 4195 307
rect 4195 273 4207 307
rect 2642 121 2696 175
<< metal1 >>
rect 5029 4872 5081 4878
rect 3472 4825 4907 4864
rect 1348 4691 1880 4734
rect 1348 4682 1398 4691
rect 1450 4682 1462 4691
rect 1348 4648 1383 4682
rect 1450 4648 1455 4682
rect 1348 4639 1398 4648
rect 1450 4639 1462 4648
rect 1514 4639 1526 4691
rect 1578 4639 1590 4691
rect 1642 4639 1654 4691
rect 1706 4639 1718 4691
rect 1770 4682 1782 4691
rect 1834 4682 1880 4691
rect 1777 4648 1782 4682
rect 1849 4648 1880 4682
rect 3472 4667 3511 4825
rect 4738 4783 4744 4790
rect 4558 4744 4744 4783
rect 1770 4639 1782 4648
rect 1834 4639 1880 4648
rect 550 4620 622 4624
rect 550 4568 560 4620
rect 612 4568 622 4620
rect 696 4618 768 4624
rect 550 4556 566 4568
rect 607 4556 622 4568
rect 682 4616 768 4618
rect 682 4564 702 4616
rect 754 4564 768 4616
rect 682 4562 710 4564
rect 550 4526 622 4556
rect 696 4556 710 4562
rect 751 4556 768 4564
rect 696 4526 768 4556
rect 840 4601 912 4630
rect 840 4561 856 4601
rect 897 4561 912 4601
rect 840 4532 912 4561
rect 994 4601 1066 4630
rect 994 4561 1009 4601
rect 1050 4561 1066 4601
rect 1348 4594 1880 4639
rect 994 4532 1066 4561
rect 564 4486 608 4526
rect 856 4466 900 4532
rect 378 4458 433 4464
rect 846 4414 852 4466
rect 904 4414 910 4466
rect 378 4173 433 4403
rect 856 4374 900 4414
rect 1008 4374 1052 4532
rect 1407 4528 1448 4594
rect 1693 4528 1735 4594
rect 1941 4591 2687 4636
rect 1404 4481 1450 4528
rect 1404 4447 1410 4481
rect 1444 4447 1450 4481
rect 1404 4409 1450 4447
rect 1404 4375 1410 4409
rect 1444 4375 1450 4409
rect 708 4330 900 4374
rect 372 4118 378 4173
rect 433 4118 439 4173
rect 708 4096 752 4330
rect 998 4322 1004 4374
rect 1056 4322 1062 4374
rect 1404 4328 1450 4375
rect 1562 4481 1608 4528
rect 1562 4447 1568 4481
rect 1602 4447 1608 4481
rect 1562 4409 1608 4447
rect 1562 4375 1568 4409
rect 1602 4375 1608 4409
rect 1562 4328 1608 4375
rect 1692 4481 1738 4528
rect 1692 4447 1698 4481
rect 1732 4447 1738 4481
rect 1692 4409 1738 4447
rect 1692 4375 1698 4409
rect 1732 4375 1738 4409
rect 1692 4328 1738 4375
rect 1850 4525 1896 4528
rect 1941 4525 1986 4591
rect 1850 4481 1986 4525
rect 1850 4447 1856 4481
rect 1890 4480 1986 4481
rect 2024 4481 2070 4528
rect 1890 4447 1896 4480
rect 1850 4409 1896 4447
rect 2024 4447 2030 4481
rect 2064 4447 2070 4481
rect 2024 4412 2070 4447
rect 1998 4410 2070 4412
rect 1850 4375 1856 4409
rect 1890 4375 1896 4409
rect 1850 4328 1896 4375
rect 1928 4409 2070 4410
rect 1928 4385 2030 4409
rect 1928 4368 1935 4385
rect 1929 4333 1935 4368
rect 1987 4375 2030 4385
rect 2064 4375 2070 4409
rect 1987 4368 2070 4375
rect 1987 4333 1993 4368
rect 2024 4328 2070 4368
rect 2182 4484 2228 4528
rect 2366 4484 2412 4528
rect 2182 4481 2412 4484
rect 2182 4447 2188 4481
rect 2222 4447 2372 4481
rect 2406 4447 2412 4481
rect 2182 4409 2412 4447
rect 2182 4375 2188 4409
rect 2222 4375 2372 4409
rect 2406 4375 2412 4409
rect 2182 4358 2412 4375
rect 2182 4328 2228 4358
rect 2366 4328 2412 4358
rect 2524 4481 2570 4528
rect 2524 4447 2530 4481
rect 2564 4447 2570 4481
rect 2642 4457 2687 4591
rect 3118 4628 3511 4667
rect 3724 4690 4264 4734
rect 3724 4638 3776 4690
rect 3828 4681 3840 4690
rect 3892 4681 3904 4690
rect 3956 4681 3968 4690
rect 4020 4681 4032 4690
rect 4084 4681 4096 4690
rect 4148 4681 4160 4690
rect 3831 4647 3840 4681
rect 3903 4647 3904 4681
rect 4084 4647 4085 4681
rect 4148 4647 4157 4681
rect 3828 4638 3840 4647
rect 3892 4638 3904 4647
rect 3956 4638 3968 4647
rect 4020 4638 4032 4647
rect 4084 4638 4096 4647
rect 4148 4638 4160 4647
rect 4212 4638 4264 4690
rect 2774 4584 2816 4585
rect 2758 4576 2816 4584
rect 2758 4524 2769 4576
rect 2821 4524 2827 4576
rect 3118 4528 3157 4628
rect 3724 4594 4264 4638
rect 3741 4538 3787 4594
rect 3736 4537 3787 4538
rect 2758 4481 2816 4524
rect 2524 4409 2570 4447
rect 2524 4375 2530 4409
rect 2564 4375 2570 4409
rect 2524 4368 2570 4375
rect 2613 4429 2715 4457
rect 2613 4395 2647 4429
rect 2681 4395 2715 4429
rect 2524 4328 2574 4368
rect 2613 4367 2715 4395
rect 2758 4447 2776 4481
rect 2810 4447 2816 4481
rect 2758 4409 2816 4447
rect 2758 4375 2776 4409
rect 2810 4375 2816 4409
rect 1008 4268 1052 4322
rect 1245 4287 1328 4306
rect 852 4224 1052 4268
rect 1148 4285 1328 4287
rect 1148 4233 1155 4285
rect 1207 4275 1328 4285
rect 1207 4241 1269 4275
rect 1303 4241 1328 4275
rect 1207 4233 1328 4241
rect 1148 4232 1328 4233
rect 852 4102 896 4224
rect 1245 4211 1328 4232
rect 1568 4294 1602 4328
rect 1568 4284 1820 4294
rect 1568 4232 1758 4284
rect 1810 4232 1820 4284
rect 1568 4222 1820 4232
rect 1568 4190 1608 4222
rect 1853 4190 1892 4328
rect 2185 4190 2224 4328
rect 2255 4291 2325 4297
rect 2255 4282 2331 4291
rect 2255 4230 2270 4282
rect 2322 4230 2331 4282
rect 2255 4221 2331 4230
rect 2255 4215 2325 4221
rect 2368 4190 2407 4328
rect 2530 4294 2574 4328
rect 2758 4328 2816 4375
rect 2928 4481 2974 4528
rect 2928 4447 2934 4481
rect 2968 4468 2974 4481
rect 3114 4481 3160 4528
rect 3114 4468 3120 4481
rect 2968 4447 3120 4468
rect 3154 4447 3160 4481
rect 3272 4481 3318 4528
rect 3272 4471 3278 4481
rect 3312 4471 3318 4481
rect 3736 4491 3782 4537
rect 2928 4409 3160 4447
rect 3262 4419 3268 4471
rect 3320 4419 3326 4471
rect 3736 4457 3742 4491
rect 3776 4457 3782 4491
rect 3736 4419 3782 4457
rect 2928 4375 2934 4409
rect 2968 4375 3120 4409
rect 3154 4375 3160 4409
rect 2928 4358 3160 4375
rect 2928 4328 2974 4358
rect 3114 4328 3160 4358
rect 3272 4409 3318 4419
rect 3272 4375 3278 4409
rect 3312 4375 3318 4409
rect 3272 4328 3318 4375
rect 3736 4385 3742 4419
rect 3776 4385 3782 4419
rect 3736 4338 3782 4385
rect 3894 4491 3940 4538
rect 3894 4457 3900 4491
rect 3934 4457 3940 4491
rect 3894 4419 3940 4457
rect 3894 4385 3900 4419
rect 3934 4385 3940 4419
rect 3894 4338 3940 4385
rect 4044 4491 4090 4594
rect 4558 4538 4597 4744
rect 4738 4738 4744 4744
rect 4796 4738 4802 4790
rect 4868 4538 4907 4825
rect 5081 4831 7015 4861
rect 5029 4814 5081 4820
rect 6862 4783 6868 4790
rect 6516 4744 6868 4783
rect 5682 4690 6222 4734
rect 5682 4638 5734 4690
rect 5786 4680 5798 4690
rect 5850 4680 5862 4690
rect 5914 4680 5926 4690
rect 5978 4680 5990 4690
rect 6042 4680 6054 4690
rect 6106 4680 6118 4690
rect 5790 4646 5798 4680
rect 6042 4646 6044 4680
rect 6106 4646 6116 4680
rect 5786 4638 5798 4646
rect 5850 4638 5862 4646
rect 5914 4638 5926 4646
rect 5978 4638 5990 4646
rect 6042 4638 6054 4646
rect 6106 4638 6118 4646
rect 6170 4638 6222 4690
rect 5682 4594 6222 4638
rect 5700 4538 5746 4594
rect 4044 4457 4050 4491
rect 4084 4457 4090 4491
rect 4044 4419 4090 4457
rect 4044 4385 4050 4419
rect 4084 4385 4090 4419
rect 4044 4338 4090 4385
rect 4202 4491 4248 4538
rect 4202 4457 4208 4491
rect 4242 4457 4248 4491
rect 4396 4491 4442 4538
rect 4396 4465 4402 4491
rect 4202 4419 4248 4457
rect 4202 4385 4208 4419
rect 4242 4385 4248 4419
rect 4285 4463 4402 4465
rect 4285 4411 4292 4463
rect 4344 4457 4402 4463
rect 4436 4457 4442 4491
rect 4344 4419 4442 4457
rect 4344 4411 4402 4419
rect 4285 4410 4402 4411
rect 4202 4338 4248 4385
rect 4396 4385 4402 4410
rect 4436 4385 4442 4419
rect 4396 4338 4442 4385
rect 4554 4491 4600 4538
rect 4554 4457 4560 4491
rect 4594 4458 4600 4491
rect 4704 4491 4750 4538
rect 4704 4458 4710 4491
rect 4594 4457 4710 4458
rect 4744 4457 4750 4491
rect 4554 4419 4750 4457
rect 4554 4385 4560 4419
rect 4594 4392 4710 4419
rect 4594 4385 4600 4392
rect 4554 4338 4600 4385
rect 4704 4385 4710 4392
rect 4744 4385 4750 4419
rect 4704 4338 4750 4385
rect 4862 4491 4908 4538
rect 4862 4457 4868 4491
rect 4902 4457 4908 4491
rect 5694 4492 5740 4538
rect 5027 4462 5057 4471
rect 4862 4419 4908 4457
rect 4862 4385 4868 4419
rect 4902 4385 4908 4419
rect 5010 4410 5016 4462
rect 5068 4410 5074 4462
rect 5694 4458 5700 4492
rect 5734 4458 5740 4492
rect 5694 4420 5740 4458
rect 4862 4338 4908 4385
rect 5026 4369 5057 4410
rect 5694 4386 5700 4420
rect 5734 4386 5740 4420
rect 2758 4294 2802 4328
rect 2530 4250 2656 4294
rect 1242 4170 1248 4174
rect 1138 4126 1248 4170
rect 1138 4102 1182 4126
rect 1242 4122 1248 4126
rect 1300 4122 1306 4174
rect 1404 4157 1450 4190
rect 1404 4123 1410 4157
rect 1444 4123 1450 4157
rect 1404 4119 1450 4123
rect 378 4074 434 4080
rect 550 4074 622 4096
rect 434 4068 622 4074
rect 434 4028 565 4068
rect 606 4028 622 4068
rect 434 4018 622 4028
rect 378 4012 434 4018
rect 550 3998 622 4018
rect 696 4068 768 4096
rect 696 4028 712 4068
rect 753 4028 768 4068
rect 696 3998 768 4028
rect 840 4073 912 4102
rect 840 4033 856 4073
rect 897 4033 912 4073
rect 840 4004 912 4033
rect 994 4074 1182 4102
rect 994 4034 1010 4074
rect 1051 4058 1182 4074
rect 1399 4090 1450 4119
rect 1562 4157 1608 4190
rect 1562 4123 1568 4157
rect 1602 4123 1608 4157
rect 1692 4157 1738 4190
rect 1692 4128 1698 4157
rect 1562 4090 1608 4123
rect 1690 4123 1698 4128
rect 1732 4128 1738 4157
rect 1850 4157 1896 4190
rect 2024 4174 2070 4190
rect 1732 4123 1740 4128
rect 1051 4034 1066 4058
rect 1399 4044 1449 4090
rect 1690 4044 1740 4123
rect 1850 4123 1856 4157
rect 1890 4123 1896 4157
rect 1850 4090 1896 4123
rect 2014 4122 2020 4174
rect 2072 4122 2078 4174
rect 2182 4157 2228 4190
rect 2182 4123 2188 4157
rect 2222 4123 2228 4157
rect 2024 4090 2070 4122
rect 2182 4090 2228 4123
rect 2366 4157 2412 4190
rect 2524 4172 2570 4190
rect 2366 4123 2372 4157
rect 2406 4123 2412 4157
rect 2366 4090 2412 4123
rect 2516 4120 2522 4172
rect 2574 4120 2580 4172
rect 2524 4090 2570 4120
rect 2024 4058 2068 4090
rect 2612 4058 2656 4250
rect 994 4004 1066 4034
rect 1324 3989 1960 4044
rect 2024 4014 2656 4058
rect 2694 4250 2802 4294
rect 2832 4280 2904 4290
rect 2694 4052 2738 4250
rect 2832 4228 2842 4280
rect 2894 4228 2904 4280
rect 2832 4218 2904 4228
rect 2933 4190 2972 4328
rect 3118 4190 3157 4328
rect 3272 4284 3316 4328
rect 3268 4278 3320 4284
rect 3555 4253 3561 4305
rect 3613 4298 3619 4305
rect 3662 4298 3713 4310
rect 3613 4295 3713 4298
rect 3613 4261 3670 4295
rect 3704 4261 3713 4295
rect 3613 4259 3713 4261
rect 3613 4253 3619 4259
rect 3662 4247 3713 4259
rect 3897 4289 3936 4338
rect 3976 4296 4027 4301
rect 3970 4289 3976 4296
rect 3897 4250 3976 4289
rect 3268 4220 3320 4226
rect 3897 4200 3936 4250
rect 3970 4244 3976 4250
rect 4028 4244 4034 4296
rect 4206 4282 4245 4338
rect 4300 4282 4347 4293
rect 4206 4280 4347 4282
rect 4206 4247 4306 4280
rect 3976 4238 4027 4244
rect 4206 4200 4245 4247
rect 4300 4246 4306 4247
rect 4340 4246 4347 4280
rect 4300 4234 4347 4246
rect 2766 4184 2818 4190
rect 2766 4126 2776 4132
rect 2770 4123 2776 4126
rect 2810 4126 2818 4132
rect 2928 4157 2974 4190
rect 2810 4123 2816 4126
rect 2770 4090 2816 4123
rect 2928 4123 2934 4157
rect 2968 4123 2974 4157
rect 2928 4090 2974 4123
rect 3114 4157 3160 4190
rect 3114 4123 3120 4157
rect 3154 4123 3160 4157
rect 3114 4090 3160 4123
rect 3272 4157 3318 4190
rect 3272 4123 3278 4157
rect 3312 4123 3318 4157
rect 3272 4090 3318 4123
rect 3274 4052 3318 4090
rect 2694 4008 3318 4052
rect 3736 4167 3782 4200
rect 3736 4133 3742 4167
rect 3776 4133 3782 4167
rect 3736 4100 3782 4133
rect 3894 4167 3940 4200
rect 3894 4133 3900 4167
rect 3934 4133 3940 4167
rect 4044 4167 4090 4200
rect 4044 4138 4050 4167
rect 3894 4100 3940 4133
rect 4042 4133 4050 4138
rect 4084 4133 4090 4167
rect 4042 4100 4090 4133
rect 4202 4167 4248 4200
rect 4202 4133 4208 4167
rect 4242 4133 4248 4167
rect 4202 4100 4248 4133
rect 3736 4044 3780 4100
rect 4042 4044 4089 4100
rect 1324 3937 1360 3989
rect 1412 3937 1424 3989
rect 1476 3980 1488 3989
rect 1540 3980 1552 3989
rect 1604 3980 1616 3989
rect 1668 3980 1680 3989
rect 1732 3980 1744 3989
rect 1796 3980 1808 3989
rect 1479 3946 1488 3980
rect 1551 3946 1552 3980
rect 1732 3946 1733 3980
rect 1796 3946 1805 3980
rect 1476 3937 1488 3946
rect 1540 3937 1552 3946
rect 1604 3937 1616 3946
rect 1668 3937 1680 3946
rect 1732 3937 1744 3946
rect 1796 3937 1808 3946
rect 1860 3937 1872 3989
rect 1924 3937 1960 3989
rect 3704 4000 4244 4044
rect 3704 3991 3756 4000
rect 3808 3991 3820 4000
rect 1324 3904 1960 3937
rect 2346 3959 2426 3984
rect 2346 3955 3517 3959
rect 2346 3921 2369 3955
rect 2403 3921 3517 3955
rect 2346 3917 3517 3921
rect 2346 3892 2426 3917
rect 2636 3859 2702 3871
rect 272 3805 278 3859
rect 332 3805 2642 3859
rect 2696 3805 2702 3859
rect 2636 3793 2702 3805
rect 3475 3764 3517 3917
rect 3704 3957 3741 3991
rect 3808 3957 3813 3991
rect 3704 3948 3756 3957
rect 3808 3948 3820 3957
rect 3872 3948 3884 4000
rect 3936 3948 3948 4000
rect 4000 3948 4012 4000
rect 4064 3948 4076 4000
rect 4128 3991 4140 4000
rect 4192 3991 4244 4000
rect 4135 3957 4140 3991
rect 4207 3957 4244 3991
rect 4128 3948 4140 3957
rect 4192 3948 4244 3957
rect 3704 3904 4244 3948
rect 3559 3799 3565 3851
rect 3617 3844 3623 3851
rect 4306 3844 4345 4234
rect 4558 4202 4597 4338
rect 4628 4307 4680 4313
rect 4625 4258 4628 4304
rect 4680 4258 4683 4304
rect 4875 4262 4904 4338
rect 4628 4249 4680 4255
rect 4875 4234 4980 4262
rect 4396 4169 4442 4202
rect 4396 4135 4402 4169
rect 4436 4135 4442 4169
rect 4396 4102 4442 4135
rect 4554 4182 4600 4202
rect 4704 4182 4750 4202
rect 4862 4182 4908 4202
rect 4554 4169 4750 4182
rect 4554 4135 4560 4169
rect 4594 4135 4710 4169
rect 4744 4135 4750 4169
rect 4554 4116 4750 4135
rect 4856 4130 4862 4182
rect 4914 4130 4920 4182
rect 4554 4102 4600 4116
rect 4704 4102 4750 4116
rect 4862 4102 4908 4130
rect 4402 3952 4430 4102
rect 4558 4057 4597 4102
rect 4552 4051 4604 4057
rect 4552 3993 4604 3999
rect 4952 3952 4980 4234
rect 5026 4184 5056 4369
rect 5694 4338 5740 4386
rect 5852 4492 5898 4538
rect 5852 4458 5858 4492
rect 5892 4458 5898 4492
rect 5852 4420 5898 4458
rect 5852 4386 5858 4420
rect 5892 4386 5898 4420
rect 5852 4338 5898 4386
rect 6002 4492 6048 4594
rect 6516 4538 6556 4744
rect 6862 4738 6868 4744
rect 6920 4738 6926 4790
rect 6985 4778 7015 4831
rect 6985 4749 7016 4778
rect 6002 4458 6008 4492
rect 6042 4458 6048 4492
rect 6002 4420 6048 4458
rect 6002 4386 6008 4420
rect 6042 4386 6048 4420
rect 6002 4338 6048 4386
rect 6160 4492 6206 4538
rect 6160 4458 6166 4492
rect 6200 4458 6206 4492
rect 6354 4492 6400 4538
rect 6354 4466 6360 4492
rect 6160 4420 6206 4458
rect 6160 4386 6166 4420
rect 6200 4386 6206 4420
rect 6244 4464 6360 4466
rect 6244 4412 6250 4464
rect 6302 4458 6360 4464
rect 6394 4458 6400 4492
rect 6302 4420 6400 4458
rect 6302 4412 6360 4420
rect 6244 4410 6360 4412
rect 6160 4338 6206 4386
rect 6354 4386 6360 4410
rect 6394 4386 6400 4420
rect 6354 4338 6400 4386
rect 6512 4492 6558 4538
rect 6512 4458 6518 4492
rect 6552 4458 6558 4492
rect 6662 4492 6708 4538
rect 6662 4458 6668 4492
rect 6702 4458 6708 4492
rect 6512 4420 6708 4458
rect 6512 4386 6518 4420
rect 6552 4392 6668 4420
rect 6552 4386 6558 4392
rect 6512 4338 6558 4386
rect 6662 4386 6668 4392
rect 6702 4386 6708 4420
rect 6662 4338 6708 4386
rect 6820 4492 6866 4538
rect 6820 4458 6826 4492
rect 6860 4458 6866 4492
rect 6986 4462 7016 4749
rect 6820 4420 6866 4458
rect 6820 4386 6826 4420
rect 6860 4386 6866 4420
rect 6968 4410 6974 4462
rect 7026 4410 7032 4462
rect 6820 4338 6866 4386
rect 6984 4370 7016 4410
rect 5111 4253 5117 4305
rect 5169 4298 5175 4305
rect 5620 4298 5672 4310
rect 5169 4296 5672 4298
rect 5169 4262 5628 4296
rect 5662 4262 5672 4296
rect 5169 4259 5672 4262
rect 5169 4253 5175 4259
rect 5620 4248 5672 4259
rect 5856 4290 5894 4338
rect 5934 4296 5986 4302
rect 5928 4290 5934 4296
rect 5856 4250 5934 4290
rect 5856 4200 5894 4250
rect 5928 4244 5934 4250
rect 5986 4244 5992 4296
rect 6164 4282 6204 4338
rect 6258 4282 6306 4294
rect 6164 4280 6306 4282
rect 6164 4248 6264 4280
rect 5934 4238 5986 4244
rect 6164 4200 6204 4248
rect 6258 4246 6264 4248
rect 6298 4246 6306 4280
rect 6258 4234 6306 4246
rect 5009 4132 5015 4184
rect 5067 4132 5073 4184
rect 5694 4168 5740 4200
rect 5694 4134 5700 4168
rect 5734 4134 5740 4168
rect 4402 3924 4980 3952
rect 3617 3805 4345 3844
rect 3617 3799 3623 3805
rect 5021 3764 5063 4132
rect 5694 4100 5740 4134
rect 5852 4168 5898 4200
rect 5852 4134 5858 4168
rect 5892 4134 5898 4168
rect 6002 4168 6048 4200
rect 6002 4138 6008 4168
rect 5852 4100 5898 4134
rect 6000 4134 6008 4138
rect 6042 4134 6048 4168
rect 5694 4044 5738 4100
rect 6000 4044 6048 4134
rect 6160 4168 6206 4200
rect 6160 4134 6166 4168
rect 6200 4134 6206 4168
rect 6160 4100 6206 4134
rect 5662 4000 6202 4044
rect 5662 3992 5714 4000
rect 5766 3992 5778 4000
rect 5662 3958 5700 3992
rect 5766 3958 5772 3992
rect 5662 3948 5714 3958
rect 5766 3948 5778 3958
rect 5830 3948 5842 4000
rect 5894 3948 5906 4000
rect 5958 3948 5970 4000
rect 6022 3948 6034 4000
rect 6086 3992 6098 4000
rect 6150 3992 6202 4000
rect 6094 3958 6098 3992
rect 6166 3958 6202 3992
rect 6086 3948 6098 3958
rect 6150 3948 6202 3958
rect 5662 3904 6202 3948
rect 5111 3799 5117 3851
rect 5169 3844 5175 3851
rect 6264 3844 6304 4234
rect 6516 4202 6556 4338
rect 6586 4308 6638 4314
rect 6584 4258 6586 4304
rect 6638 4258 6642 4304
rect 6834 4262 6862 4338
rect 6586 4250 6638 4256
rect 6834 4234 6936 4262
rect 6354 4170 6400 4202
rect 6354 4136 6360 4170
rect 6394 4136 6400 4170
rect 6354 4102 6400 4136
rect 6512 4182 6558 4202
rect 6662 4182 6708 4202
rect 6820 4182 6866 4202
rect 6512 4170 6708 4182
rect 6512 4136 6518 4170
rect 6552 4136 6668 4170
rect 6702 4136 6708 4170
rect 6512 4116 6708 4136
rect 6814 4130 6820 4182
rect 6872 4130 6878 4182
rect 6512 4102 6558 4116
rect 6662 4102 6708 4116
rect 6820 4102 6866 4130
rect 6360 3952 6388 4102
rect 6516 4058 6556 4102
rect 6510 4052 6562 4058
rect 6510 3994 6562 4000
rect 6908 3952 6936 4234
rect 6984 4184 7014 4370
rect 6968 4132 6974 4184
rect 7026 4132 7032 4184
rect 6360 3924 6936 3952
rect 6908 3860 6936 3924
rect 5169 3806 6304 3844
rect 6346 3832 6936 3860
rect 5169 3805 5572 3806
rect 5169 3799 5175 3805
rect 3475 3722 5063 3764
rect 5035 3681 5087 3687
rect 3472 3597 4907 3636
rect 6346 3669 6374 3832
rect 6908 3830 6936 3832
rect 6512 3766 6564 3772
rect 6512 3708 6564 3714
rect 5087 3641 6374 3669
rect 6523 3651 6553 3708
rect 5035 3623 5087 3629
rect 6523 3621 7015 3651
rect 1348 3463 1880 3506
rect 1348 3454 1398 3463
rect 1450 3454 1462 3463
rect 1348 3420 1383 3454
rect 1450 3420 1455 3454
rect 1348 3411 1398 3420
rect 1450 3411 1462 3420
rect 1514 3411 1526 3463
rect 1578 3411 1590 3463
rect 1642 3411 1654 3463
rect 1706 3411 1718 3463
rect 1770 3454 1782 3463
rect 1834 3454 1880 3463
rect 1777 3420 1782 3454
rect 1849 3420 1880 3454
rect 3472 3439 3511 3597
rect 4738 3555 4744 3562
rect 4558 3516 4744 3555
rect 1770 3411 1782 3420
rect 1834 3411 1880 3420
rect 550 3392 622 3396
rect 550 3340 560 3392
rect 612 3340 622 3392
rect 696 3390 768 3396
rect 550 3328 566 3340
rect 607 3328 622 3340
rect 682 3388 768 3390
rect 682 3336 702 3388
rect 754 3336 768 3388
rect 682 3334 710 3336
rect 550 3298 622 3328
rect 696 3328 710 3334
rect 751 3328 768 3336
rect 696 3298 768 3328
rect 840 3373 912 3402
rect 840 3333 856 3373
rect 897 3333 912 3373
rect 840 3304 912 3333
rect 994 3373 1066 3402
rect 994 3333 1009 3373
rect 1050 3333 1066 3373
rect 1348 3366 1880 3411
rect 994 3304 1066 3333
rect 564 3258 608 3298
rect 856 3238 900 3304
rect 378 3230 433 3236
rect 846 3186 852 3238
rect 904 3186 910 3238
rect 378 2945 433 3175
rect 856 3146 900 3186
rect 1008 3146 1052 3304
rect 1407 3300 1448 3366
rect 1693 3300 1735 3366
rect 1941 3363 2687 3408
rect 1404 3253 1450 3300
rect 1404 3219 1410 3253
rect 1444 3219 1450 3253
rect 1404 3181 1450 3219
rect 1404 3147 1410 3181
rect 1444 3147 1450 3181
rect 708 3102 900 3146
rect 372 2890 378 2945
rect 433 2890 439 2945
rect 708 2868 752 3102
rect 998 3094 1004 3146
rect 1056 3094 1062 3146
rect 1404 3100 1450 3147
rect 1562 3253 1608 3300
rect 1562 3219 1568 3253
rect 1602 3219 1608 3253
rect 1562 3181 1608 3219
rect 1562 3147 1568 3181
rect 1602 3147 1608 3181
rect 1562 3100 1608 3147
rect 1692 3253 1738 3300
rect 1692 3219 1698 3253
rect 1732 3219 1738 3253
rect 1692 3181 1738 3219
rect 1692 3147 1698 3181
rect 1732 3147 1738 3181
rect 1692 3100 1738 3147
rect 1850 3297 1896 3300
rect 1941 3297 1986 3363
rect 1850 3253 1986 3297
rect 1850 3219 1856 3253
rect 1890 3252 1986 3253
rect 2024 3253 2070 3300
rect 1890 3219 1896 3252
rect 1850 3181 1896 3219
rect 2024 3219 2030 3253
rect 2064 3219 2070 3253
rect 2024 3184 2070 3219
rect 1998 3182 2070 3184
rect 1850 3147 1856 3181
rect 1890 3147 1896 3181
rect 1850 3100 1896 3147
rect 1928 3181 2070 3182
rect 1928 3157 2030 3181
rect 1928 3140 1935 3157
rect 1929 3105 1935 3140
rect 1987 3147 2030 3157
rect 2064 3147 2070 3181
rect 1987 3140 2070 3147
rect 1987 3105 1993 3140
rect 2024 3100 2070 3140
rect 2182 3256 2228 3300
rect 2366 3256 2412 3300
rect 2182 3253 2412 3256
rect 2182 3219 2188 3253
rect 2222 3219 2372 3253
rect 2406 3219 2412 3253
rect 2182 3181 2412 3219
rect 2182 3147 2188 3181
rect 2222 3147 2372 3181
rect 2406 3147 2412 3181
rect 2182 3130 2412 3147
rect 2182 3100 2228 3130
rect 2366 3100 2412 3130
rect 2524 3253 2570 3300
rect 2524 3219 2530 3253
rect 2564 3219 2570 3253
rect 2642 3229 2687 3363
rect 3118 3400 3511 3439
rect 3724 3462 4264 3506
rect 3724 3410 3776 3462
rect 3828 3453 3840 3462
rect 3892 3453 3904 3462
rect 3956 3453 3968 3462
rect 4020 3453 4032 3462
rect 4084 3453 4096 3462
rect 4148 3453 4160 3462
rect 3831 3419 3840 3453
rect 3903 3419 3904 3453
rect 4084 3419 4085 3453
rect 4148 3419 4157 3453
rect 3828 3410 3840 3419
rect 3892 3410 3904 3419
rect 3956 3410 3968 3419
rect 4020 3410 4032 3419
rect 4084 3410 4096 3419
rect 4148 3410 4160 3419
rect 4212 3410 4264 3462
rect 2774 3356 2816 3357
rect 2758 3348 2816 3356
rect 2758 3296 2769 3348
rect 2821 3296 2827 3348
rect 3118 3300 3157 3400
rect 3724 3366 4264 3410
rect 3741 3310 3787 3366
rect 3736 3309 3787 3310
rect 2758 3253 2816 3296
rect 2524 3181 2570 3219
rect 2524 3147 2530 3181
rect 2564 3147 2570 3181
rect 2524 3140 2570 3147
rect 2613 3201 2715 3229
rect 2613 3167 2647 3201
rect 2681 3167 2715 3201
rect 2524 3100 2574 3140
rect 2613 3139 2715 3167
rect 2758 3219 2776 3253
rect 2810 3219 2816 3253
rect 2758 3181 2816 3219
rect 2758 3147 2776 3181
rect 2810 3147 2816 3181
rect 1008 3040 1052 3094
rect 1245 3059 1328 3078
rect 852 2996 1052 3040
rect 1148 3057 1328 3059
rect 1148 3005 1155 3057
rect 1207 3047 1328 3057
rect 1207 3013 1269 3047
rect 1303 3013 1328 3047
rect 1207 3005 1328 3013
rect 1148 3004 1328 3005
rect 852 2874 896 2996
rect 1245 2983 1328 3004
rect 1568 3066 1602 3100
rect 1568 3056 1820 3066
rect 1568 3004 1758 3056
rect 1810 3004 1820 3056
rect 1568 2994 1820 3004
rect 1568 2962 1608 2994
rect 1853 2962 1892 3100
rect 2185 2962 2224 3100
rect 2255 3063 2325 3069
rect 2255 3054 2331 3063
rect 2255 3002 2270 3054
rect 2322 3002 2331 3054
rect 2255 2993 2331 3002
rect 2255 2987 2325 2993
rect 2368 2962 2407 3100
rect 2530 3066 2574 3100
rect 2758 3100 2816 3147
rect 2928 3253 2974 3300
rect 2928 3219 2934 3253
rect 2968 3240 2974 3253
rect 3114 3253 3160 3300
rect 3114 3240 3120 3253
rect 2968 3219 3120 3240
rect 3154 3219 3160 3253
rect 3272 3253 3318 3300
rect 3272 3243 3278 3253
rect 3312 3243 3318 3253
rect 3736 3263 3782 3309
rect 2928 3181 3160 3219
rect 3262 3191 3268 3243
rect 3320 3191 3326 3243
rect 3736 3229 3742 3263
rect 3776 3229 3782 3263
rect 3736 3191 3782 3229
rect 2928 3147 2934 3181
rect 2968 3147 3120 3181
rect 3154 3147 3160 3181
rect 2928 3130 3160 3147
rect 2928 3100 2974 3130
rect 3114 3100 3160 3130
rect 3272 3181 3318 3191
rect 3272 3147 3278 3181
rect 3312 3147 3318 3181
rect 3272 3100 3318 3147
rect 3736 3157 3742 3191
rect 3776 3157 3782 3191
rect 3736 3110 3782 3157
rect 3894 3263 3940 3310
rect 3894 3229 3900 3263
rect 3934 3229 3940 3263
rect 3894 3191 3940 3229
rect 3894 3157 3900 3191
rect 3934 3157 3940 3191
rect 3894 3110 3940 3157
rect 4044 3263 4090 3366
rect 4558 3310 4597 3516
rect 4738 3510 4744 3516
rect 4796 3510 4802 3562
rect 4868 3310 4907 3597
rect 6837 3555 6843 3562
rect 6516 3516 6843 3555
rect 5682 3462 6222 3506
rect 5682 3410 5734 3462
rect 5786 3452 5798 3462
rect 5850 3452 5862 3462
rect 5914 3452 5926 3462
rect 5978 3452 5990 3462
rect 6042 3452 6054 3462
rect 6106 3452 6118 3462
rect 5790 3418 5798 3452
rect 6042 3418 6044 3452
rect 6106 3418 6116 3452
rect 5786 3410 5798 3418
rect 5850 3410 5862 3418
rect 5914 3410 5926 3418
rect 5978 3410 5990 3418
rect 6042 3410 6054 3418
rect 6106 3410 6118 3418
rect 6170 3410 6222 3462
rect 5682 3366 6222 3410
rect 5700 3310 5746 3366
rect 4044 3229 4050 3263
rect 4084 3229 4090 3263
rect 4044 3191 4090 3229
rect 4044 3157 4050 3191
rect 4084 3157 4090 3191
rect 4044 3110 4090 3157
rect 4202 3263 4248 3310
rect 4202 3229 4208 3263
rect 4242 3229 4248 3263
rect 4396 3263 4442 3310
rect 4396 3237 4402 3263
rect 4202 3191 4248 3229
rect 4202 3157 4208 3191
rect 4242 3157 4248 3191
rect 4285 3235 4402 3237
rect 4285 3183 4292 3235
rect 4344 3229 4402 3235
rect 4436 3229 4442 3263
rect 4344 3191 4442 3229
rect 4344 3183 4402 3191
rect 4285 3182 4402 3183
rect 4202 3110 4248 3157
rect 4396 3157 4402 3182
rect 4436 3157 4442 3191
rect 4396 3110 4442 3157
rect 4554 3263 4600 3310
rect 4554 3229 4560 3263
rect 4594 3230 4600 3263
rect 4704 3263 4750 3310
rect 4704 3230 4710 3263
rect 4594 3229 4710 3230
rect 4744 3229 4750 3263
rect 4554 3191 4750 3229
rect 4554 3157 4560 3191
rect 4594 3164 4710 3191
rect 4594 3157 4600 3164
rect 4554 3110 4600 3157
rect 4704 3157 4710 3164
rect 4744 3157 4750 3191
rect 4704 3110 4750 3157
rect 4862 3263 4908 3310
rect 4862 3229 4868 3263
rect 4902 3229 4908 3263
rect 5694 3264 5740 3310
rect 5027 3234 5057 3243
rect 4862 3191 4908 3229
rect 4862 3157 4868 3191
rect 4902 3157 4908 3191
rect 5010 3182 5016 3234
rect 5068 3182 5074 3234
rect 5694 3230 5700 3264
rect 5734 3230 5740 3264
rect 5694 3192 5740 3230
rect 4862 3110 4908 3157
rect 5026 3141 5057 3182
rect 5694 3158 5700 3192
rect 5734 3158 5740 3192
rect 2758 3066 2802 3100
rect 2530 3022 2656 3066
rect 1242 2942 1248 2946
rect 1138 2898 1248 2942
rect 1138 2874 1182 2898
rect 1242 2894 1248 2898
rect 1300 2894 1306 2946
rect 1404 2929 1450 2962
rect 1404 2895 1410 2929
rect 1444 2895 1450 2929
rect 1404 2891 1450 2895
rect 378 2846 434 2852
rect 550 2846 622 2868
rect 434 2840 622 2846
rect 434 2800 565 2840
rect 606 2800 622 2840
rect 434 2790 622 2800
rect 378 2784 434 2790
rect 550 2770 622 2790
rect 696 2840 768 2868
rect 696 2800 712 2840
rect 753 2800 768 2840
rect 696 2770 768 2800
rect 840 2845 912 2874
rect 840 2805 856 2845
rect 897 2805 912 2845
rect 840 2776 912 2805
rect 994 2846 1182 2874
rect 994 2806 1010 2846
rect 1051 2830 1182 2846
rect 1399 2862 1450 2891
rect 1562 2929 1608 2962
rect 1562 2895 1568 2929
rect 1602 2895 1608 2929
rect 1692 2929 1738 2962
rect 1692 2900 1698 2929
rect 1562 2862 1608 2895
rect 1690 2895 1698 2900
rect 1732 2900 1738 2929
rect 1850 2929 1896 2962
rect 2024 2946 2070 2962
rect 1732 2895 1740 2900
rect 1051 2806 1066 2830
rect 1399 2816 1449 2862
rect 1690 2816 1740 2895
rect 1850 2895 1856 2929
rect 1890 2895 1896 2929
rect 1850 2862 1896 2895
rect 2014 2894 2020 2946
rect 2072 2894 2078 2946
rect 2182 2929 2228 2962
rect 2182 2895 2188 2929
rect 2222 2895 2228 2929
rect 2024 2862 2070 2894
rect 2182 2862 2228 2895
rect 2366 2929 2412 2962
rect 2524 2944 2570 2962
rect 2366 2895 2372 2929
rect 2406 2895 2412 2929
rect 2366 2862 2412 2895
rect 2516 2892 2522 2944
rect 2574 2892 2580 2944
rect 2524 2862 2570 2892
rect 2024 2830 2068 2862
rect 2612 2830 2656 3022
rect 994 2776 1066 2806
rect 1324 2761 1960 2816
rect 2024 2786 2656 2830
rect 2694 3022 2802 3066
rect 2832 3052 2904 3062
rect 2694 2824 2738 3022
rect 2832 3000 2842 3052
rect 2894 3000 2904 3052
rect 2832 2990 2904 3000
rect 2933 2962 2972 3100
rect 3118 2962 3157 3100
rect 3272 3056 3316 3100
rect 3268 3050 3320 3056
rect 3555 3025 3561 3077
rect 3613 3070 3619 3077
rect 3662 3070 3713 3082
rect 3613 3067 3713 3070
rect 3613 3033 3670 3067
rect 3704 3033 3713 3067
rect 3613 3031 3713 3033
rect 3613 3025 3619 3031
rect 3662 3019 3713 3031
rect 3897 3061 3936 3110
rect 3976 3068 4027 3073
rect 3970 3061 3976 3068
rect 3897 3022 3976 3061
rect 3268 2992 3320 2998
rect 3897 2972 3936 3022
rect 3970 3016 3976 3022
rect 4028 3016 4034 3068
rect 4206 3054 4245 3110
rect 4300 3054 4347 3065
rect 4206 3052 4347 3054
rect 4206 3019 4306 3052
rect 3976 3010 4027 3016
rect 4206 2972 4245 3019
rect 4300 3018 4306 3019
rect 4340 3018 4347 3052
rect 4300 3006 4347 3018
rect 2766 2956 2818 2962
rect 2766 2898 2776 2904
rect 2770 2895 2776 2898
rect 2810 2898 2818 2904
rect 2928 2929 2974 2962
rect 2810 2895 2816 2898
rect 2770 2862 2816 2895
rect 2928 2895 2934 2929
rect 2968 2895 2974 2929
rect 2928 2862 2974 2895
rect 3114 2929 3160 2962
rect 3114 2895 3120 2929
rect 3154 2895 3160 2929
rect 3114 2862 3160 2895
rect 3272 2929 3318 2962
rect 3272 2895 3278 2929
rect 3312 2895 3318 2929
rect 3272 2862 3318 2895
rect 3274 2824 3318 2862
rect 2694 2780 3318 2824
rect 3736 2939 3782 2972
rect 3736 2905 3742 2939
rect 3776 2905 3782 2939
rect 3736 2872 3782 2905
rect 3894 2939 3940 2972
rect 3894 2905 3900 2939
rect 3934 2905 3940 2939
rect 4044 2939 4090 2972
rect 4044 2910 4050 2939
rect 3894 2872 3940 2905
rect 4042 2905 4050 2910
rect 4084 2905 4090 2939
rect 4042 2872 4090 2905
rect 4202 2939 4248 2972
rect 4202 2905 4208 2939
rect 4242 2905 4248 2939
rect 4202 2872 4248 2905
rect 3736 2816 3780 2872
rect 4042 2816 4089 2872
rect 1324 2709 1360 2761
rect 1412 2709 1424 2761
rect 1476 2752 1488 2761
rect 1540 2752 1552 2761
rect 1604 2752 1616 2761
rect 1668 2752 1680 2761
rect 1732 2752 1744 2761
rect 1796 2752 1808 2761
rect 1479 2718 1488 2752
rect 1551 2718 1552 2752
rect 1732 2718 1733 2752
rect 1796 2718 1805 2752
rect 1476 2709 1488 2718
rect 1540 2709 1552 2718
rect 1604 2709 1616 2718
rect 1668 2709 1680 2718
rect 1732 2709 1744 2718
rect 1796 2709 1808 2718
rect 1860 2709 1872 2761
rect 1924 2709 1960 2761
rect 3704 2772 4244 2816
rect 3704 2763 3756 2772
rect 3808 2763 3820 2772
rect 1324 2676 1960 2709
rect 2346 2731 2426 2756
rect 2346 2727 3517 2731
rect 2346 2693 2369 2727
rect 2403 2693 3517 2727
rect 2346 2689 3517 2693
rect 2346 2664 2426 2689
rect 2636 2631 2702 2643
rect 272 2577 278 2631
rect 332 2577 2642 2631
rect 2696 2577 2702 2631
rect 2636 2565 2702 2577
rect 3475 2536 3517 2689
rect 3704 2729 3741 2763
rect 3808 2729 3813 2763
rect 3704 2720 3756 2729
rect 3808 2720 3820 2729
rect 3872 2720 3884 2772
rect 3936 2720 3948 2772
rect 4000 2720 4012 2772
rect 4064 2720 4076 2772
rect 4128 2763 4140 2772
rect 4192 2763 4244 2772
rect 4135 2729 4140 2763
rect 4207 2729 4244 2763
rect 4128 2720 4140 2729
rect 4192 2720 4244 2729
rect 3704 2676 4244 2720
rect 3559 2571 3565 2623
rect 3617 2616 3623 2623
rect 4306 2616 4345 3006
rect 4558 2974 4597 3110
rect 4628 3079 4680 3085
rect 4625 3030 4628 3076
rect 4680 3030 4683 3076
rect 4875 3034 4904 3110
rect 4628 3021 4680 3027
rect 4875 3006 4980 3034
rect 4396 2941 4442 2974
rect 4396 2907 4402 2941
rect 4436 2907 4442 2941
rect 4396 2874 4442 2907
rect 4554 2954 4600 2974
rect 4704 2954 4750 2974
rect 4862 2954 4908 2974
rect 4554 2941 4750 2954
rect 4554 2907 4560 2941
rect 4594 2907 4710 2941
rect 4744 2907 4750 2941
rect 4554 2888 4750 2907
rect 4856 2902 4862 2954
rect 4914 2902 4920 2954
rect 4554 2874 4600 2888
rect 4704 2874 4750 2888
rect 4862 2874 4908 2902
rect 4402 2724 4430 2874
rect 4558 2829 4597 2874
rect 4552 2823 4604 2829
rect 4552 2765 4604 2771
rect 4952 2724 4980 3006
rect 5026 2956 5056 3141
rect 5694 3110 5740 3158
rect 5852 3264 5898 3310
rect 5852 3230 5858 3264
rect 5892 3230 5898 3264
rect 5852 3192 5898 3230
rect 5852 3158 5858 3192
rect 5892 3158 5898 3192
rect 5852 3110 5898 3158
rect 6002 3264 6048 3366
rect 6516 3310 6556 3516
rect 6837 3510 6843 3516
rect 6895 3510 6901 3562
rect 6985 3550 7015 3621
rect 6985 3521 7016 3550
rect 6002 3230 6008 3264
rect 6042 3230 6048 3264
rect 6002 3192 6048 3230
rect 6002 3158 6008 3192
rect 6042 3158 6048 3192
rect 6002 3110 6048 3158
rect 6160 3264 6206 3310
rect 6160 3230 6166 3264
rect 6200 3230 6206 3264
rect 6354 3264 6400 3310
rect 6354 3238 6360 3264
rect 6160 3192 6206 3230
rect 6160 3158 6166 3192
rect 6200 3158 6206 3192
rect 6244 3236 6360 3238
rect 6244 3184 6250 3236
rect 6302 3230 6360 3236
rect 6394 3230 6400 3264
rect 6302 3192 6400 3230
rect 6302 3184 6360 3192
rect 6244 3182 6360 3184
rect 6160 3110 6206 3158
rect 6354 3158 6360 3182
rect 6394 3158 6400 3192
rect 6354 3110 6400 3158
rect 6512 3264 6558 3310
rect 6512 3230 6518 3264
rect 6552 3230 6558 3264
rect 6662 3264 6708 3310
rect 6662 3230 6668 3264
rect 6702 3230 6708 3264
rect 6512 3192 6708 3230
rect 6512 3158 6518 3192
rect 6552 3164 6668 3192
rect 6552 3158 6558 3164
rect 6512 3110 6558 3158
rect 6662 3158 6668 3164
rect 6702 3158 6708 3192
rect 6662 3110 6708 3158
rect 6820 3264 6866 3310
rect 6820 3230 6826 3264
rect 6860 3230 6866 3264
rect 6986 3234 7016 3521
rect 6820 3192 6866 3230
rect 6820 3158 6826 3192
rect 6860 3158 6866 3192
rect 6968 3182 6974 3234
rect 7026 3182 7032 3234
rect 6820 3110 6866 3158
rect 6984 3142 7016 3182
rect 5191 3025 5197 3077
rect 5249 3070 5255 3077
rect 5620 3070 5672 3082
rect 5249 3068 5672 3070
rect 5249 3034 5628 3068
rect 5662 3034 5672 3068
rect 5249 3031 5672 3034
rect 5249 3025 5255 3031
rect 5620 3020 5672 3031
rect 5856 3062 5894 3110
rect 5934 3068 5986 3074
rect 5928 3062 5934 3068
rect 5856 3022 5934 3062
rect 5856 2972 5894 3022
rect 5928 3016 5934 3022
rect 5986 3016 5992 3068
rect 6164 3054 6204 3110
rect 6258 3054 6306 3066
rect 6164 3052 6306 3054
rect 6164 3020 6264 3052
rect 5934 3010 5986 3016
rect 6164 2972 6204 3020
rect 6258 3018 6264 3020
rect 6298 3018 6306 3052
rect 6258 3006 6306 3018
rect 5009 2904 5015 2956
rect 5067 2904 5073 2956
rect 5694 2940 5740 2972
rect 5694 2906 5700 2940
rect 5734 2906 5740 2940
rect 4402 2696 4980 2724
rect 3617 2577 4345 2616
rect 3617 2571 3623 2577
rect 5021 2536 5063 2904
rect 5694 2872 5740 2906
rect 5852 2940 5898 2972
rect 5852 2906 5858 2940
rect 5892 2906 5898 2940
rect 6002 2940 6048 2972
rect 6002 2910 6008 2940
rect 5852 2872 5898 2906
rect 6000 2906 6008 2910
rect 6042 2906 6048 2940
rect 5694 2816 5738 2872
rect 6000 2816 6048 2906
rect 6160 2940 6206 2972
rect 6160 2906 6166 2940
rect 6200 2906 6206 2940
rect 6160 2872 6206 2906
rect 5662 2772 6202 2816
rect 5662 2764 5714 2772
rect 5766 2764 5778 2772
rect 5662 2730 5700 2764
rect 5766 2730 5772 2764
rect 5662 2720 5714 2730
rect 5766 2720 5778 2730
rect 5830 2720 5842 2772
rect 5894 2720 5906 2772
rect 5958 2720 5970 2772
rect 6022 2720 6034 2772
rect 6086 2764 6098 2772
rect 6150 2764 6202 2772
rect 6094 2730 6098 2764
rect 6166 2730 6202 2764
rect 6086 2720 6098 2730
rect 6150 2720 6202 2730
rect 5662 2676 6202 2720
rect 5191 2571 5197 2623
rect 5249 2616 5255 2623
rect 6264 2616 6304 3006
rect 6516 2974 6556 3110
rect 6586 3080 6638 3086
rect 6584 3030 6586 3076
rect 6638 3030 6642 3076
rect 6834 3034 6862 3110
rect 6586 3022 6638 3028
rect 6834 3006 6936 3034
rect 6354 2942 6400 2974
rect 6354 2908 6360 2942
rect 6394 2908 6400 2942
rect 6354 2874 6400 2908
rect 6512 2954 6558 2974
rect 6662 2954 6708 2974
rect 6820 2954 6866 2974
rect 6512 2942 6708 2954
rect 6512 2908 6518 2942
rect 6552 2908 6668 2942
rect 6702 2908 6708 2942
rect 6512 2888 6708 2908
rect 6814 2902 6820 2954
rect 6872 2902 6878 2954
rect 6512 2874 6558 2888
rect 6662 2874 6708 2888
rect 6820 2874 6866 2902
rect 6360 2724 6388 2874
rect 6516 2830 6556 2874
rect 6510 2824 6562 2830
rect 6510 2766 6562 2772
rect 6908 2724 6936 3006
rect 6984 2956 7014 3142
rect 6968 2904 6974 2956
rect 7026 2904 7032 2956
rect 6360 2696 6936 2724
rect 5249 2578 6304 2616
rect 5249 2577 5587 2578
rect 5249 2571 5255 2577
rect 3475 2494 5063 2536
rect 6908 2524 6936 2696
rect 7107 2536 7159 2542
rect 6908 2496 7107 2524
rect 7107 2478 7159 2484
rect 5029 2416 5081 2422
rect 3472 2369 4907 2408
rect 1348 2235 1880 2278
rect 1348 2226 1398 2235
rect 1450 2226 1462 2235
rect 1348 2192 1383 2226
rect 1450 2192 1455 2226
rect 1348 2183 1398 2192
rect 1450 2183 1462 2192
rect 1514 2183 1526 2235
rect 1578 2183 1590 2235
rect 1642 2183 1654 2235
rect 1706 2183 1718 2235
rect 1770 2226 1782 2235
rect 1834 2226 1880 2235
rect 1777 2192 1782 2226
rect 1849 2192 1880 2226
rect 3472 2211 3511 2369
rect 4738 2327 4744 2334
rect 4558 2288 4744 2327
rect 1770 2183 1782 2192
rect 1834 2183 1880 2192
rect 550 2164 622 2168
rect 550 2112 560 2164
rect 612 2112 622 2164
rect 696 2162 768 2168
rect 550 2100 566 2112
rect 607 2100 622 2112
rect 682 2160 768 2162
rect 682 2108 702 2160
rect 754 2108 768 2160
rect 682 2106 710 2108
rect 550 2070 622 2100
rect 696 2100 710 2106
rect 751 2100 768 2108
rect 696 2070 768 2100
rect 840 2145 912 2174
rect 840 2105 856 2145
rect 897 2105 912 2145
rect 840 2076 912 2105
rect 994 2145 1066 2174
rect 994 2105 1009 2145
rect 1050 2105 1066 2145
rect 1348 2138 1880 2183
rect 994 2076 1066 2105
rect 564 2030 608 2070
rect 856 2010 900 2076
rect 378 2002 433 2008
rect 846 1958 852 2010
rect 904 1958 910 2010
rect 378 1717 433 1947
rect 856 1918 900 1958
rect 1008 1918 1052 2076
rect 1407 2072 1448 2138
rect 1693 2072 1735 2138
rect 1941 2135 2687 2180
rect 1404 2025 1450 2072
rect 1404 1991 1410 2025
rect 1444 1991 1450 2025
rect 1404 1953 1450 1991
rect 1404 1919 1410 1953
rect 1444 1919 1450 1953
rect 708 1874 900 1918
rect 372 1662 378 1717
rect 433 1662 439 1717
rect 708 1640 752 1874
rect 998 1866 1004 1918
rect 1056 1866 1062 1918
rect 1404 1872 1450 1919
rect 1562 2025 1608 2072
rect 1562 1991 1568 2025
rect 1602 1991 1608 2025
rect 1562 1953 1608 1991
rect 1562 1919 1568 1953
rect 1602 1919 1608 1953
rect 1562 1872 1608 1919
rect 1692 2025 1738 2072
rect 1692 1991 1698 2025
rect 1732 1991 1738 2025
rect 1692 1953 1738 1991
rect 1692 1919 1698 1953
rect 1732 1919 1738 1953
rect 1692 1872 1738 1919
rect 1850 2069 1896 2072
rect 1941 2069 1986 2135
rect 1850 2025 1986 2069
rect 1850 1991 1856 2025
rect 1890 2024 1986 2025
rect 2024 2025 2070 2072
rect 1890 1991 1896 2024
rect 1850 1953 1896 1991
rect 2024 1991 2030 2025
rect 2064 1991 2070 2025
rect 2024 1956 2070 1991
rect 1998 1954 2070 1956
rect 1850 1919 1856 1953
rect 1890 1919 1896 1953
rect 1850 1872 1896 1919
rect 1928 1953 2070 1954
rect 1928 1929 2030 1953
rect 1928 1912 1935 1929
rect 1929 1877 1935 1912
rect 1987 1919 2030 1929
rect 2064 1919 2070 1953
rect 1987 1912 2070 1919
rect 1987 1877 1993 1912
rect 2024 1872 2070 1912
rect 2182 2028 2228 2072
rect 2366 2028 2412 2072
rect 2182 2025 2412 2028
rect 2182 1991 2188 2025
rect 2222 1991 2372 2025
rect 2406 1991 2412 2025
rect 2182 1953 2412 1991
rect 2182 1919 2188 1953
rect 2222 1919 2372 1953
rect 2406 1919 2412 1953
rect 2182 1902 2412 1919
rect 2182 1872 2228 1902
rect 2366 1872 2412 1902
rect 2524 2025 2570 2072
rect 2524 1991 2530 2025
rect 2564 1991 2570 2025
rect 2642 2001 2687 2135
rect 3118 2172 3511 2211
rect 3724 2234 4264 2278
rect 3724 2182 3776 2234
rect 3828 2225 3840 2234
rect 3892 2225 3904 2234
rect 3956 2225 3968 2234
rect 4020 2225 4032 2234
rect 4084 2225 4096 2234
rect 4148 2225 4160 2234
rect 3831 2191 3840 2225
rect 3903 2191 3904 2225
rect 4084 2191 4085 2225
rect 4148 2191 4157 2225
rect 3828 2182 3840 2191
rect 3892 2182 3904 2191
rect 3956 2182 3968 2191
rect 4020 2182 4032 2191
rect 4084 2182 4096 2191
rect 4148 2182 4160 2191
rect 4212 2182 4264 2234
rect 2774 2128 2816 2129
rect 2758 2120 2816 2128
rect 2758 2068 2769 2120
rect 2821 2068 2827 2120
rect 3118 2072 3157 2172
rect 3724 2138 4264 2182
rect 3741 2082 3787 2138
rect 3736 2081 3787 2082
rect 2758 2025 2816 2068
rect 2524 1953 2570 1991
rect 2524 1919 2530 1953
rect 2564 1919 2570 1953
rect 2524 1912 2570 1919
rect 2613 1973 2715 2001
rect 2613 1939 2647 1973
rect 2681 1939 2715 1973
rect 2524 1872 2574 1912
rect 2613 1911 2715 1939
rect 2758 1991 2776 2025
rect 2810 1991 2816 2025
rect 2758 1953 2816 1991
rect 2758 1919 2776 1953
rect 2810 1919 2816 1953
rect 1008 1812 1052 1866
rect 1245 1831 1328 1850
rect 852 1768 1052 1812
rect 1148 1829 1328 1831
rect 1148 1777 1155 1829
rect 1207 1819 1328 1829
rect 1207 1785 1269 1819
rect 1303 1785 1328 1819
rect 1207 1777 1328 1785
rect 1148 1776 1328 1777
rect 852 1646 896 1768
rect 1245 1755 1328 1776
rect 1568 1838 1602 1872
rect 1568 1828 1820 1838
rect 1568 1776 1758 1828
rect 1810 1776 1820 1828
rect 1568 1766 1820 1776
rect 1568 1734 1608 1766
rect 1853 1734 1892 1872
rect 2185 1734 2224 1872
rect 2255 1835 2325 1841
rect 2255 1826 2331 1835
rect 2255 1774 2270 1826
rect 2322 1774 2331 1826
rect 2255 1765 2331 1774
rect 2255 1759 2325 1765
rect 2368 1734 2407 1872
rect 2530 1838 2574 1872
rect 2758 1872 2816 1919
rect 2928 2025 2974 2072
rect 2928 1991 2934 2025
rect 2968 2012 2974 2025
rect 3114 2025 3160 2072
rect 3114 2012 3120 2025
rect 2968 1991 3120 2012
rect 3154 1991 3160 2025
rect 3272 2025 3318 2072
rect 3272 2015 3278 2025
rect 3312 2015 3318 2025
rect 3736 2035 3782 2081
rect 2928 1953 3160 1991
rect 3262 1963 3268 2015
rect 3320 1963 3326 2015
rect 3736 2001 3742 2035
rect 3776 2001 3782 2035
rect 3736 1963 3782 2001
rect 2928 1919 2934 1953
rect 2968 1919 3120 1953
rect 3154 1919 3160 1953
rect 2928 1902 3160 1919
rect 2928 1872 2974 1902
rect 3114 1872 3160 1902
rect 3272 1953 3318 1963
rect 3272 1919 3278 1953
rect 3312 1919 3318 1953
rect 3272 1872 3318 1919
rect 3736 1929 3742 1963
rect 3776 1929 3782 1963
rect 3736 1882 3782 1929
rect 3894 2035 3940 2082
rect 3894 2001 3900 2035
rect 3934 2001 3940 2035
rect 3894 1963 3940 2001
rect 3894 1929 3900 1963
rect 3934 1929 3940 1963
rect 3894 1882 3940 1929
rect 4044 2035 4090 2138
rect 4558 2082 4597 2288
rect 4738 2282 4744 2288
rect 4796 2282 4802 2334
rect 4868 2082 4907 2369
rect 5081 2375 7015 2405
rect 5029 2358 5081 2364
rect 6862 2327 6868 2334
rect 6516 2288 6868 2327
rect 5682 2234 6222 2278
rect 5682 2182 5734 2234
rect 5786 2224 5798 2234
rect 5850 2224 5862 2234
rect 5914 2224 5926 2234
rect 5978 2224 5990 2234
rect 6042 2224 6054 2234
rect 6106 2224 6118 2234
rect 5790 2190 5798 2224
rect 6042 2190 6044 2224
rect 6106 2190 6116 2224
rect 5786 2182 5798 2190
rect 5850 2182 5862 2190
rect 5914 2182 5926 2190
rect 5978 2182 5990 2190
rect 6042 2182 6054 2190
rect 6106 2182 6118 2190
rect 6170 2182 6222 2234
rect 5682 2138 6222 2182
rect 5700 2082 5746 2138
rect 4044 2001 4050 2035
rect 4084 2001 4090 2035
rect 4044 1963 4090 2001
rect 4044 1929 4050 1963
rect 4084 1929 4090 1963
rect 4044 1882 4090 1929
rect 4202 2035 4248 2082
rect 4202 2001 4208 2035
rect 4242 2001 4248 2035
rect 4396 2035 4442 2082
rect 4396 2009 4402 2035
rect 4202 1963 4248 2001
rect 4202 1929 4208 1963
rect 4242 1929 4248 1963
rect 4285 2007 4402 2009
rect 4285 1955 4292 2007
rect 4344 2001 4402 2007
rect 4436 2001 4442 2035
rect 4344 1963 4442 2001
rect 4344 1955 4402 1963
rect 4285 1954 4402 1955
rect 4202 1882 4248 1929
rect 4396 1929 4402 1954
rect 4436 1929 4442 1963
rect 4396 1882 4442 1929
rect 4554 2035 4600 2082
rect 4554 2001 4560 2035
rect 4594 2002 4600 2035
rect 4704 2035 4750 2082
rect 4704 2002 4710 2035
rect 4594 2001 4710 2002
rect 4744 2001 4750 2035
rect 4554 1963 4750 2001
rect 4554 1929 4560 1963
rect 4594 1936 4710 1963
rect 4594 1929 4600 1936
rect 4554 1882 4600 1929
rect 4704 1929 4710 1936
rect 4744 1929 4750 1963
rect 4704 1882 4750 1929
rect 4862 2035 4908 2082
rect 4862 2001 4868 2035
rect 4902 2001 4908 2035
rect 5694 2036 5740 2082
rect 5027 2006 5057 2015
rect 4862 1963 4908 2001
rect 4862 1929 4868 1963
rect 4902 1929 4908 1963
rect 5010 1954 5016 2006
rect 5068 1954 5074 2006
rect 5694 2002 5700 2036
rect 5734 2002 5740 2036
rect 5694 1964 5740 2002
rect 4862 1882 4908 1929
rect 5026 1913 5057 1954
rect 5694 1930 5700 1964
rect 5734 1930 5740 1964
rect 2758 1838 2802 1872
rect 2530 1794 2656 1838
rect 1242 1714 1248 1718
rect 1138 1670 1248 1714
rect 1138 1646 1182 1670
rect 1242 1666 1248 1670
rect 1300 1666 1306 1718
rect 1404 1701 1450 1734
rect 1404 1667 1410 1701
rect 1444 1667 1450 1701
rect 1404 1663 1450 1667
rect 378 1618 434 1624
rect 550 1618 622 1640
rect 434 1612 622 1618
rect 434 1572 565 1612
rect 606 1572 622 1612
rect 434 1562 622 1572
rect 378 1556 434 1562
rect 550 1542 622 1562
rect 696 1612 768 1640
rect 696 1572 712 1612
rect 753 1572 768 1612
rect 696 1542 768 1572
rect 840 1617 912 1646
rect 840 1577 856 1617
rect 897 1577 912 1617
rect 840 1548 912 1577
rect 994 1618 1182 1646
rect 994 1578 1010 1618
rect 1051 1602 1182 1618
rect 1399 1634 1450 1663
rect 1562 1701 1608 1734
rect 1562 1667 1568 1701
rect 1602 1667 1608 1701
rect 1692 1701 1738 1734
rect 1692 1672 1698 1701
rect 1562 1634 1608 1667
rect 1690 1667 1698 1672
rect 1732 1672 1738 1701
rect 1850 1701 1896 1734
rect 2024 1718 2070 1734
rect 1732 1667 1740 1672
rect 1051 1578 1066 1602
rect 1399 1588 1449 1634
rect 1690 1588 1740 1667
rect 1850 1667 1856 1701
rect 1890 1667 1896 1701
rect 1850 1634 1896 1667
rect 2014 1666 2020 1718
rect 2072 1666 2078 1718
rect 2182 1701 2228 1734
rect 2182 1667 2188 1701
rect 2222 1667 2228 1701
rect 2024 1634 2070 1666
rect 2182 1634 2228 1667
rect 2366 1701 2412 1734
rect 2524 1716 2570 1734
rect 2366 1667 2372 1701
rect 2406 1667 2412 1701
rect 2366 1634 2412 1667
rect 2516 1664 2522 1716
rect 2574 1664 2580 1716
rect 2524 1634 2570 1664
rect 2024 1602 2068 1634
rect 2612 1602 2656 1794
rect 994 1548 1066 1578
rect 1324 1533 1960 1588
rect 2024 1558 2656 1602
rect 2694 1794 2802 1838
rect 2832 1824 2904 1834
rect 2694 1596 2738 1794
rect 2832 1772 2842 1824
rect 2894 1772 2904 1824
rect 2832 1762 2904 1772
rect 2933 1734 2972 1872
rect 3118 1734 3157 1872
rect 3272 1828 3316 1872
rect 3268 1822 3320 1828
rect 3555 1797 3561 1849
rect 3613 1842 3619 1849
rect 3662 1842 3713 1854
rect 3613 1839 3713 1842
rect 3613 1805 3670 1839
rect 3704 1805 3713 1839
rect 3613 1803 3713 1805
rect 3613 1797 3619 1803
rect 3662 1791 3713 1803
rect 3897 1833 3936 1882
rect 3976 1840 4027 1845
rect 3970 1833 3976 1840
rect 3897 1794 3976 1833
rect 3268 1764 3320 1770
rect 3897 1744 3936 1794
rect 3970 1788 3976 1794
rect 4028 1788 4034 1840
rect 4206 1826 4245 1882
rect 4300 1826 4347 1837
rect 4206 1824 4347 1826
rect 4206 1791 4306 1824
rect 3976 1782 4027 1788
rect 4206 1744 4245 1791
rect 4300 1790 4306 1791
rect 4340 1790 4347 1824
rect 4300 1778 4347 1790
rect 2766 1728 2818 1734
rect 2766 1670 2776 1676
rect 2770 1667 2776 1670
rect 2810 1670 2818 1676
rect 2928 1701 2974 1734
rect 2810 1667 2816 1670
rect 2770 1634 2816 1667
rect 2928 1667 2934 1701
rect 2968 1667 2974 1701
rect 2928 1634 2974 1667
rect 3114 1701 3160 1734
rect 3114 1667 3120 1701
rect 3154 1667 3160 1701
rect 3114 1634 3160 1667
rect 3272 1701 3318 1734
rect 3272 1667 3278 1701
rect 3312 1667 3318 1701
rect 3272 1634 3318 1667
rect 3274 1596 3318 1634
rect 2694 1552 3318 1596
rect 3736 1711 3782 1744
rect 3736 1677 3742 1711
rect 3776 1677 3782 1711
rect 3736 1644 3782 1677
rect 3894 1711 3940 1744
rect 3894 1677 3900 1711
rect 3934 1677 3940 1711
rect 4044 1711 4090 1744
rect 4044 1682 4050 1711
rect 3894 1644 3940 1677
rect 4042 1677 4050 1682
rect 4084 1677 4090 1711
rect 4042 1644 4090 1677
rect 4202 1711 4248 1744
rect 4202 1677 4208 1711
rect 4242 1677 4248 1711
rect 4202 1644 4248 1677
rect 3736 1588 3780 1644
rect 4042 1588 4089 1644
rect 1324 1481 1360 1533
rect 1412 1481 1424 1533
rect 1476 1524 1488 1533
rect 1540 1524 1552 1533
rect 1604 1524 1616 1533
rect 1668 1524 1680 1533
rect 1732 1524 1744 1533
rect 1796 1524 1808 1533
rect 1479 1490 1488 1524
rect 1551 1490 1552 1524
rect 1732 1490 1733 1524
rect 1796 1490 1805 1524
rect 1476 1481 1488 1490
rect 1540 1481 1552 1490
rect 1604 1481 1616 1490
rect 1668 1481 1680 1490
rect 1732 1481 1744 1490
rect 1796 1481 1808 1490
rect 1860 1481 1872 1533
rect 1924 1481 1960 1533
rect 3704 1544 4244 1588
rect 3704 1535 3756 1544
rect 3808 1535 3820 1544
rect 1324 1448 1960 1481
rect 2346 1503 2426 1528
rect 2346 1499 3517 1503
rect 2346 1465 2369 1499
rect 2403 1465 3517 1499
rect 2346 1461 3517 1465
rect 2346 1436 2426 1461
rect 2636 1403 2702 1415
rect 272 1349 278 1403
rect 332 1349 2642 1403
rect 2696 1349 2702 1403
rect 2636 1337 2702 1349
rect 3475 1308 3517 1461
rect 3704 1501 3741 1535
rect 3808 1501 3813 1535
rect 3704 1492 3756 1501
rect 3808 1492 3820 1501
rect 3872 1492 3884 1544
rect 3936 1492 3948 1544
rect 4000 1492 4012 1544
rect 4064 1492 4076 1544
rect 4128 1535 4140 1544
rect 4192 1535 4244 1544
rect 4135 1501 4140 1535
rect 4207 1501 4244 1535
rect 4128 1492 4140 1501
rect 4192 1492 4244 1501
rect 3704 1448 4244 1492
rect 3559 1343 3565 1395
rect 3617 1388 3623 1395
rect 4306 1388 4345 1778
rect 4558 1746 4597 1882
rect 4628 1851 4680 1857
rect 4625 1802 4628 1848
rect 4680 1802 4683 1848
rect 4875 1806 4904 1882
rect 4628 1793 4680 1799
rect 4875 1778 4980 1806
rect 4396 1713 4442 1746
rect 4396 1679 4402 1713
rect 4436 1679 4442 1713
rect 4396 1646 4442 1679
rect 4554 1726 4600 1746
rect 4704 1726 4750 1746
rect 4862 1726 4908 1746
rect 4554 1713 4750 1726
rect 4554 1679 4560 1713
rect 4594 1679 4710 1713
rect 4744 1679 4750 1713
rect 4554 1660 4750 1679
rect 4856 1674 4862 1726
rect 4914 1674 4920 1726
rect 4554 1646 4600 1660
rect 4704 1646 4750 1660
rect 4862 1646 4908 1674
rect 4402 1496 4430 1646
rect 4558 1601 4597 1646
rect 4552 1595 4604 1601
rect 4552 1537 4604 1543
rect 4952 1496 4980 1778
rect 5026 1728 5056 1913
rect 5694 1882 5740 1930
rect 5852 2036 5898 2082
rect 5852 2002 5858 2036
rect 5892 2002 5898 2036
rect 5852 1964 5898 2002
rect 5852 1930 5858 1964
rect 5892 1930 5898 1964
rect 5852 1882 5898 1930
rect 6002 2036 6048 2138
rect 6516 2082 6556 2288
rect 6862 2282 6868 2288
rect 6920 2282 6926 2334
rect 6985 2322 7015 2375
rect 6985 2293 7016 2322
rect 6002 2002 6008 2036
rect 6042 2002 6048 2036
rect 6002 1964 6048 2002
rect 6002 1930 6008 1964
rect 6042 1930 6048 1964
rect 6002 1882 6048 1930
rect 6160 2036 6206 2082
rect 6160 2002 6166 2036
rect 6200 2002 6206 2036
rect 6354 2036 6400 2082
rect 6354 2010 6360 2036
rect 6160 1964 6206 2002
rect 6160 1930 6166 1964
rect 6200 1930 6206 1964
rect 6244 2008 6360 2010
rect 6244 1956 6250 2008
rect 6302 2002 6360 2008
rect 6394 2002 6400 2036
rect 6302 1964 6400 2002
rect 6302 1956 6360 1964
rect 6244 1954 6360 1956
rect 6160 1882 6206 1930
rect 6354 1930 6360 1954
rect 6394 1930 6400 1964
rect 6354 1882 6400 1930
rect 6512 2036 6558 2082
rect 6512 2002 6518 2036
rect 6552 2002 6558 2036
rect 6662 2036 6708 2082
rect 6662 2002 6668 2036
rect 6702 2002 6708 2036
rect 6512 1964 6708 2002
rect 6512 1930 6518 1964
rect 6552 1936 6668 1964
rect 6552 1930 6558 1936
rect 6512 1882 6558 1930
rect 6662 1930 6668 1936
rect 6702 1930 6708 1964
rect 6662 1882 6708 1930
rect 6820 2036 6866 2082
rect 6820 2002 6826 2036
rect 6860 2002 6866 2036
rect 6986 2006 7016 2293
rect 6820 1964 6866 2002
rect 6820 1930 6826 1964
rect 6860 1930 6866 1964
rect 6968 1954 6974 2006
rect 7026 1954 7032 2006
rect 6820 1882 6866 1930
rect 6984 1914 7016 1954
rect 5111 1797 5117 1849
rect 5169 1842 5175 1849
rect 5620 1842 5672 1854
rect 5169 1840 5672 1842
rect 5169 1806 5628 1840
rect 5662 1806 5672 1840
rect 5169 1803 5672 1806
rect 5169 1797 5175 1803
rect 5620 1792 5672 1803
rect 5856 1834 5894 1882
rect 5934 1840 5986 1846
rect 5928 1834 5934 1840
rect 5856 1794 5934 1834
rect 5856 1744 5894 1794
rect 5928 1788 5934 1794
rect 5986 1788 5992 1840
rect 6164 1826 6204 1882
rect 6258 1826 6306 1838
rect 6164 1824 6306 1826
rect 6164 1792 6264 1824
rect 5934 1782 5986 1788
rect 6164 1744 6204 1792
rect 6258 1790 6264 1792
rect 6298 1790 6306 1824
rect 6258 1778 6306 1790
rect 5009 1676 5015 1728
rect 5067 1676 5073 1728
rect 5694 1712 5740 1744
rect 5694 1678 5700 1712
rect 5734 1678 5740 1712
rect 4402 1468 4980 1496
rect 3617 1349 4345 1388
rect 3617 1343 3623 1349
rect 5021 1308 5063 1676
rect 5694 1644 5740 1678
rect 5852 1712 5898 1744
rect 5852 1678 5858 1712
rect 5892 1678 5898 1712
rect 6002 1712 6048 1744
rect 6002 1682 6008 1712
rect 5852 1644 5898 1678
rect 6000 1678 6008 1682
rect 6042 1678 6048 1712
rect 5694 1588 5738 1644
rect 6000 1588 6048 1678
rect 6160 1712 6206 1744
rect 6160 1678 6166 1712
rect 6200 1678 6206 1712
rect 6160 1644 6206 1678
rect 5662 1544 6202 1588
rect 5662 1536 5714 1544
rect 5766 1536 5778 1544
rect 5662 1502 5700 1536
rect 5766 1502 5772 1536
rect 5662 1492 5714 1502
rect 5766 1492 5778 1502
rect 5830 1492 5842 1544
rect 5894 1492 5906 1544
rect 5958 1492 5970 1544
rect 6022 1492 6034 1544
rect 6086 1536 6098 1544
rect 6150 1536 6202 1544
rect 6094 1502 6098 1536
rect 6166 1502 6202 1536
rect 6086 1492 6098 1502
rect 6150 1492 6202 1502
rect 5662 1448 6202 1492
rect 5111 1343 5117 1395
rect 5169 1388 5175 1395
rect 6264 1388 6304 1778
rect 6516 1746 6556 1882
rect 6586 1852 6638 1858
rect 6584 1802 6586 1848
rect 6638 1802 6642 1848
rect 6834 1806 6862 1882
rect 6586 1794 6638 1800
rect 6834 1778 6936 1806
rect 6354 1714 6400 1746
rect 6354 1680 6360 1714
rect 6394 1680 6400 1714
rect 6354 1646 6400 1680
rect 6512 1726 6558 1746
rect 6662 1726 6708 1746
rect 6820 1726 6866 1746
rect 6512 1714 6708 1726
rect 6512 1680 6518 1714
rect 6552 1680 6668 1714
rect 6702 1680 6708 1714
rect 6512 1660 6708 1680
rect 6814 1674 6820 1726
rect 6872 1674 6878 1726
rect 6512 1646 6558 1660
rect 6662 1646 6708 1660
rect 6820 1646 6866 1674
rect 6360 1496 6388 1646
rect 6516 1602 6556 1646
rect 6510 1596 6562 1602
rect 6510 1538 6562 1544
rect 6908 1496 6936 1778
rect 6984 1728 7014 1914
rect 6968 1676 6974 1728
rect 7026 1676 7032 1728
rect 6360 1468 6936 1496
rect 6908 1404 6936 1468
rect 5169 1350 6304 1388
rect 6346 1376 6936 1404
rect 5169 1349 5572 1350
rect 5169 1343 5175 1349
rect 3475 1266 5063 1308
rect 5035 1225 5087 1231
rect 3472 1141 4907 1180
rect 6346 1213 6374 1376
rect 6908 1374 6936 1376
rect 5087 1185 6374 1213
rect 5035 1167 5087 1173
rect 1348 1007 1880 1050
rect 1348 998 1398 1007
rect 1450 998 1462 1007
rect 1348 964 1383 998
rect 1450 964 1455 998
rect 1348 955 1398 964
rect 1450 955 1462 964
rect 1514 955 1526 1007
rect 1578 955 1590 1007
rect 1642 955 1654 1007
rect 1706 955 1718 1007
rect 1770 998 1782 1007
rect 1834 998 1880 1007
rect 1777 964 1782 998
rect 1849 964 1880 998
rect 3472 983 3511 1141
rect 4738 1099 4744 1106
rect 4558 1060 4744 1099
rect 1770 955 1782 964
rect 1834 955 1880 964
rect 550 936 622 940
rect 550 884 560 936
rect 612 884 622 936
rect 696 934 768 940
rect 550 872 566 884
rect 607 872 622 884
rect 682 932 768 934
rect 682 880 702 932
rect 754 880 768 932
rect 682 878 710 880
rect 550 842 622 872
rect 696 872 710 878
rect 751 872 768 880
rect 696 842 768 872
rect 840 917 912 946
rect 840 877 856 917
rect 897 877 912 917
rect 840 848 912 877
rect 994 917 1066 946
rect 994 877 1009 917
rect 1050 877 1066 917
rect 1348 910 1880 955
rect 994 848 1066 877
rect 564 802 608 842
rect 856 782 900 848
rect 378 774 433 780
rect 846 730 852 782
rect 904 730 910 782
rect 378 489 433 719
rect 856 690 900 730
rect 1008 690 1052 848
rect 1407 844 1448 910
rect 1693 844 1735 910
rect 1941 907 2687 952
rect 1404 797 1450 844
rect 1404 763 1410 797
rect 1444 763 1450 797
rect 1404 725 1450 763
rect 1404 691 1410 725
rect 1444 691 1450 725
rect 708 646 900 690
rect 372 434 378 489
rect 433 434 439 489
rect 708 412 752 646
rect 998 638 1004 690
rect 1056 638 1062 690
rect 1404 644 1450 691
rect 1562 797 1608 844
rect 1562 763 1568 797
rect 1602 763 1608 797
rect 1562 725 1608 763
rect 1562 691 1568 725
rect 1602 691 1608 725
rect 1562 644 1608 691
rect 1692 797 1738 844
rect 1692 763 1698 797
rect 1732 763 1738 797
rect 1692 725 1738 763
rect 1692 691 1698 725
rect 1732 691 1738 725
rect 1692 644 1738 691
rect 1850 841 1896 844
rect 1941 841 1986 907
rect 1850 797 1986 841
rect 1850 763 1856 797
rect 1890 796 1986 797
rect 2024 797 2070 844
rect 1890 763 1896 796
rect 1850 725 1896 763
rect 2024 763 2030 797
rect 2064 763 2070 797
rect 2024 728 2070 763
rect 1998 726 2070 728
rect 1850 691 1856 725
rect 1890 691 1896 725
rect 1850 644 1896 691
rect 1928 725 2070 726
rect 1928 701 2030 725
rect 1928 684 1935 701
rect 1929 649 1935 684
rect 1987 691 2030 701
rect 2064 691 2070 725
rect 1987 684 2070 691
rect 1987 649 1993 684
rect 2024 644 2070 684
rect 2182 800 2228 844
rect 2366 800 2412 844
rect 2182 797 2412 800
rect 2182 763 2188 797
rect 2222 763 2372 797
rect 2406 763 2412 797
rect 2182 725 2412 763
rect 2182 691 2188 725
rect 2222 691 2372 725
rect 2406 691 2412 725
rect 2182 674 2412 691
rect 2182 644 2228 674
rect 2366 644 2412 674
rect 2524 797 2570 844
rect 2524 763 2530 797
rect 2564 763 2570 797
rect 2642 773 2687 907
rect 3118 944 3511 983
rect 3724 1006 4264 1050
rect 3724 954 3776 1006
rect 3828 997 3840 1006
rect 3892 997 3904 1006
rect 3956 997 3968 1006
rect 4020 997 4032 1006
rect 4084 997 4096 1006
rect 4148 997 4160 1006
rect 3831 963 3840 997
rect 3903 963 3904 997
rect 4084 963 4085 997
rect 4148 963 4157 997
rect 3828 954 3840 963
rect 3892 954 3904 963
rect 3956 954 3968 963
rect 4020 954 4032 963
rect 4084 954 4096 963
rect 4148 954 4160 963
rect 4212 954 4264 1006
rect 2774 900 2816 901
rect 2758 892 2816 900
rect 2758 840 2769 892
rect 2821 840 2827 892
rect 3118 844 3157 944
rect 3724 910 4264 954
rect 3741 854 3787 910
rect 3736 853 3787 854
rect 2758 797 2816 840
rect 2524 725 2570 763
rect 2524 691 2530 725
rect 2564 691 2570 725
rect 2524 684 2570 691
rect 2613 745 2715 773
rect 2613 711 2647 745
rect 2681 711 2715 745
rect 2524 644 2574 684
rect 2613 683 2715 711
rect 2758 763 2776 797
rect 2810 763 2816 797
rect 2758 725 2816 763
rect 2758 691 2776 725
rect 2810 691 2816 725
rect 1008 584 1052 638
rect 1245 603 1328 622
rect 852 540 1052 584
rect 1148 601 1328 603
rect 1148 549 1155 601
rect 1207 591 1328 601
rect 1207 557 1269 591
rect 1303 557 1328 591
rect 1207 549 1328 557
rect 1148 548 1328 549
rect 852 418 896 540
rect 1245 527 1328 548
rect 1568 610 1602 644
rect 1568 600 1820 610
rect 1568 548 1758 600
rect 1810 548 1820 600
rect 1568 538 1820 548
rect 1568 506 1608 538
rect 1853 506 1892 644
rect 2185 506 2224 644
rect 2255 607 2325 613
rect 2255 598 2331 607
rect 2255 546 2270 598
rect 2322 546 2331 598
rect 2255 537 2331 546
rect 2255 531 2325 537
rect 2368 506 2407 644
rect 2530 610 2574 644
rect 2758 644 2816 691
rect 2928 797 2974 844
rect 2928 763 2934 797
rect 2968 784 2974 797
rect 3114 797 3160 844
rect 3114 784 3120 797
rect 2968 763 3120 784
rect 3154 763 3160 797
rect 3272 797 3318 844
rect 3272 787 3278 797
rect 3312 787 3318 797
rect 3736 807 3782 853
rect 2928 725 3160 763
rect 3262 735 3268 787
rect 3320 735 3326 787
rect 3736 773 3742 807
rect 3776 773 3782 807
rect 3736 735 3782 773
rect 2928 691 2934 725
rect 2968 691 3120 725
rect 3154 691 3160 725
rect 2928 674 3160 691
rect 2928 644 2974 674
rect 3114 644 3160 674
rect 3272 725 3318 735
rect 3272 691 3278 725
rect 3312 691 3318 725
rect 3272 644 3318 691
rect 3736 701 3742 735
rect 3776 701 3782 735
rect 3736 654 3782 701
rect 3894 807 3940 854
rect 3894 773 3900 807
rect 3934 773 3940 807
rect 3894 735 3940 773
rect 3894 701 3900 735
rect 3934 701 3940 735
rect 3894 654 3940 701
rect 4044 807 4090 910
rect 4558 854 4597 1060
rect 4738 1054 4744 1060
rect 4796 1054 4802 1106
rect 4868 854 4907 1141
rect 4044 773 4050 807
rect 4084 773 4090 807
rect 4044 735 4090 773
rect 4044 701 4050 735
rect 4084 701 4090 735
rect 4044 654 4090 701
rect 4202 807 4248 854
rect 4202 773 4208 807
rect 4242 773 4248 807
rect 4396 807 4442 854
rect 4396 781 4402 807
rect 4202 735 4248 773
rect 4202 701 4208 735
rect 4242 701 4248 735
rect 4285 779 4402 781
rect 4285 727 4292 779
rect 4344 773 4402 779
rect 4436 773 4442 807
rect 4344 735 4442 773
rect 4344 727 4402 735
rect 4285 726 4402 727
rect 4202 654 4248 701
rect 4396 701 4402 726
rect 4436 701 4442 735
rect 4396 654 4442 701
rect 4554 807 4600 854
rect 4554 773 4560 807
rect 4594 774 4600 807
rect 4704 807 4750 854
rect 4704 774 4710 807
rect 4594 773 4710 774
rect 4744 773 4750 807
rect 4554 735 4750 773
rect 4554 701 4560 735
rect 4594 708 4710 735
rect 4594 701 4600 708
rect 4554 654 4600 701
rect 4704 701 4710 708
rect 4744 701 4750 735
rect 4704 654 4750 701
rect 4862 807 4908 854
rect 4862 773 4868 807
rect 4902 773 4908 807
rect 5027 778 5057 787
rect 4862 735 4908 773
rect 4862 701 4868 735
rect 4902 701 4908 735
rect 5010 726 5016 778
rect 5068 726 5074 778
rect 4862 654 4908 701
rect 5026 685 5057 726
rect 2758 610 2802 644
rect 2530 566 2656 610
rect 1242 486 1248 490
rect 1138 442 1248 486
rect 1138 418 1182 442
rect 1242 438 1248 442
rect 1300 438 1306 490
rect 1404 473 1450 506
rect 1404 439 1410 473
rect 1444 439 1450 473
rect 1404 435 1450 439
rect 378 390 434 396
rect 550 390 622 412
rect 434 384 622 390
rect 434 344 565 384
rect 606 344 622 384
rect 434 334 622 344
rect 378 328 434 334
rect 550 314 622 334
rect 696 384 768 412
rect 696 344 712 384
rect 753 344 768 384
rect 696 314 768 344
rect 840 389 912 418
rect 840 349 856 389
rect 897 349 912 389
rect 840 320 912 349
rect 994 390 1182 418
rect 994 350 1010 390
rect 1051 374 1182 390
rect 1399 406 1450 435
rect 1562 473 1608 506
rect 1562 439 1568 473
rect 1602 439 1608 473
rect 1692 473 1738 506
rect 1692 444 1698 473
rect 1562 406 1608 439
rect 1690 439 1698 444
rect 1732 444 1738 473
rect 1850 473 1896 506
rect 2024 490 2070 506
rect 1732 439 1740 444
rect 1051 350 1066 374
rect 1399 360 1449 406
rect 1690 360 1740 439
rect 1850 439 1856 473
rect 1890 439 1896 473
rect 1850 406 1896 439
rect 2014 438 2020 490
rect 2072 438 2078 490
rect 2182 473 2228 506
rect 2182 439 2188 473
rect 2222 439 2228 473
rect 2024 406 2070 438
rect 2182 406 2228 439
rect 2366 473 2412 506
rect 2524 488 2570 506
rect 2366 439 2372 473
rect 2406 439 2412 473
rect 2366 406 2412 439
rect 2516 436 2522 488
rect 2574 436 2580 488
rect 2524 406 2570 436
rect 2024 374 2068 406
rect 2612 374 2656 566
rect 994 320 1066 350
rect 1324 305 1960 360
rect 2024 330 2656 374
rect 2694 566 2802 610
rect 2832 596 2904 606
rect 2694 368 2738 566
rect 2832 544 2842 596
rect 2894 544 2904 596
rect 2832 534 2904 544
rect 2933 506 2972 644
rect 3118 506 3157 644
rect 3272 600 3316 644
rect 3268 594 3320 600
rect 3555 569 3561 621
rect 3613 614 3619 621
rect 3662 614 3713 626
rect 3613 611 3713 614
rect 3613 577 3670 611
rect 3704 577 3713 611
rect 3613 575 3713 577
rect 3613 569 3619 575
rect 3662 563 3713 575
rect 3897 605 3936 654
rect 3976 612 4027 617
rect 3970 605 3976 612
rect 3897 566 3976 605
rect 3268 536 3320 542
rect 3897 516 3936 566
rect 3970 560 3976 566
rect 4028 560 4034 612
rect 4206 598 4245 654
rect 4300 598 4347 609
rect 4206 596 4347 598
rect 4206 563 4306 596
rect 3976 554 4027 560
rect 4206 516 4245 563
rect 4300 562 4306 563
rect 4340 562 4347 596
rect 4300 550 4347 562
rect 2766 500 2818 506
rect 2766 442 2776 448
rect 2770 439 2776 442
rect 2810 442 2818 448
rect 2928 473 2974 506
rect 2810 439 2816 442
rect 2770 406 2816 439
rect 2928 439 2934 473
rect 2968 439 2974 473
rect 2928 406 2974 439
rect 3114 473 3160 506
rect 3114 439 3120 473
rect 3154 439 3160 473
rect 3114 406 3160 439
rect 3272 473 3318 506
rect 3272 439 3278 473
rect 3312 439 3318 473
rect 3272 406 3318 439
rect 3274 368 3318 406
rect 2694 324 3318 368
rect 3736 483 3782 516
rect 3736 449 3742 483
rect 3776 449 3782 483
rect 3736 416 3782 449
rect 3894 483 3940 516
rect 3894 449 3900 483
rect 3934 449 3940 483
rect 4044 483 4090 516
rect 4044 454 4050 483
rect 3894 416 3940 449
rect 4042 449 4050 454
rect 4084 449 4090 483
rect 4042 416 4090 449
rect 4202 483 4248 516
rect 4202 449 4208 483
rect 4242 449 4248 483
rect 4202 416 4248 449
rect 3736 360 3780 416
rect 4042 360 4089 416
rect 1324 253 1360 305
rect 1412 253 1424 305
rect 1476 296 1488 305
rect 1540 296 1552 305
rect 1604 296 1616 305
rect 1668 296 1680 305
rect 1732 296 1744 305
rect 1796 296 1808 305
rect 1479 262 1488 296
rect 1551 262 1552 296
rect 1732 262 1733 296
rect 1796 262 1805 296
rect 1476 253 1488 262
rect 1540 253 1552 262
rect 1604 253 1616 262
rect 1668 253 1680 262
rect 1732 253 1744 262
rect 1796 253 1808 262
rect 1860 253 1872 305
rect 1924 253 1960 305
rect 3704 316 4244 360
rect 3704 307 3756 316
rect 3808 307 3820 316
rect 1324 220 1960 253
rect 2346 275 2426 300
rect 2346 271 3517 275
rect 2346 237 2369 271
rect 2403 237 3517 271
rect 2346 233 3517 237
rect 2346 208 2426 233
rect 2636 175 2702 187
rect 272 121 278 175
rect 332 121 2642 175
rect 2696 121 2702 175
rect 2636 109 2702 121
rect 3475 80 3517 233
rect 3704 273 3741 307
rect 3808 273 3813 307
rect 3704 264 3756 273
rect 3808 264 3820 273
rect 3872 264 3884 316
rect 3936 264 3948 316
rect 4000 264 4012 316
rect 4064 264 4076 316
rect 4128 307 4140 316
rect 4192 307 4244 316
rect 4135 273 4140 307
rect 4207 273 4244 307
rect 4128 264 4140 273
rect 4192 264 4244 273
rect 3704 220 4244 264
rect 3559 115 3565 167
rect 3617 160 3623 167
rect 4306 160 4345 550
rect 4558 518 4597 654
rect 4628 623 4680 629
rect 4625 574 4628 620
rect 4680 574 4683 620
rect 4875 578 4904 654
rect 4628 565 4680 571
rect 4875 550 4980 578
rect 4396 485 4442 518
rect 4396 451 4402 485
rect 4436 451 4442 485
rect 4396 418 4442 451
rect 4554 498 4600 518
rect 4704 498 4750 518
rect 4862 498 4908 518
rect 4554 485 4750 498
rect 4554 451 4560 485
rect 4594 451 4710 485
rect 4744 451 4750 485
rect 4554 432 4750 451
rect 4856 446 4862 498
rect 4914 446 4920 498
rect 4554 418 4600 432
rect 4704 418 4750 432
rect 4862 418 4908 446
rect 4402 268 4430 418
rect 4558 373 4597 418
rect 4552 367 4604 373
rect 4552 309 4604 315
rect 4952 268 4980 550
rect 5026 500 5056 685
rect 5009 448 5015 500
rect 5067 448 5073 500
rect 4402 240 4980 268
rect 3617 121 4345 160
rect 3617 115 3623 121
rect 5021 80 5063 448
rect 3475 38 5063 80
<< via1 >>
rect 1398 4682 1450 4691
rect 1462 4682 1514 4691
rect 1398 4648 1417 4682
rect 1417 4648 1450 4682
rect 1462 4648 1489 4682
rect 1489 4648 1514 4682
rect 1398 4639 1450 4648
rect 1462 4639 1514 4648
rect 1526 4682 1578 4691
rect 1526 4648 1527 4682
rect 1527 4648 1561 4682
rect 1561 4648 1578 4682
rect 1526 4639 1578 4648
rect 1590 4682 1642 4691
rect 1590 4648 1599 4682
rect 1599 4648 1633 4682
rect 1633 4648 1642 4682
rect 1590 4639 1642 4648
rect 1654 4682 1706 4691
rect 1654 4648 1671 4682
rect 1671 4648 1705 4682
rect 1705 4648 1706 4682
rect 1654 4639 1706 4648
rect 1718 4682 1770 4691
rect 1782 4682 1834 4691
rect 1718 4648 1743 4682
rect 1743 4648 1770 4682
rect 1782 4648 1815 4682
rect 1815 4648 1834 4682
rect 1718 4639 1770 4648
rect 1782 4639 1834 4648
rect 560 4596 612 4620
rect 560 4568 566 4596
rect 566 4568 607 4596
rect 607 4568 612 4596
rect 702 4596 754 4616
rect 702 4564 710 4596
rect 710 4564 751 4596
rect 751 4564 754 4596
rect 378 4403 433 4458
rect 852 4414 904 4466
rect 378 4118 433 4173
rect 1004 4322 1056 4374
rect 1935 4333 1987 4385
rect 3776 4681 3828 4690
rect 3840 4681 3892 4690
rect 3904 4681 3956 4690
rect 3968 4681 4020 4690
rect 4032 4681 4084 4690
rect 4096 4681 4148 4690
rect 4160 4681 4212 4690
rect 3776 4647 3797 4681
rect 3797 4647 3828 4681
rect 3840 4647 3869 4681
rect 3869 4647 3892 4681
rect 3904 4647 3941 4681
rect 3941 4647 3956 4681
rect 3968 4647 3975 4681
rect 3975 4647 4013 4681
rect 4013 4647 4020 4681
rect 4032 4647 4047 4681
rect 4047 4647 4084 4681
rect 4096 4647 4119 4681
rect 4119 4647 4148 4681
rect 4160 4647 4191 4681
rect 4191 4647 4212 4681
rect 3776 4638 3828 4647
rect 3840 4638 3892 4647
rect 3904 4638 3956 4647
rect 3968 4638 4020 4647
rect 4032 4638 4084 4647
rect 4096 4638 4148 4647
rect 4160 4638 4212 4647
rect 2769 4524 2821 4576
rect 1155 4233 1207 4285
rect 1758 4275 1810 4284
rect 1758 4241 1773 4275
rect 1773 4241 1807 4275
rect 1807 4241 1810 4275
rect 1758 4232 1810 4241
rect 2270 4273 2322 4282
rect 2270 4239 2273 4273
rect 2273 4239 2307 4273
rect 2307 4239 2322 4273
rect 2270 4230 2322 4239
rect 3268 4447 3278 4471
rect 3278 4447 3312 4471
rect 3312 4447 3320 4471
rect 3268 4419 3320 4447
rect 4744 4738 4796 4790
rect 5029 4820 5081 4872
rect 5734 4680 5786 4690
rect 5798 4680 5850 4690
rect 5862 4680 5914 4690
rect 5926 4680 5978 4690
rect 5990 4680 6042 4690
rect 6054 4680 6106 4690
rect 6118 4680 6170 4690
rect 5734 4646 5756 4680
rect 5756 4646 5786 4680
rect 5798 4646 5828 4680
rect 5828 4646 5850 4680
rect 5862 4646 5900 4680
rect 5900 4646 5914 4680
rect 5926 4646 5934 4680
rect 5934 4646 5972 4680
rect 5972 4646 5978 4680
rect 5990 4646 6006 4680
rect 6006 4646 6042 4680
rect 6054 4646 6078 4680
rect 6078 4646 6106 4680
rect 6118 4646 6150 4680
rect 6150 4646 6170 4680
rect 5734 4638 5786 4646
rect 5798 4638 5850 4646
rect 5862 4638 5914 4646
rect 5926 4638 5978 4646
rect 5990 4638 6042 4646
rect 6054 4638 6106 4646
rect 6118 4638 6170 4646
rect 4292 4411 4344 4463
rect 5016 4410 5068 4462
rect 1248 4122 1300 4174
rect 378 4018 434 4074
rect 2020 4157 2072 4174
rect 2020 4123 2030 4157
rect 2030 4123 2064 4157
rect 2064 4123 2072 4157
rect 2020 4122 2072 4123
rect 2522 4157 2574 4172
rect 2522 4123 2530 4157
rect 2530 4123 2564 4157
rect 2564 4123 2574 4157
rect 2522 4120 2574 4123
rect 2842 4271 2894 4280
rect 2842 4237 2857 4271
rect 2857 4237 2891 4271
rect 2891 4237 2894 4271
rect 2842 4228 2894 4237
rect 3268 4226 3320 4278
rect 3561 4253 3613 4305
rect 3976 4286 4028 4296
rect 3976 4252 3984 4286
rect 3984 4252 4018 4286
rect 4018 4252 4028 4286
rect 3976 4244 4028 4252
rect 2766 4157 2818 4184
rect 2766 4132 2776 4157
rect 2776 4132 2810 4157
rect 2810 4132 2818 4157
rect 1360 3980 1412 3989
rect 1360 3946 1373 3980
rect 1373 3946 1407 3980
rect 1407 3946 1412 3980
rect 1360 3937 1412 3946
rect 1424 3980 1476 3989
rect 1488 3980 1540 3989
rect 1552 3980 1604 3989
rect 1616 3980 1668 3989
rect 1680 3980 1732 3989
rect 1744 3980 1796 3989
rect 1808 3980 1860 3989
rect 1424 3946 1445 3980
rect 1445 3946 1476 3980
rect 1488 3946 1517 3980
rect 1517 3946 1540 3980
rect 1552 3946 1589 3980
rect 1589 3946 1604 3980
rect 1616 3946 1623 3980
rect 1623 3946 1661 3980
rect 1661 3946 1668 3980
rect 1680 3946 1695 3980
rect 1695 3946 1732 3980
rect 1744 3946 1767 3980
rect 1767 3946 1796 3980
rect 1808 3946 1839 3980
rect 1839 3946 1860 3980
rect 1424 3937 1476 3946
rect 1488 3937 1540 3946
rect 1552 3937 1604 3946
rect 1616 3937 1668 3946
rect 1680 3937 1732 3946
rect 1744 3937 1796 3946
rect 1808 3937 1860 3946
rect 1872 3980 1924 3989
rect 1872 3946 1877 3980
rect 1877 3946 1911 3980
rect 1911 3946 1924 3980
rect 1872 3937 1924 3946
rect 3756 3991 3808 4000
rect 3820 3991 3872 4000
rect 278 3805 332 3859
rect 3756 3957 3775 3991
rect 3775 3957 3808 3991
rect 3820 3957 3847 3991
rect 3847 3957 3872 3991
rect 3756 3948 3808 3957
rect 3820 3948 3872 3957
rect 3884 3991 3936 4000
rect 3884 3957 3885 3991
rect 3885 3957 3919 3991
rect 3919 3957 3936 3991
rect 3884 3948 3936 3957
rect 3948 3991 4000 4000
rect 3948 3957 3957 3991
rect 3957 3957 3991 3991
rect 3991 3957 4000 3991
rect 3948 3948 4000 3957
rect 4012 3991 4064 4000
rect 4012 3957 4029 3991
rect 4029 3957 4063 3991
rect 4063 3957 4064 3991
rect 4012 3948 4064 3957
rect 4076 3991 4128 4000
rect 4140 3991 4192 4000
rect 4076 3957 4101 3991
rect 4101 3957 4128 3991
rect 4140 3957 4173 3991
rect 4173 3957 4192 3991
rect 4076 3948 4128 3957
rect 4140 3948 4192 3957
rect 3565 3799 3617 3851
rect 4628 4298 4680 4307
rect 4628 4264 4637 4298
rect 4637 4264 4671 4298
rect 4671 4264 4680 4298
rect 4628 4255 4680 4264
rect 4862 4169 4914 4182
rect 4862 4135 4868 4169
rect 4868 4135 4902 4169
rect 4902 4135 4914 4169
rect 4862 4130 4914 4135
rect 4552 3999 4604 4051
rect 6868 4738 6920 4790
rect 6250 4412 6302 4464
rect 6974 4410 7026 4462
rect 5117 4253 5169 4305
rect 5934 4286 5986 4296
rect 5934 4252 5942 4286
rect 5942 4252 5976 4286
rect 5976 4252 5986 4286
rect 5934 4244 5986 4252
rect 5015 4132 5067 4184
rect 5714 3992 5766 4000
rect 5778 3992 5830 4000
rect 5714 3958 5734 3992
rect 5734 3958 5766 3992
rect 5778 3958 5806 3992
rect 5806 3958 5830 3992
rect 5714 3948 5766 3958
rect 5778 3948 5830 3958
rect 5842 3992 5894 4000
rect 5842 3958 5844 3992
rect 5844 3958 5878 3992
rect 5878 3958 5894 3992
rect 5842 3948 5894 3958
rect 5906 3992 5958 4000
rect 5906 3958 5916 3992
rect 5916 3958 5950 3992
rect 5950 3958 5958 3992
rect 5906 3948 5958 3958
rect 5970 3992 6022 4000
rect 5970 3958 5988 3992
rect 5988 3958 6022 3992
rect 5970 3948 6022 3958
rect 6034 3992 6086 4000
rect 6098 3992 6150 4000
rect 6034 3958 6060 3992
rect 6060 3958 6086 3992
rect 6098 3958 6132 3992
rect 6132 3958 6150 3992
rect 6034 3948 6086 3958
rect 6098 3948 6150 3958
rect 5117 3799 5169 3851
rect 6586 4298 6638 4308
rect 6586 4264 6596 4298
rect 6596 4264 6630 4298
rect 6630 4264 6638 4298
rect 6586 4256 6638 4264
rect 6820 4170 6872 4182
rect 6820 4136 6826 4170
rect 6826 4136 6860 4170
rect 6860 4136 6872 4170
rect 6820 4130 6872 4136
rect 6510 4000 6562 4052
rect 6974 4132 7026 4184
rect 5035 3629 5087 3681
rect 6512 3714 6564 3766
rect 1398 3454 1450 3463
rect 1462 3454 1514 3463
rect 1398 3420 1417 3454
rect 1417 3420 1450 3454
rect 1462 3420 1489 3454
rect 1489 3420 1514 3454
rect 1398 3411 1450 3420
rect 1462 3411 1514 3420
rect 1526 3454 1578 3463
rect 1526 3420 1527 3454
rect 1527 3420 1561 3454
rect 1561 3420 1578 3454
rect 1526 3411 1578 3420
rect 1590 3454 1642 3463
rect 1590 3420 1599 3454
rect 1599 3420 1633 3454
rect 1633 3420 1642 3454
rect 1590 3411 1642 3420
rect 1654 3454 1706 3463
rect 1654 3420 1671 3454
rect 1671 3420 1705 3454
rect 1705 3420 1706 3454
rect 1654 3411 1706 3420
rect 1718 3454 1770 3463
rect 1782 3454 1834 3463
rect 1718 3420 1743 3454
rect 1743 3420 1770 3454
rect 1782 3420 1815 3454
rect 1815 3420 1834 3454
rect 1718 3411 1770 3420
rect 1782 3411 1834 3420
rect 560 3368 612 3392
rect 560 3340 566 3368
rect 566 3340 607 3368
rect 607 3340 612 3368
rect 702 3368 754 3388
rect 702 3336 710 3368
rect 710 3336 751 3368
rect 751 3336 754 3368
rect 378 3175 433 3230
rect 852 3186 904 3238
rect 378 2890 433 2945
rect 1004 3094 1056 3146
rect 1935 3105 1987 3157
rect 3776 3453 3828 3462
rect 3840 3453 3892 3462
rect 3904 3453 3956 3462
rect 3968 3453 4020 3462
rect 4032 3453 4084 3462
rect 4096 3453 4148 3462
rect 4160 3453 4212 3462
rect 3776 3419 3797 3453
rect 3797 3419 3828 3453
rect 3840 3419 3869 3453
rect 3869 3419 3892 3453
rect 3904 3419 3941 3453
rect 3941 3419 3956 3453
rect 3968 3419 3975 3453
rect 3975 3419 4013 3453
rect 4013 3419 4020 3453
rect 4032 3419 4047 3453
rect 4047 3419 4084 3453
rect 4096 3419 4119 3453
rect 4119 3419 4148 3453
rect 4160 3419 4191 3453
rect 4191 3419 4212 3453
rect 3776 3410 3828 3419
rect 3840 3410 3892 3419
rect 3904 3410 3956 3419
rect 3968 3410 4020 3419
rect 4032 3410 4084 3419
rect 4096 3410 4148 3419
rect 4160 3410 4212 3419
rect 2769 3296 2821 3348
rect 1155 3005 1207 3057
rect 1758 3047 1810 3056
rect 1758 3013 1773 3047
rect 1773 3013 1807 3047
rect 1807 3013 1810 3047
rect 1758 3004 1810 3013
rect 2270 3045 2322 3054
rect 2270 3011 2273 3045
rect 2273 3011 2307 3045
rect 2307 3011 2322 3045
rect 2270 3002 2322 3011
rect 3268 3219 3278 3243
rect 3278 3219 3312 3243
rect 3312 3219 3320 3243
rect 3268 3191 3320 3219
rect 4744 3510 4796 3562
rect 5734 3452 5786 3462
rect 5798 3452 5850 3462
rect 5862 3452 5914 3462
rect 5926 3452 5978 3462
rect 5990 3452 6042 3462
rect 6054 3452 6106 3462
rect 6118 3452 6170 3462
rect 5734 3418 5756 3452
rect 5756 3418 5786 3452
rect 5798 3418 5828 3452
rect 5828 3418 5850 3452
rect 5862 3418 5900 3452
rect 5900 3418 5914 3452
rect 5926 3418 5934 3452
rect 5934 3418 5972 3452
rect 5972 3418 5978 3452
rect 5990 3418 6006 3452
rect 6006 3418 6042 3452
rect 6054 3418 6078 3452
rect 6078 3418 6106 3452
rect 6118 3418 6150 3452
rect 6150 3418 6170 3452
rect 5734 3410 5786 3418
rect 5798 3410 5850 3418
rect 5862 3410 5914 3418
rect 5926 3410 5978 3418
rect 5990 3410 6042 3418
rect 6054 3410 6106 3418
rect 6118 3410 6170 3418
rect 4292 3183 4344 3235
rect 5016 3182 5068 3234
rect 1248 2894 1300 2946
rect 378 2790 434 2846
rect 2020 2929 2072 2946
rect 2020 2895 2030 2929
rect 2030 2895 2064 2929
rect 2064 2895 2072 2929
rect 2020 2894 2072 2895
rect 2522 2929 2574 2944
rect 2522 2895 2530 2929
rect 2530 2895 2564 2929
rect 2564 2895 2574 2929
rect 2522 2892 2574 2895
rect 2842 3043 2894 3052
rect 2842 3009 2857 3043
rect 2857 3009 2891 3043
rect 2891 3009 2894 3043
rect 2842 3000 2894 3009
rect 3268 2998 3320 3050
rect 3561 3025 3613 3077
rect 3976 3058 4028 3068
rect 3976 3024 3984 3058
rect 3984 3024 4018 3058
rect 4018 3024 4028 3058
rect 3976 3016 4028 3024
rect 2766 2929 2818 2956
rect 2766 2904 2776 2929
rect 2776 2904 2810 2929
rect 2810 2904 2818 2929
rect 1360 2752 1412 2761
rect 1360 2718 1373 2752
rect 1373 2718 1407 2752
rect 1407 2718 1412 2752
rect 1360 2709 1412 2718
rect 1424 2752 1476 2761
rect 1488 2752 1540 2761
rect 1552 2752 1604 2761
rect 1616 2752 1668 2761
rect 1680 2752 1732 2761
rect 1744 2752 1796 2761
rect 1808 2752 1860 2761
rect 1424 2718 1445 2752
rect 1445 2718 1476 2752
rect 1488 2718 1517 2752
rect 1517 2718 1540 2752
rect 1552 2718 1589 2752
rect 1589 2718 1604 2752
rect 1616 2718 1623 2752
rect 1623 2718 1661 2752
rect 1661 2718 1668 2752
rect 1680 2718 1695 2752
rect 1695 2718 1732 2752
rect 1744 2718 1767 2752
rect 1767 2718 1796 2752
rect 1808 2718 1839 2752
rect 1839 2718 1860 2752
rect 1424 2709 1476 2718
rect 1488 2709 1540 2718
rect 1552 2709 1604 2718
rect 1616 2709 1668 2718
rect 1680 2709 1732 2718
rect 1744 2709 1796 2718
rect 1808 2709 1860 2718
rect 1872 2752 1924 2761
rect 1872 2718 1877 2752
rect 1877 2718 1911 2752
rect 1911 2718 1924 2752
rect 1872 2709 1924 2718
rect 3756 2763 3808 2772
rect 3820 2763 3872 2772
rect 278 2577 332 2631
rect 3756 2729 3775 2763
rect 3775 2729 3808 2763
rect 3820 2729 3847 2763
rect 3847 2729 3872 2763
rect 3756 2720 3808 2729
rect 3820 2720 3872 2729
rect 3884 2763 3936 2772
rect 3884 2729 3885 2763
rect 3885 2729 3919 2763
rect 3919 2729 3936 2763
rect 3884 2720 3936 2729
rect 3948 2763 4000 2772
rect 3948 2729 3957 2763
rect 3957 2729 3991 2763
rect 3991 2729 4000 2763
rect 3948 2720 4000 2729
rect 4012 2763 4064 2772
rect 4012 2729 4029 2763
rect 4029 2729 4063 2763
rect 4063 2729 4064 2763
rect 4012 2720 4064 2729
rect 4076 2763 4128 2772
rect 4140 2763 4192 2772
rect 4076 2729 4101 2763
rect 4101 2729 4128 2763
rect 4140 2729 4173 2763
rect 4173 2729 4192 2763
rect 4076 2720 4128 2729
rect 4140 2720 4192 2729
rect 3565 2571 3617 2623
rect 4628 3070 4680 3079
rect 4628 3036 4637 3070
rect 4637 3036 4671 3070
rect 4671 3036 4680 3070
rect 4628 3027 4680 3036
rect 4862 2941 4914 2954
rect 4862 2907 4868 2941
rect 4868 2907 4902 2941
rect 4902 2907 4914 2941
rect 4862 2902 4914 2907
rect 4552 2771 4604 2823
rect 6843 3510 6895 3562
rect 6250 3184 6302 3236
rect 6974 3182 7026 3234
rect 5197 3025 5249 3077
rect 5934 3058 5986 3068
rect 5934 3024 5942 3058
rect 5942 3024 5976 3058
rect 5976 3024 5986 3058
rect 5934 3016 5986 3024
rect 5015 2904 5067 2956
rect 5714 2764 5766 2772
rect 5778 2764 5830 2772
rect 5714 2730 5734 2764
rect 5734 2730 5766 2764
rect 5778 2730 5806 2764
rect 5806 2730 5830 2764
rect 5714 2720 5766 2730
rect 5778 2720 5830 2730
rect 5842 2764 5894 2772
rect 5842 2730 5844 2764
rect 5844 2730 5878 2764
rect 5878 2730 5894 2764
rect 5842 2720 5894 2730
rect 5906 2764 5958 2772
rect 5906 2730 5916 2764
rect 5916 2730 5950 2764
rect 5950 2730 5958 2764
rect 5906 2720 5958 2730
rect 5970 2764 6022 2772
rect 5970 2730 5988 2764
rect 5988 2730 6022 2764
rect 5970 2720 6022 2730
rect 6034 2764 6086 2772
rect 6098 2764 6150 2772
rect 6034 2730 6060 2764
rect 6060 2730 6086 2764
rect 6098 2730 6132 2764
rect 6132 2730 6150 2764
rect 6034 2720 6086 2730
rect 6098 2720 6150 2730
rect 5197 2571 5249 2623
rect 6586 3070 6638 3080
rect 6586 3036 6596 3070
rect 6596 3036 6630 3070
rect 6630 3036 6638 3070
rect 6586 3028 6638 3036
rect 6820 2942 6872 2954
rect 6820 2908 6826 2942
rect 6826 2908 6860 2942
rect 6860 2908 6872 2942
rect 6820 2902 6872 2908
rect 6510 2772 6562 2824
rect 6974 2904 7026 2956
rect 7107 2484 7159 2536
rect 1398 2226 1450 2235
rect 1462 2226 1514 2235
rect 1398 2192 1417 2226
rect 1417 2192 1450 2226
rect 1462 2192 1489 2226
rect 1489 2192 1514 2226
rect 1398 2183 1450 2192
rect 1462 2183 1514 2192
rect 1526 2226 1578 2235
rect 1526 2192 1527 2226
rect 1527 2192 1561 2226
rect 1561 2192 1578 2226
rect 1526 2183 1578 2192
rect 1590 2226 1642 2235
rect 1590 2192 1599 2226
rect 1599 2192 1633 2226
rect 1633 2192 1642 2226
rect 1590 2183 1642 2192
rect 1654 2226 1706 2235
rect 1654 2192 1671 2226
rect 1671 2192 1705 2226
rect 1705 2192 1706 2226
rect 1654 2183 1706 2192
rect 1718 2226 1770 2235
rect 1782 2226 1834 2235
rect 1718 2192 1743 2226
rect 1743 2192 1770 2226
rect 1782 2192 1815 2226
rect 1815 2192 1834 2226
rect 1718 2183 1770 2192
rect 1782 2183 1834 2192
rect 560 2140 612 2164
rect 560 2112 566 2140
rect 566 2112 607 2140
rect 607 2112 612 2140
rect 702 2140 754 2160
rect 702 2108 710 2140
rect 710 2108 751 2140
rect 751 2108 754 2140
rect 378 1947 433 2002
rect 852 1958 904 2010
rect 378 1662 433 1717
rect 1004 1866 1056 1918
rect 1935 1877 1987 1929
rect 3776 2225 3828 2234
rect 3840 2225 3892 2234
rect 3904 2225 3956 2234
rect 3968 2225 4020 2234
rect 4032 2225 4084 2234
rect 4096 2225 4148 2234
rect 4160 2225 4212 2234
rect 3776 2191 3797 2225
rect 3797 2191 3828 2225
rect 3840 2191 3869 2225
rect 3869 2191 3892 2225
rect 3904 2191 3941 2225
rect 3941 2191 3956 2225
rect 3968 2191 3975 2225
rect 3975 2191 4013 2225
rect 4013 2191 4020 2225
rect 4032 2191 4047 2225
rect 4047 2191 4084 2225
rect 4096 2191 4119 2225
rect 4119 2191 4148 2225
rect 4160 2191 4191 2225
rect 4191 2191 4212 2225
rect 3776 2182 3828 2191
rect 3840 2182 3892 2191
rect 3904 2182 3956 2191
rect 3968 2182 4020 2191
rect 4032 2182 4084 2191
rect 4096 2182 4148 2191
rect 4160 2182 4212 2191
rect 2769 2068 2821 2120
rect 1155 1777 1207 1829
rect 1758 1819 1810 1828
rect 1758 1785 1773 1819
rect 1773 1785 1807 1819
rect 1807 1785 1810 1819
rect 1758 1776 1810 1785
rect 2270 1817 2322 1826
rect 2270 1783 2273 1817
rect 2273 1783 2307 1817
rect 2307 1783 2322 1817
rect 2270 1774 2322 1783
rect 3268 1991 3278 2015
rect 3278 1991 3312 2015
rect 3312 1991 3320 2015
rect 3268 1963 3320 1991
rect 4744 2282 4796 2334
rect 5029 2364 5081 2416
rect 5734 2224 5786 2234
rect 5798 2224 5850 2234
rect 5862 2224 5914 2234
rect 5926 2224 5978 2234
rect 5990 2224 6042 2234
rect 6054 2224 6106 2234
rect 6118 2224 6170 2234
rect 5734 2190 5756 2224
rect 5756 2190 5786 2224
rect 5798 2190 5828 2224
rect 5828 2190 5850 2224
rect 5862 2190 5900 2224
rect 5900 2190 5914 2224
rect 5926 2190 5934 2224
rect 5934 2190 5972 2224
rect 5972 2190 5978 2224
rect 5990 2190 6006 2224
rect 6006 2190 6042 2224
rect 6054 2190 6078 2224
rect 6078 2190 6106 2224
rect 6118 2190 6150 2224
rect 6150 2190 6170 2224
rect 5734 2182 5786 2190
rect 5798 2182 5850 2190
rect 5862 2182 5914 2190
rect 5926 2182 5978 2190
rect 5990 2182 6042 2190
rect 6054 2182 6106 2190
rect 6118 2182 6170 2190
rect 4292 1955 4344 2007
rect 5016 1954 5068 2006
rect 1248 1666 1300 1718
rect 378 1562 434 1618
rect 2020 1701 2072 1718
rect 2020 1667 2030 1701
rect 2030 1667 2064 1701
rect 2064 1667 2072 1701
rect 2020 1666 2072 1667
rect 2522 1701 2574 1716
rect 2522 1667 2530 1701
rect 2530 1667 2564 1701
rect 2564 1667 2574 1701
rect 2522 1664 2574 1667
rect 2842 1815 2894 1824
rect 2842 1781 2857 1815
rect 2857 1781 2891 1815
rect 2891 1781 2894 1815
rect 2842 1772 2894 1781
rect 3268 1770 3320 1822
rect 3561 1797 3613 1849
rect 3976 1830 4028 1840
rect 3976 1796 3984 1830
rect 3984 1796 4018 1830
rect 4018 1796 4028 1830
rect 3976 1788 4028 1796
rect 2766 1701 2818 1728
rect 2766 1676 2776 1701
rect 2776 1676 2810 1701
rect 2810 1676 2818 1701
rect 1360 1524 1412 1533
rect 1360 1490 1373 1524
rect 1373 1490 1407 1524
rect 1407 1490 1412 1524
rect 1360 1481 1412 1490
rect 1424 1524 1476 1533
rect 1488 1524 1540 1533
rect 1552 1524 1604 1533
rect 1616 1524 1668 1533
rect 1680 1524 1732 1533
rect 1744 1524 1796 1533
rect 1808 1524 1860 1533
rect 1424 1490 1445 1524
rect 1445 1490 1476 1524
rect 1488 1490 1517 1524
rect 1517 1490 1540 1524
rect 1552 1490 1589 1524
rect 1589 1490 1604 1524
rect 1616 1490 1623 1524
rect 1623 1490 1661 1524
rect 1661 1490 1668 1524
rect 1680 1490 1695 1524
rect 1695 1490 1732 1524
rect 1744 1490 1767 1524
rect 1767 1490 1796 1524
rect 1808 1490 1839 1524
rect 1839 1490 1860 1524
rect 1424 1481 1476 1490
rect 1488 1481 1540 1490
rect 1552 1481 1604 1490
rect 1616 1481 1668 1490
rect 1680 1481 1732 1490
rect 1744 1481 1796 1490
rect 1808 1481 1860 1490
rect 1872 1524 1924 1533
rect 1872 1490 1877 1524
rect 1877 1490 1911 1524
rect 1911 1490 1924 1524
rect 1872 1481 1924 1490
rect 3756 1535 3808 1544
rect 3820 1535 3872 1544
rect 278 1349 332 1403
rect 3756 1501 3775 1535
rect 3775 1501 3808 1535
rect 3820 1501 3847 1535
rect 3847 1501 3872 1535
rect 3756 1492 3808 1501
rect 3820 1492 3872 1501
rect 3884 1535 3936 1544
rect 3884 1501 3885 1535
rect 3885 1501 3919 1535
rect 3919 1501 3936 1535
rect 3884 1492 3936 1501
rect 3948 1535 4000 1544
rect 3948 1501 3957 1535
rect 3957 1501 3991 1535
rect 3991 1501 4000 1535
rect 3948 1492 4000 1501
rect 4012 1535 4064 1544
rect 4012 1501 4029 1535
rect 4029 1501 4063 1535
rect 4063 1501 4064 1535
rect 4012 1492 4064 1501
rect 4076 1535 4128 1544
rect 4140 1535 4192 1544
rect 4076 1501 4101 1535
rect 4101 1501 4128 1535
rect 4140 1501 4173 1535
rect 4173 1501 4192 1535
rect 4076 1492 4128 1501
rect 4140 1492 4192 1501
rect 3565 1343 3617 1395
rect 4628 1842 4680 1851
rect 4628 1808 4637 1842
rect 4637 1808 4671 1842
rect 4671 1808 4680 1842
rect 4628 1799 4680 1808
rect 4862 1713 4914 1726
rect 4862 1679 4868 1713
rect 4868 1679 4902 1713
rect 4902 1679 4914 1713
rect 4862 1674 4914 1679
rect 4552 1543 4604 1595
rect 6868 2282 6920 2334
rect 6250 1956 6302 2008
rect 6974 1954 7026 2006
rect 5117 1797 5169 1849
rect 5934 1830 5986 1840
rect 5934 1796 5942 1830
rect 5942 1796 5976 1830
rect 5976 1796 5986 1830
rect 5934 1788 5986 1796
rect 5015 1676 5067 1728
rect 5714 1536 5766 1544
rect 5778 1536 5830 1544
rect 5714 1502 5734 1536
rect 5734 1502 5766 1536
rect 5778 1502 5806 1536
rect 5806 1502 5830 1536
rect 5714 1492 5766 1502
rect 5778 1492 5830 1502
rect 5842 1536 5894 1544
rect 5842 1502 5844 1536
rect 5844 1502 5878 1536
rect 5878 1502 5894 1536
rect 5842 1492 5894 1502
rect 5906 1536 5958 1544
rect 5906 1502 5916 1536
rect 5916 1502 5950 1536
rect 5950 1502 5958 1536
rect 5906 1492 5958 1502
rect 5970 1536 6022 1544
rect 5970 1502 5988 1536
rect 5988 1502 6022 1536
rect 5970 1492 6022 1502
rect 6034 1536 6086 1544
rect 6098 1536 6150 1544
rect 6034 1502 6060 1536
rect 6060 1502 6086 1536
rect 6098 1502 6132 1536
rect 6132 1502 6150 1536
rect 6034 1492 6086 1502
rect 6098 1492 6150 1502
rect 5117 1343 5169 1395
rect 6586 1842 6638 1852
rect 6586 1808 6596 1842
rect 6596 1808 6630 1842
rect 6630 1808 6638 1842
rect 6586 1800 6638 1808
rect 6820 1714 6872 1726
rect 6820 1680 6826 1714
rect 6826 1680 6860 1714
rect 6860 1680 6872 1714
rect 6820 1674 6872 1680
rect 6510 1544 6562 1596
rect 6974 1676 7026 1728
rect 5035 1173 5087 1225
rect 1398 998 1450 1007
rect 1462 998 1514 1007
rect 1398 964 1417 998
rect 1417 964 1450 998
rect 1462 964 1489 998
rect 1489 964 1514 998
rect 1398 955 1450 964
rect 1462 955 1514 964
rect 1526 998 1578 1007
rect 1526 964 1527 998
rect 1527 964 1561 998
rect 1561 964 1578 998
rect 1526 955 1578 964
rect 1590 998 1642 1007
rect 1590 964 1599 998
rect 1599 964 1633 998
rect 1633 964 1642 998
rect 1590 955 1642 964
rect 1654 998 1706 1007
rect 1654 964 1671 998
rect 1671 964 1705 998
rect 1705 964 1706 998
rect 1654 955 1706 964
rect 1718 998 1770 1007
rect 1782 998 1834 1007
rect 1718 964 1743 998
rect 1743 964 1770 998
rect 1782 964 1815 998
rect 1815 964 1834 998
rect 1718 955 1770 964
rect 1782 955 1834 964
rect 560 912 612 936
rect 560 884 566 912
rect 566 884 607 912
rect 607 884 612 912
rect 702 912 754 932
rect 702 880 710 912
rect 710 880 751 912
rect 751 880 754 912
rect 378 719 433 774
rect 852 730 904 782
rect 378 434 433 489
rect 1004 638 1056 690
rect 1935 649 1987 701
rect 3776 997 3828 1006
rect 3840 997 3892 1006
rect 3904 997 3956 1006
rect 3968 997 4020 1006
rect 4032 997 4084 1006
rect 4096 997 4148 1006
rect 4160 997 4212 1006
rect 3776 963 3797 997
rect 3797 963 3828 997
rect 3840 963 3869 997
rect 3869 963 3892 997
rect 3904 963 3941 997
rect 3941 963 3956 997
rect 3968 963 3975 997
rect 3975 963 4013 997
rect 4013 963 4020 997
rect 4032 963 4047 997
rect 4047 963 4084 997
rect 4096 963 4119 997
rect 4119 963 4148 997
rect 4160 963 4191 997
rect 4191 963 4212 997
rect 3776 954 3828 963
rect 3840 954 3892 963
rect 3904 954 3956 963
rect 3968 954 4020 963
rect 4032 954 4084 963
rect 4096 954 4148 963
rect 4160 954 4212 963
rect 2769 840 2821 892
rect 1155 549 1207 601
rect 1758 591 1810 600
rect 1758 557 1773 591
rect 1773 557 1807 591
rect 1807 557 1810 591
rect 1758 548 1810 557
rect 2270 589 2322 598
rect 2270 555 2273 589
rect 2273 555 2307 589
rect 2307 555 2322 589
rect 2270 546 2322 555
rect 3268 763 3278 787
rect 3278 763 3312 787
rect 3312 763 3320 787
rect 3268 735 3320 763
rect 4744 1054 4796 1106
rect 4292 727 4344 779
rect 5016 726 5068 778
rect 1248 438 1300 490
rect 378 334 434 390
rect 2020 473 2072 490
rect 2020 439 2030 473
rect 2030 439 2064 473
rect 2064 439 2072 473
rect 2020 438 2072 439
rect 2522 473 2574 488
rect 2522 439 2530 473
rect 2530 439 2564 473
rect 2564 439 2574 473
rect 2522 436 2574 439
rect 2842 587 2894 596
rect 2842 553 2857 587
rect 2857 553 2891 587
rect 2891 553 2894 587
rect 2842 544 2894 553
rect 3268 542 3320 594
rect 3561 569 3613 621
rect 3976 602 4028 612
rect 3976 568 3984 602
rect 3984 568 4018 602
rect 4018 568 4028 602
rect 3976 560 4028 568
rect 2766 473 2818 500
rect 2766 448 2776 473
rect 2776 448 2810 473
rect 2810 448 2818 473
rect 1360 296 1412 305
rect 1360 262 1373 296
rect 1373 262 1407 296
rect 1407 262 1412 296
rect 1360 253 1412 262
rect 1424 296 1476 305
rect 1488 296 1540 305
rect 1552 296 1604 305
rect 1616 296 1668 305
rect 1680 296 1732 305
rect 1744 296 1796 305
rect 1808 296 1860 305
rect 1424 262 1445 296
rect 1445 262 1476 296
rect 1488 262 1517 296
rect 1517 262 1540 296
rect 1552 262 1589 296
rect 1589 262 1604 296
rect 1616 262 1623 296
rect 1623 262 1661 296
rect 1661 262 1668 296
rect 1680 262 1695 296
rect 1695 262 1732 296
rect 1744 262 1767 296
rect 1767 262 1796 296
rect 1808 262 1839 296
rect 1839 262 1860 296
rect 1424 253 1476 262
rect 1488 253 1540 262
rect 1552 253 1604 262
rect 1616 253 1668 262
rect 1680 253 1732 262
rect 1744 253 1796 262
rect 1808 253 1860 262
rect 1872 296 1924 305
rect 1872 262 1877 296
rect 1877 262 1911 296
rect 1911 262 1924 296
rect 1872 253 1924 262
rect 3756 307 3808 316
rect 3820 307 3872 316
rect 278 121 332 175
rect 3756 273 3775 307
rect 3775 273 3808 307
rect 3820 273 3847 307
rect 3847 273 3872 307
rect 3756 264 3808 273
rect 3820 264 3872 273
rect 3884 307 3936 316
rect 3884 273 3885 307
rect 3885 273 3919 307
rect 3919 273 3936 307
rect 3884 264 3936 273
rect 3948 307 4000 316
rect 3948 273 3957 307
rect 3957 273 3991 307
rect 3991 273 4000 307
rect 3948 264 4000 273
rect 4012 307 4064 316
rect 4012 273 4029 307
rect 4029 273 4063 307
rect 4063 273 4064 307
rect 4012 264 4064 273
rect 4076 307 4128 316
rect 4140 307 4192 316
rect 4076 273 4101 307
rect 4101 273 4128 307
rect 4140 273 4173 307
rect 4173 273 4192 307
rect 4076 264 4128 273
rect 4140 264 4192 273
rect 3565 115 3617 167
rect 4628 614 4680 623
rect 4628 580 4637 614
rect 4637 580 4671 614
rect 4671 580 4680 614
rect 4628 571 4680 580
rect 4862 485 4914 498
rect 4862 451 4868 485
rect 4868 451 4902 485
rect 4902 451 4914 485
rect 4862 446 4914 451
rect 4552 315 4604 367
rect 5015 448 5067 500
<< metal2 >>
rect 42 4690 110 4699
rect 42 3484 110 4622
rect 274 4287 329 4912
rect 378 4458 433 4912
rect 1348 4693 1880 4734
rect 1348 4637 1388 4693
rect 1444 4691 1468 4693
rect 1524 4691 1548 4693
rect 1604 4691 1628 4693
rect 1684 4691 1708 4693
rect 1764 4691 1788 4693
rect 1450 4639 1462 4691
rect 1524 4639 1526 4691
rect 1706 4639 1708 4691
rect 1770 4639 1782 4691
rect 1444 4637 1468 4639
rect 1524 4637 1548 4639
rect 1604 4637 1628 4639
rect 1684 4637 1708 4639
rect 1764 4637 1788 4639
rect 1844 4637 1880 4693
rect 560 4620 612 4626
rect 700 4618 756 4624
rect 612 4616 976 4618
rect 612 4568 702 4616
rect 560 4564 702 4568
rect 754 4564 976 4616
rect 1348 4594 1880 4637
rect 2759 4576 2827 4584
rect 560 4562 1268 4564
rect 700 4556 756 4562
rect 920 4556 1268 4562
rect 2759 4556 2769 4576
rect 920 4524 2769 4556
rect 2821 4524 2827 4576
rect 920 4512 2827 4524
rect 920 4508 1268 4512
rect 852 4466 904 4472
rect 372 4403 378 4458
rect 433 4403 439 4458
rect 1396 4467 2851 4476
rect 3268 4471 3320 4477
rect 1396 4462 3268 4467
rect 904 4432 3268 4462
rect 904 4418 1440 4432
rect 2851 4423 3268 4432
rect 852 4408 904 4414
rect 3268 4413 3320 4419
rect 1930 4386 1990 4397
rect 1004 4374 1056 4380
rect 1930 4375 1932 4386
rect 1056 4363 1242 4370
rect 1599 4363 1932 4375
rect 1056 4341 1932 4363
rect 1056 4329 1633 4341
rect 1930 4330 1932 4341
rect 1988 4375 1990 4386
rect 1988 4341 1991 4375
rect 1988 4330 1990 4341
rect 1056 4326 1242 4329
rect 1004 4316 1056 4322
rect 1930 4319 1990 4330
rect 3564 4311 3605 4912
rect 5023 4820 5029 4872
rect 5081 4820 5087 4872
rect 5122 4824 5163 4912
rect 5202 4824 5243 4912
rect 5282 4824 5323 4912
rect 5362 4824 5403 4912
rect 5442 4824 5483 4912
rect 5522 4824 5563 4912
rect 4744 4790 4796 4796
rect 5036 4784 5075 4820
rect 4796 4745 5075 4784
rect 3724 4692 4264 4734
rect 4744 4732 4796 4738
rect 3724 4636 3766 4692
rect 3822 4690 3846 4692
rect 3902 4690 3926 4692
rect 3982 4690 4006 4692
rect 4062 4690 4086 4692
rect 4142 4690 4166 4692
rect 3828 4638 3840 4690
rect 3902 4638 3904 4690
rect 4084 4638 4086 4690
rect 4148 4638 4160 4690
rect 3822 4636 3846 4638
rect 3902 4636 3926 4638
rect 3982 4636 4006 4638
rect 4062 4636 4086 4638
rect 4142 4636 4166 4638
rect 4222 4636 4264 4692
rect 3724 4594 4264 4636
rect 4291 4465 4346 4471
rect 5016 4465 5068 4468
rect 4291 4463 5084 4465
rect 4291 4411 4292 4463
rect 4344 4462 5084 4463
rect 4344 4411 5016 4462
rect 4291 4410 5016 4411
rect 5068 4410 5084 4462
rect 4291 4404 4346 4410
rect 5016 4404 5068 4410
rect 5122 4311 5164 4824
rect 3561 4305 3613 4311
rect 1154 4287 1209 4293
rect 274 4285 1209 4287
rect 274 4233 1155 4285
rect 1207 4233 1209 4285
rect 274 4232 1209 4233
rect 1154 4226 1209 4232
rect 1754 4288 1814 4294
rect 2267 4288 2325 4297
rect 1754 4285 2325 4288
rect 2838 4285 2898 4290
rect 1754 4284 2898 4285
rect 1754 4232 1758 4284
rect 1810 4282 2908 4284
rect 1810 4232 2270 4282
rect 1754 4230 2270 4232
rect 2322 4280 2908 4282
rect 2322 4230 2842 4280
rect 1754 4228 2842 4230
rect 2894 4228 2908 4280
rect 1754 4222 1814 4228
rect 2267 4227 2908 4228
rect 2267 4215 2325 4227
rect 2838 4224 2908 4227
rect 3262 4226 3268 4278
rect 3320 4226 3326 4278
rect 3976 4296 4028 4302
rect 3561 4247 3613 4253
rect 3975 4247 3976 4290
rect 2838 4218 2898 4224
rect 2768 4184 2816 4188
rect 378 4173 433 4179
rect 1248 4174 1300 4180
rect 433 4170 619 4173
rect 433 4126 1248 4170
rect 433 4118 619 4126
rect 2020 4174 2072 4180
rect 2522 4176 2574 4178
rect 1300 4126 2020 4170
rect 378 4112 433 4118
rect 1248 4116 1300 4122
rect 2020 4116 2072 4122
rect 2509 4174 2587 4176
rect 2509 4118 2520 4174
rect 2576 4118 2587 4174
rect 2760 4132 2766 4184
rect 2818 4180 2824 4184
rect 3270 4180 3314 4226
rect 3564 4208 3605 4247
rect 4622 4255 4628 4307
rect 4680 4255 4686 4307
rect 5117 4305 5169 4311
rect 3976 4238 4028 4244
rect 2818 4136 3314 4180
rect 3979 4191 4018 4238
rect 4637 4191 4671 4255
rect 5117 4247 5169 4253
rect 5122 4208 5164 4247
rect 5202 4208 5244 4824
rect 5282 4208 5324 4824
rect 5362 4208 5404 4824
rect 5442 4208 5484 4824
rect 5522 4208 5564 4824
rect 6868 4790 6920 4796
rect 6920 4745 7147 4784
rect 5682 4692 6222 4734
rect 6868 4732 6920 4738
rect 5682 4636 5724 4692
rect 5780 4690 5804 4692
rect 5860 4690 5884 4692
rect 5940 4690 5964 4692
rect 6020 4690 6044 4692
rect 6100 4690 6124 4692
rect 5786 4638 5798 4690
rect 5860 4638 5862 4690
rect 6042 4638 6044 4690
rect 6106 4638 6118 4690
rect 5780 4636 5804 4638
rect 5860 4636 5884 4638
rect 5940 4636 5964 4638
rect 6020 4636 6044 4638
rect 6100 4636 6124 4638
rect 6180 4636 6222 4692
rect 5682 4594 6222 4636
rect 6250 4466 6304 4472
rect 6974 4466 7026 4468
rect 6250 4464 7042 4466
rect 6302 4462 7042 4464
rect 6302 4412 6974 4462
rect 6250 4410 6974 4412
rect 7026 4410 7042 4462
rect 6250 4404 6304 4410
rect 6974 4404 7026 4410
rect 5934 4296 5986 4302
rect 6580 4256 6586 4308
rect 6638 4256 6644 4308
rect 5934 4238 5986 4244
rect 3979 4152 4673 4191
rect 4862 4182 4914 4188
rect 2818 4132 2824 4136
rect 2509 4116 2587 4118
rect 2522 4114 2574 4116
rect 2768 4092 2812 4132
rect 5015 4184 5067 4190
rect 4914 4142 5015 4171
rect 42 2234 110 3416
rect 42 1028 110 2166
rect 42 951 110 960
rect 144 4014 212 4023
rect 144 2778 212 3946
rect 274 3865 329 4054
rect 372 4018 378 4074
rect 434 4018 440 4074
rect 274 3859 332 3865
rect 274 3805 278 3859
rect 277 3684 332 3805
rect 378 3846 434 4018
rect 1324 3991 1960 4044
rect 1324 3989 1374 3991
rect 1430 3989 1454 3991
rect 1510 3989 1534 3991
rect 1590 3989 1614 3991
rect 1670 3989 1694 3991
rect 1750 3989 1774 3991
rect 1830 3989 1854 3991
rect 1910 3989 1960 3991
rect 1324 3937 1360 3989
rect 1604 3937 1614 3989
rect 1670 3937 1680 3989
rect 1924 3937 1960 3989
rect 1324 3935 1374 3937
rect 1430 3935 1454 3937
rect 1510 3935 1534 3937
rect 1590 3935 1614 3937
rect 1670 3935 1694 3937
rect 1750 3935 1774 3937
rect 1830 3935 1854 3937
rect 1910 3935 1960 3937
rect 1324 3904 1960 3935
rect 3564 3857 3605 4128
rect 4862 4124 4914 4130
rect 5015 4126 5067 4132
rect 5202 4128 5243 4208
rect 5282 4128 5323 4208
rect 5362 4128 5403 4208
rect 5442 4128 5483 4208
rect 5522 4128 5563 4208
rect 5938 4192 5976 4238
rect 6596 4192 6630 4256
rect 5938 4152 6632 4192
rect 6820 4182 6872 4188
rect 6974 4184 7026 4190
rect 6872 4142 6974 4172
rect 3704 4002 4244 4044
rect 3704 3946 3746 4002
rect 3802 4000 3826 4002
rect 3882 4000 3906 4002
rect 3962 4000 3986 4002
rect 4042 4000 4066 4002
rect 4122 4000 4146 4002
rect 3808 3948 3820 4000
rect 3882 3948 3884 4000
rect 4064 3948 4066 4000
rect 4128 3948 4140 4000
rect 3802 3946 3826 3948
rect 3882 3946 3906 3948
rect 3962 3946 3986 3948
rect 4042 3946 4066 3948
rect 4122 3946 4146 3948
rect 4202 3946 4244 4002
rect 4546 3999 4552 4051
rect 4604 3999 4610 4051
rect 3704 3904 4244 3946
rect 3564 3851 3617 3857
rect 274 3059 329 3684
rect 378 3230 433 3846
rect 3564 3799 3565 3851
rect 4559 3835 4598 3999
rect 5122 3857 5164 4128
rect 5117 3851 5169 3857
rect 3564 3793 3617 3799
rect 5117 3793 5169 3799
rect 1348 3465 1880 3506
rect 1348 3409 1388 3465
rect 1444 3463 1468 3465
rect 1524 3463 1548 3465
rect 1604 3463 1628 3465
rect 1684 3463 1708 3465
rect 1764 3463 1788 3465
rect 1450 3411 1462 3463
rect 1524 3411 1526 3463
rect 1706 3411 1708 3463
rect 1770 3411 1782 3463
rect 1444 3409 1468 3411
rect 1524 3409 1548 3411
rect 1604 3409 1628 3411
rect 1684 3409 1708 3411
rect 1764 3409 1788 3411
rect 1844 3409 1880 3465
rect 560 3392 612 3398
rect 700 3390 756 3396
rect 612 3388 976 3390
rect 612 3340 702 3388
rect 560 3336 702 3340
rect 754 3336 976 3388
rect 1348 3366 1880 3409
rect 2759 3348 2827 3356
rect 560 3334 1268 3336
rect 700 3328 756 3334
rect 920 3328 1268 3334
rect 2759 3328 2769 3348
rect 920 3296 2769 3328
rect 2821 3296 2827 3348
rect 920 3284 2827 3296
rect 920 3280 1268 3284
rect 852 3238 904 3244
rect 372 3175 378 3230
rect 433 3175 439 3230
rect 1396 3239 2851 3248
rect 3268 3243 3320 3249
rect 1396 3234 3268 3239
rect 904 3204 3268 3234
rect 904 3190 1440 3204
rect 2851 3195 3268 3204
rect 852 3180 904 3186
rect 3268 3185 3320 3191
rect 1930 3158 1990 3169
rect 1004 3146 1056 3152
rect 1930 3147 1932 3158
rect 1056 3135 1242 3142
rect 1599 3135 1932 3147
rect 1056 3113 1932 3135
rect 1056 3101 1633 3113
rect 1930 3102 1932 3113
rect 1988 3147 1990 3158
rect 1988 3113 1991 3147
rect 1988 3102 1990 3113
rect 1056 3098 1242 3101
rect 1004 3088 1056 3094
rect 1930 3091 1990 3102
rect 3564 3083 3605 3793
rect 5029 3629 5035 3681
rect 5087 3629 5093 3681
rect 4744 3562 4796 3568
rect 5047 3556 5075 3629
rect 4796 3517 5075 3556
rect 3724 3464 4264 3506
rect 4744 3504 4796 3510
rect 3724 3408 3766 3464
rect 3822 3462 3846 3464
rect 3902 3462 3926 3464
rect 3982 3462 4006 3464
rect 4062 3462 4086 3464
rect 4142 3462 4166 3464
rect 3828 3410 3840 3462
rect 3902 3410 3904 3462
rect 4084 3410 4086 3462
rect 4148 3410 4160 3462
rect 3822 3408 3846 3410
rect 3902 3408 3926 3410
rect 3982 3408 4006 3410
rect 4062 3408 4086 3410
rect 4142 3408 4166 3410
rect 4222 3408 4264 3464
rect 3724 3366 4264 3408
rect 4291 3237 4346 3243
rect 5016 3237 5068 3240
rect 4291 3235 5084 3237
rect 4291 3183 4292 3235
rect 4344 3234 5084 3235
rect 4344 3183 5016 3234
rect 4291 3182 5016 3183
rect 5068 3182 5084 3234
rect 4291 3176 4346 3182
rect 5016 3176 5068 3182
rect 3561 3077 3613 3083
rect 1154 3059 1209 3065
rect 274 3057 1209 3059
rect 274 3005 1155 3057
rect 1207 3005 1209 3057
rect 274 3004 1209 3005
rect 1154 2998 1209 3004
rect 1754 3060 1814 3066
rect 2267 3060 2325 3069
rect 1754 3057 2325 3060
rect 2838 3057 2898 3062
rect 1754 3056 2898 3057
rect 1754 3004 1758 3056
rect 1810 3054 2908 3056
rect 1810 3004 2270 3054
rect 1754 3002 2270 3004
rect 2322 3052 2908 3054
rect 2322 3002 2842 3052
rect 1754 3000 2842 3002
rect 2894 3000 2908 3052
rect 1754 2994 1814 3000
rect 2267 2999 2908 3000
rect 2267 2987 2325 2999
rect 2838 2996 2908 2999
rect 3262 2998 3268 3050
rect 3320 2998 3326 3050
rect 3976 3068 4028 3074
rect 3561 3019 3613 3025
rect 3975 3019 3976 3062
rect 2838 2990 2898 2996
rect 2768 2956 2816 2960
rect 378 2945 433 2951
rect 1248 2946 1300 2952
rect 433 2942 619 2945
rect 433 2898 1248 2942
rect 433 2890 619 2898
rect 2020 2946 2072 2952
rect 2522 2948 2574 2950
rect 1300 2898 2020 2942
rect 378 2884 433 2890
rect 1248 2888 1300 2894
rect 2020 2888 2072 2894
rect 2509 2946 2587 2948
rect 2509 2890 2520 2946
rect 2576 2890 2587 2946
rect 2760 2904 2766 2956
rect 2818 2952 2824 2956
rect 3270 2952 3314 2998
rect 3564 2980 3605 3019
rect 4622 3027 4628 3079
rect 4680 3027 4686 3079
rect 3976 3010 4028 3016
rect 2818 2908 3314 2952
rect 3979 2963 4018 3010
rect 4637 2963 4671 3027
rect 5122 2980 5164 3793
rect 5202 3083 5244 4128
rect 5197 3077 5249 3083
rect 5197 3019 5249 3025
rect 5202 2980 5244 3019
rect 5282 2980 5324 4128
rect 5362 2980 5404 4128
rect 5442 2980 5484 4128
rect 5522 2980 5564 4128
rect 6820 4124 6872 4130
rect 6974 4126 7026 4132
rect 5662 4002 6202 4044
rect 5662 3946 5704 4002
rect 5760 4000 5784 4002
rect 5840 4000 5864 4002
rect 5920 4000 5944 4002
rect 6000 4000 6024 4002
rect 6080 4000 6104 4002
rect 5766 3948 5778 4000
rect 5840 3948 5842 4000
rect 6022 3948 6024 4000
rect 6086 3948 6098 4000
rect 5760 3946 5784 3948
rect 5840 3946 5864 3948
rect 5920 3946 5944 3948
rect 6000 3946 6024 3948
rect 6080 3946 6104 3948
rect 6160 3946 6202 4002
rect 6504 4000 6510 4052
rect 6562 4000 6568 4052
rect 5662 3904 6202 3946
rect 6518 3836 6556 4000
rect 6523 3766 6553 3836
rect 6506 3714 6512 3766
rect 6564 3714 6570 3766
rect 6843 3562 6895 3568
rect 6895 3517 7150 3556
rect 5682 3464 6222 3506
rect 6843 3504 6895 3510
rect 5682 3408 5724 3464
rect 5780 3462 5804 3464
rect 5860 3462 5884 3464
rect 5940 3462 5964 3464
rect 6020 3462 6044 3464
rect 6100 3462 6124 3464
rect 5786 3410 5798 3462
rect 5860 3410 5862 3462
rect 6042 3410 6044 3462
rect 6106 3410 6118 3462
rect 5780 3408 5804 3410
rect 5860 3408 5884 3410
rect 5940 3408 5964 3410
rect 6020 3408 6044 3410
rect 6100 3408 6124 3410
rect 6180 3408 6222 3464
rect 5682 3366 6222 3408
rect 6250 3238 6304 3244
rect 6974 3238 7026 3240
rect 6250 3236 7042 3238
rect 6302 3234 7042 3236
rect 6302 3184 6974 3234
rect 6250 3182 6974 3184
rect 7026 3182 7042 3234
rect 6250 3176 6304 3182
rect 6974 3176 7026 3182
rect 5934 3068 5986 3074
rect 6580 3028 6586 3080
rect 6638 3028 6644 3080
rect 5934 3010 5986 3016
rect 3979 2924 4673 2963
rect 4862 2954 4914 2960
rect 2818 2904 2824 2908
rect 2509 2888 2587 2890
rect 2522 2886 2574 2888
rect 2768 2864 2812 2904
rect 5015 2956 5067 2962
rect 4914 2914 5015 2943
rect 144 1558 212 2710
rect 274 2637 329 2826
rect 372 2790 378 2846
rect 434 2790 440 2846
rect 274 2631 332 2637
rect 274 2577 278 2631
rect 277 2456 332 2577
rect 378 2618 434 2790
rect 1324 2763 1960 2816
rect 1324 2761 1374 2763
rect 1430 2761 1454 2763
rect 1510 2761 1534 2763
rect 1590 2761 1614 2763
rect 1670 2761 1694 2763
rect 1750 2761 1774 2763
rect 1830 2761 1854 2763
rect 1910 2761 1960 2763
rect 1324 2709 1360 2761
rect 1604 2709 1614 2761
rect 1670 2709 1680 2761
rect 1924 2709 1960 2761
rect 1324 2707 1374 2709
rect 1430 2707 1454 2709
rect 1510 2707 1534 2709
rect 1590 2707 1614 2709
rect 1670 2707 1694 2709
rect 1750 2707 1774 2709
rect 1830 2707 1854 2709
rect 1910 2707 1960 2709
rect 1324 2676 1960 2707
rect 3564 2629 3605 2900
rect 4862 2896 4914 2902
rect 5015 2898 5067 2904
rect 5122 2900 5163 2980
rect 5282 2900 5323 2980
rect 5362 2900 5403 2980
rect 5442 2900 5483 2980
rect 5522 2900 5563 2980
rect 5938 2964 5976 3010
rect 6596 2964 6630 3028
rect 5938 2924 6632 2964
rect 6820 2954 6872 2960
rect 6974 2956 7026 2962
rect 6872 2914 6974 2944
rect 3704 2774 4244 2816
rect 3704 2718 3746 2774
rect 3802 2772 3826 2774
rect 3882 2772 3906 2774
rect 3962 2772 3986 2774
rect 4042 2772 4066 2774
rect 4122 2772 4146 2774
rect 3808 2720 3820 2772
rect 3882 2720 3884 2772
rect 4064 2720 4066 2772
rect 4128 2720 4140 2772
rect 3802 2718 3826 2720
rect 3882 2718 3906 2720
rect 3962 2718 3986 2720
rect 4042 2718 4066 2720
rect 4122 2718 4146 2720
rect 4202 2718 4244 2774
rect 4546 2771 4552 2823
rect 4604 2771 4610 2823
rect 3704 2676 4244 2718
rect 3564 2623 3617 2629
rect 274 1831 329 2456
rect 378 2002 433 2618
rect 3564 2571 3565 2623
rect 4559 2607 4598 2771
rect 3564 2565 3617 2571
rect 1348 2237 1880 2278
rect 1348 2181 1388 2237
rect 1444 2235 1468 2237
rect 1524 2235 1548 2237
rect 1604 2235 1628 2237
rect 1684 2235 1708 2237
rect 1764 2235 1788 2237
rect 1450 2183 1462 2235
rect 1524 2183 1526 2235
rect 1706 2183 1708 2235
rect 1770 2183 1782 2235
rect 1444 2181 1468 2183
rect 1524 2181 1548 2183
rect 1604 2181 1628 2183
rect 1684 2181 1708 2183
rect 1764 2181 1788 2183
rect 1844 2181 1880 2237
rect 560 2164 612 2170
rect 700 2162 756 2168
rect 612 2160 976 2162
rect 612 2112 702 2160
rect 560 2108 702 2112
rect 754 2108 976 2160
rect 1348 2138 1880 2181
rect 2759 2120 2827 2128
rect 560 2106 1268 2108
rect 700 2100 756 2106
rect 920 2100 1268 2106
rect 2759 2100 2769 2120
rect 920 2068 2769 2100
rect 2821 2068 2827 2120
rect 920 2056 2827 2068
rect 920 2052 1268 2056
rect 852 2010 904 2016
rect 372 1947 378 2002
rect 433 1947 439 2002
rect 1396 2011 2851 2020
rect 3268 2015 3320 2021
rect 1396 2006 3268 2011
rect 904 1976 3268 2006
rect 904 1962 1440 1976
rect 2851 1967 3268 1976
rect 852 1952 904 1958
rect 3268 1957 3320 1963
rect 1930 1930 1990 1941
rect 1004 1918 1056 1924
rect 1930 1919 1932 1930
rect 1056 1907 1242 1914
rect 1599 1907 1932 1919
rect 1056 1885 1932 1907
rect 1056 1873 1633 1885
rect 1930 1874 1932 1885
rect 1988 1919 1990 1930
rect 1988 1885 1991 1919
rect 1988 1874 1990 1885
rect 1056 1870 1242 1873
rect 1004 1860 1056 1866
rect 1930 1863 1990 1874
rect 3564 1855 3605 2565
rect 5023 2364 5029 2416
rect 5081 2364 5087 2416
rect 4744 2334 4796 2340
rect 5036 2328 5075 2364
rect 4796 2289 5075 2328
rect 3724 2236 4264 2278
rect 4744 2276 4796 2282
rect 3724 2180 3766 2236
rect 3822 2234 3846 2236
rect 3902 2234 3926 2236
rect 3982 2234 4006 2236
rect 4062 2234 4086 2236
rect 4142 2234 4166 2236
rect 3828 2182 3840 2234
rect 3902 2182 3904 2234
rect 4084 2182 4086 2234
rect 4148 2182 4160 2234
rect 3822 2180 3846 2182
rect 3902 2180 3926 2182
rect 3982 2180 4006 2182
rect 4062 2180 4086 2182
rect 4142 2180 4166 2182
rect 4222 2180 4264 2236
rect 3724 2138 4264 2180
rect 4291 2009 4346 2015
rect 5016 2009 5068 2012
rect 4291 2007 5084 2009
rect 4291 1955 4292 2007
rect 4344 2006 5084 2007
rect 4344 1955 5016 2006
rect 4291 1954 5016 1955
rect 5068 1954 5084 2006
rect 4291 1948 4346 1954
rect 5016 1948 5068 1954
rect 5122 1855 5164 2900
rect 5202 2629 5244 2900
rect 5197 2623 5249 2629
rect 5197 2565 5249 2571
rect 3561 1849 3613 1855
rect 1154 1831 1209 1837
rect 274 1829 1209 1831
rect 274 1777 1155 1829
rect 1207 1777 1209 1829
rect 274 1776 1209 1777
rect 1154 1770 1209 1776
rect 1754 1832 1814 1838
rect 2267 1832 2325 1841
rect 1754 1829 2325 1832
rect 2838 1829 2898 1834
rect 1754 1828 2898 1829
rect 1754 1776 1758 1828
rect 1810 1826 2908 1828
rect 1810 1776 2270 1826
rect 1754 1774 2270 1776
rect 2322 1824 2908 1826
rect 2322 1774 2842 1824
rect 1754 1772 2842 1774
rect 2894 1772 2908 1824
rect 1754 1766 1814 1772
rect 2267 1771 2908 1772
rect 2267 1759 2325 1771
rect 2838 1768 2908 1771
rect 3262 1770 3268 1822
rect 3320 1770 3326 1822
rect 3976 1840 4028 1846
rect 3561 1791 3613 1797
rect 3975 1791 3976 1834
rect 2838 1762 2898 1768
rect 2768 1728 2816 1732
rect 378 1717 433 1723
rect 1248 1718 1300 1724
rect 433 1714 619 1717
rect 433 1670 1248 1714
rect 433 1662 619 1670
rect 2020 1718 2072 1724
rect 2522 1720 2574 1722
rect 1300 1670 2020 1714
rect 378 1656 433 1662
rect 1248 1660 1300 1666
rect 2020 1660 2072 1666
rect 2509 1718 2587 1720
rect 2509 1662 2520 1718
rect 2576 1662 2587 1718
rect 2760 1676 2766 1728
rect 2818 1724 2824 1728
rect 3270 1724 3314 1770
rect 3564 1752 3605 1791
rect 4622 1799 4628 1851
rect 4680 1799 4686 1851
rect 5117 1849 5169 1855
rect 3976 1782 4028 1788
rect 2818 1680 3314 1724
rect 3979 1735 4018 1782
rect 4637 1735 4671 1799
rect 5117 1791 5169 1797
rect 5122 1752 5164 1791
rect 5202 1752 5244 2565
rect 5282 1752 5324 2900
rect 5362 1752 5404 2900
rect 5442 1752 5484 2900
rect 5522 1752 5564 2900
rect 6820 2896 6872 2902
rect 6974 2898 7026 2904
rect 5662 2774 6202 2816
rect 5662 2718 5704 2774
rect 5760 2772 5784 2774
rect 5840 2772 5864 2774
rect 5920 2772 5944 2774
rect 6000 2772 6024 2774
rect 6080 2772 6104 2774
rect 5766 2720 5778 2772
rect 5840 2720 5842 2772
rect 6022 2720 6024 2772
rect 6086 2720 6098 2772
rect 5760 2718 5784 2720
rect 5840 2718 5864 2720
rect 5920 2718 5944 2720
rect 6000 2718 6024 2720
rect 6080 2718 6104 2720
rect 6160 2718 6202 2774
rect 6504 2772 6510 2824
rect 6562 2772 6568 2824
rect 5662 2676 6202 2718
rect 6518 2608 6556 2772
rect 7101 2484 7107 2536
rect 7159 2484 7165 2536
rect 6868 2334 6920 2340
rect 7119 2328 7147 2484
rect 6920 2289 7147 2328
rect 5682 2236 6222 2278
rect 6868 2276 6920 2282
rect 5682 2180 5724 2236
rect 5780 2234 5804 2236
rect 5860 2234 5884 2236
rect 5940 2234 5964 2236
rect 6020 2234 6044 2236
rect 6100 2234 6124 2236
rect 5786 2182 5798 2234
rect 5860 2182 5862 2234
rect 6042 2182 6044 2234
rect 6106 2182 6118 2234
rect 5780 2180 5804 2182
rect 5860 2180 5884 2182
rect 5940 2180 5964 2182
rect 6020 2180 6044 2182
rect 6100 2180 6124 2182
rect 6180 2180 6222 2236
rect 5682 2138 6222 2180
rect 6250 2010 6304 2016
rect 6974 2010 7026 2012
rect 6250 2008 7042 2010
rect 6302 2006 7042 2008
rect 6302 1956 6974 2006
rect 6250 1954 6974 1956
rect 7026 1954 7042 2006
rect 6250 1948 6304 1954
rect 6974 1948 7026 1954
rect 5934 1840 5986 1846
rect 6580 1800 6586 1852
rect 6638 1800 6644 1852
rect 5934 1782 5986 1788
rect 3979 1696 4673 1735
rect 4862 1726 4914 1732
rect 2818 1676 2824 1680
rect 2509 1660 2587 1662
rect 2522 1658 2574 1660
rect 2768 1636 2812 1676
rect 5015 1728 5067 1734
rect 4914 1686 5015 1715
rect 144 322 212 1490
rect 274 1409 329 1598
rect 372 1562 378 1618
rect 434 1562 440 1618
rect 274 1403 332 1409
rect 274 1349 278 1403
rect 277 1228 332 1349
rect 378 1390 434 1562
rect 1324 1535 1960 1588
rect 1324 1533 1374 1535
rect 1430 1533 1454 1535
rect 1510 1533 1534 1535
rect 1590 1533 1614 1535
rect 1670 1533 1694 1535
rect 1750 1533 1774 1535
rect 1830 1533 1854 1535
rect 1910 1533 1960 1535
rect 1324 1481 1360 1533
rect 1604 1481 1614 1533
rect 1670 1481 1680 1533
rect 1924 1481 1960 1533
rect 1324 1479 1374 1481
rect 1430 1479 1454 1481
rect 1510 1479 1534 1481
rect 1590 1479 1614 1481
rect 1670 1479 1694 1481
rect 1750 1479 1774 1481
rect 1830 1479 1854 1481
rect 1910 1479 1960 1481
rect 1324 1448 1960 1479
rect 3564 1401 3605 1672
rect 4862 1668 4914 1674
rect 5015 1670 5067 1676
rect 5202 1672 5243 1752
rect 5282 1672 5323 1752
rect 5362 1672 5403 1752
rect 5442 1672 5483 1752
rect 5522 1672 5563 1752
rect 5938 1736 5976 1782
rect 6596 1736 6630 1800
rect 5938 1696 6632 1736
rect 6820 1726 6872 1732
rect 6974 1728 7026 1734
rect 6872 1686 6974 1716
rect 3704 1546 4244 1588
rect 3704 1490 3746 1546
rect 3802 1544 3826 1546
rect 3882 1544 3906 1546
rect 3962 1544 3986 1546
rect 4042 1544 4066 1546
rect 4122 1544 4146 1546
rect 3808 1492 3820 1544
rect 3882 1492 3884 1544
rect 4064 1492 4066 1544
rect 4128 1492 4140 1544
rect 3802 1490 3826 1492
rect 3882 1490 3906 1492
rect 3962 1490 3986 1492
rect 4042 1490 4066 1492
rect 4122 1490 4146 1492
rect 4202 1490 4244 1546
rect 4546 1543 4552 1595
rect 4604 1543 4610 1595
rect 3704 1448 4244 1490
rect 3564 1395 3617 1401
rect 274 603 329 1228
rect 378 774 433 1390
rect 3564 1343 3565 1395
rect 4559 1379 4598 1543
rect 5122 1401 5164 1672
rect 5117 1395 5169 1401
rect 3564 1337 3617 1343
rect 5117 1337 5169 1343
rect 1348 1009 1880 1050
rect 1348 953 1388 1009
rect 1444 1007 1468 1009
rect 1524 1007 1548 1009
rect 1604 1007 1628 1009
rect 1684 1007 1708 1009
rect 1764 1007 1788 1009
rect 1450 955 1462 1007
rect 1524 955 1526 1007
rect 1706 955 1708 1007
rect 1770 955 1782 1007
rect 1444 953 1468 955
rect 1524 953 1548 955
rect 1604 953 1628 955
rect 1684 953 1708 955
rect 1764 953 1788 955
rect 1844 953 1880 1009
rect 560 936 612 942
rect 700 934 756 940
rect 612 932 976 934
rect 612 884 702 932
rect 560 880 702 884
rect 754 880 976 932
rect 1348 910 1880 953
rect 2759 892 2827 900
rect 560 878 1268 880
rect 700 872 756 878
rect 920 872 1268 878
rect 2759 872 2769 892
rect 920 840 2769 872
rect 2821 840 2827 892
rect 920 828 2827 840
rect 920 824 1268 828
rect 852 782 904 788
rect 372 719 378 774
rect 433 719 439 774
rect 1396 783 2851 792
rect 3268 787 3320 793
rect 1396 778 3268 783
rect 904 748 3268 778
rect 904 734 1440 748
rect 2851 739 3268 748
rect 852 724 904 730
rect 3268 729 3320 735
rect 1930 702 1990 713
rect 1004 690 1056 696
rect 1930 691 1932 702
rect 1056 679 1242 686
rect 1599 679 1932 691
rect 1056 657 1932 679
rect 1056 645 1633 657
rect 1930 646 1932 657
rect 1988 691 1990 702
rect 1988 657 1991 691
rect 1988 646 1990 657
rect 1056 642 1242 645
rect 1004 632 1056 638
rect 1930 635 1990 646
rect 3564 627 3605 1337
rect 5029 1173 5035 1225
rect 5087 1173 5093 1225
rect 4744 1106 4796 1112
rect 5047 1100 5075 1173
rect 5122 1142 5164 1337
rect 5202 1142 5244 1672
rect 5282 1142 5324 1672
rect 5362 1142 5404 1672
rect 5442 1142 5484 1672
rect 5522 1142 5564 1672
rect 6820 1668 6872 1674
rect 6974 1670 7026 1676
rect 5662 1546 6202 1588
rect 5662 1490 5704 1546
rect 5760 1544 5784 1546
rect 5840 1544 5864 1546
rect 5920 1544 5944 1546
rect 6000 1544 6024 1546
rect 6080 1544 6104 1546
rect 5766 1492 5778 1544
rect 5840 1492 5842 1544
rect 6022 1492 6024 1544
rect 6086 1492 6098 1544
rect 5760 1490 5784 1492
rect 5840 1490 5864 1492
rect 5920 1490 5944 1492
rect 6000 1490 6024 1492
rect 6080 1490 6104 1492
rect 6160 1490 6202 1546
rect 6504 1544 6510 1596
rect 6562 1544 6568 1596
rect 5662 1448 6202 1490
rect 6518 1380 6556 1544
rect 4796 1061 5075 1100
rect 3724 1008 4264 1050
rect 4744 1048 4796 1054
rect 3724 952 3766 1008
rect 3822 1006 3846 1008
rect 3902 1006 3926 1008
rect 3982 1006 4006 1008
rect 4062 1006 4086 1008
rect 4142 1006 4166 1008
rect 3828 954 3840 1006
rect 3902 954 3904 1006
rect 4084 954 4086 1006
rect 4148 954 4160 1006
rect 3822 952 3846 954
rect 3902 952 3926 954
rect 3982 952 4006 954
rect 4062 952 4086 954
rect 4142 952 4166 954
rect 4222 952 4264 1008
rect 3724 910 4264 952
rect 4291 781 4346 787
rect 5016 781 5068 784
rect 4291 779 5084 781
rect 4291 727 4292 779
rect 4344 778 5084 779
rect 4344 727 5016 778
rect 4291 726 5016 727
rect 5068 726 5084 778
rect 4291 720 4346 726
rect 5016 720 5068 726
rect 3561 621 3613 627
rect 1154 603 1209 609
rect 274 601 1209 603
rect 274 549 1155 601
rect 1207 549 1209 601
rect 274 548 1209 549
rect 1154 542 1209 548
rect 1754 604 1814 610
rect 2267 604 2325 613
rect 1754 601 2325 604
rect 2838 601 2898 606
rect 1754 600 2898 601
rect 1754 548 1758 600
rect 1810 598 2908 600
rect 1810 548 2270 598
rect 1754 546 2270 548
rect 2322 596 2908 598
rect 2322 546 2842 596
rect 1754 544 2842 546
rect 2894 544 2908 596
rect 1754 538 1814 544
rect 2267 543 2908 544
rect 2267 531 2325 543
rect 2838 540 2908 543
rect 3262 542 3268 594
rect 3320 542 3326 594
rect 3976 612 4028 618
rect 3561 563 3613 569
rect 3975 563 3976 606
rect 2838 534 2898 540
rect 2768 500 2816 504
rect 378 489 433 495
rect 1248 490 1300 496
rect 433 486 619 489
rect 433 442 1248 486
rect 433 434 619 442
rect 2020 490 2072 496
rect 2522 492 2574 494
rect 1300 442 2020 486
rect 378 428 433 434
rect 1248 432 1300 438
rect 2020 432 2072 438
rect 2509 490 2587 492
rect 2509 434 2520 490
rect 2576 434 2587 490
rect 2760 448 2766 500
rect 2818 496 2824 500
rect 3270 496 3314 542
rect 3564 524 3605 563
rect 4622 571 4628 623
rect 4680 571 4686 623
rect 3976 554 4028 560
rect 2818 452 3314 496
rect 3979 507 4018 554
rect 4637 507 4671 571
rect 3979 468 4673 507
rect 4862 498 4914 504
rect 2818 448 2824 452
rect 2509 432 2587 434
rect 2522 430 2574 432
rect 2768 408 2812 448
rect 5015 500 5067 506
rect 4914 458 5015 487
rect 144 245 212 254
rect 274 181 329 370
rect 372 334 378 390
rect 434 334 440 390
rect 274 175 332 181
rect 274 121 278 175
rect 277 0 332 121
rect 378 162 434 334
rect 1324 307 1960 360
rect 1324 305 1374 307
rect 1430 305 1454 307
rect 1510 305 1534 307
rect 1590 305 1614 307
rect 1670 305 1694 307
rect 1750 305 1774 307
rect 1830 305 1854 307
rect 1910 305 1960 307
rect 1324 253 1360 305
rect 1604 253 1614 305
rect 1670 253 1680 305
rect 1924 253 1960 305
rect 1324 251 1374 253
rect 1430 251 1454 253
rect 1510 251 1534 253
rect 1590 251 1614 253
rect 1670 251 1694 253
rect 1750 251 1774 253
rect 1830 251 1854 253
rect 1910 251 1960 253
rect 1324 220 1960 251
rect 3564 173 3605 444
rect 4862 440 4914 446
rect 5015 442 5067 448
rect 3704 318 4244 360
rect 3704 262 3746 318
rect 3802 316 3826 318
rect 3882 316 3906 318
rect 3962 316 3986 318
rect 4042 316 4066 318
rect 4122 316 4146 318
rect 3808 264 3820 316
rect 3882 264 3884 316
rect 4064 264 4066 316
rect 4128 264 4140 316
rect 3802 262 3826 264
rect 3882 262 3906 264
rect 3962 262 3986 264
rect 4042 262 4066 264
rect 4122 262 4146 264
rect 4202 262 4244 318
rect 4546 315 4552 367
rect 4604 315 4610 367
rect 3704 220 4244 262
rect 3564 167 3617 173
rect 378 0 433 162
rect 3564 115 3565 167
rect 4559 151 4598 315
rect 3564 109 3617 115
rect 3564 0 3605 109
<< via2 >>
rect 42 4622 110 4690
rect 1388 4691 1444 4693
rect 1468 4691 1524 4693
rect 1548 4691 1604 4693
rect 1628 4691 1684 4693
rect 1708 4691 1764 4693
rect 1788 4691 1844 4693
rect 1388 4639 1398 4691
rect 1398 4639 1444 4691
rect 1468 4639 1514 4691
rect 1514 4639 1524 4691
rect 1548 4639 1578 4691
rect 1578 4639 1590 4691
rect 1590 4639 1604 4691
rect 1628 4639 1642 4691
rect 1642 4639 1654 4691
rect 1654 4639 1684 4691
rect 1708 4639 1718 4691
rect 1718 4639 1764 4691
rect 1788 4639 1834 4691
rect 1834 4639 1844 4691
rect 1388 4637 1444 4639
rect 1468 4637 1524 4639
rect 1548 4637 1604 4639
rect 1628 4637 1684 4639
rect 1708 4637 1764 4639
rect 1788 4637 1844 4639
rect 1932 4385 1988 4386
rect 1932 4333 1935 4385
rect 1935 4333 1987 4385
rect 1987 4333 1988 4385
rect 1932 4330 1988 4333
rect 3766 4690 3822 4692
rect 3846 4690 3902 4692
rect 3926 4690 3982 4692
rect 4006 4690 4062 4692
rect 4086 4690 4142 4692
rect 4166 4690 4222 4692
rect 3766 4638 3776 4690
rect 3776 4638 3822 4690
rect 3846 4638 3892 4690
rect 3892 4638 3902 4690
rect 3926 4638 3956 4690
rect 3956 4638 3968 4690
rect 3968 4638 3982 4690
rect 4006 4638 4020 4690
rect 4020 4638 4032 4690
rect 4032 4638 4062 4690
rect 4086 4638 4096 4690
rect 4096 4638 4142 4690
rect 4166 4638 4212 4690
rect 4212 4638 4222 4690
rect 3766 4636 3822 4638
rect 3846 4636 3902 4638
rect 3926 4636 3982 4638
rect 4006 4636 4062 4638
rect 4086 4636 4142 4638
rect 4166 4636 4222 4638
rect 2520 4172 2576 4174
rect 2520 4120 2522 4172
rect 2522 4120 2574 4172
rect 2574 4120 2576 4172
rect 2520 4118 2576 4120
rect 5724 4690 5780 4692
rect 5804 4690 5860 4692
rect 5884 4690 5940 4692
rect 5964 4690 6020 4692
rect 6044 4690 6100 4692
rect 6124 4690 6180 4692
rect 5724 4638 5734 4690
rect 5734 4638 5780 4690
rect 5804 4638 5850 4690
rect 5850 4638 5860 4690
rect 5884 4638 5914 4690
rect 5914 4638 5926 4690
rect 5926 4638 5940 4690
rect 5964 4638 5978 4690
rect 5978 4638 5990 4690
rect 5990 4638 6020 4690
rect 6044 4638 6054 4690
rect 6054 4638 6100 4690
rect 6124 4638 6170 4690
rect 6170 4638 6180 4690
rect 5724 4636 5780 4638
rect 5804 4636 5860 4638
rect 5884 4636 5940 4638
rect 5964 4636 6020 4638
rect 6044 4636 6100 4638
rect 6124 4636 6180 4638
rect 42 3416 110 3484
rect 42 2166 110 2234
rect 42 960 110 1028
rect 144 3946 212 4014
rect 1374 3989 1430 3991
rect 1454 3989 1510 3991
rect 1534 3989 1590 3991
rect 1614 3989 1670 3991
rect 1694 3989 1750 3991
rect 1774 3989 1830 3991
rect 1854 3989 1910 3991
rect 1374 3937 1412 3989
rect 1412 3937 1424 3989
rect 1424 3937 1430 3989
rect 1454 3937 1476 3989
rect 1476 3937 1488 3989
rect 1488 3937 1510 3989
rect 1534 3937 1540 3989
rect 1540 3937 1552 3989
rect 1552 3937 1590 3989
rect 1614 3937 1616 3989
rect 1616 3937 1668 3989
rect 1668 3937 1670 3989
rect 1694 3937 1732 3989
rect 1732 3937 1744 3989
rect 1744 3937 1750 3989
rect 1774 3937 1796 3989
rect 1796 3937 1808 3989
rect 1808 3937 1830 3989
rect 1854 3937 1860 3989
rect 1860 3937 1872 3989
rect 1872 3937 1910 3989
rect 1374 3935 1430 3937
rect 1454 3935 1510 3937
rect 1534 3935 1590 3937
rect 1614 3935 1670 3937
rect 1694 3935 1750 3937
rect 1774 3935 1830 3937
rect 1854 3935 1910 3937
rect 3746 4000 3802 4002
rect 3826 4000 3882 4002
rect 3906 4000 3962 4002
rect 3986 4000 4042 4002
rect 4066 4000 4122 4002
rect 4146 4000 4202 4002
rect 3746 3948 3756 4000
rect 3756 3948 3802 4000
rect 3826 3948 3872 4000
rect 3872 3948 3882 4000
rect 3906 3948 3936 4000
rect 3936 3948 3948 4000
rect 3948 3948 3962 4000
rect 3986 3948 4000 4000
rect 4000 3948 4012 4000
rect 4012 3948 4042 4000
rect 4066 3948 4076 4000
rect 4076 3948 4122 4000
rect 4146 3948 4192 4000
rect 4192 3948 4202 4000
rect 3746 3946 3802 3948
rect 3826 3946 3882 3948
rect 3906 3946 3962 3948
rect 3986 3946 4042 3948
rect 4066 3946 4122 3948
rect 4146 3946 4202 3948
rect 1388 3463 1444 3465
rect 1468 3463 1524 3465
rect 1548 3463 1604 3465
rect 1628 3463 1684 3465
rect 1708 3463 1764 3465
rect 1788 3463 1844 3465
rect 1388 3411 1398 3463
rect 1398 3411 1444 3463
rect 1468 3411 1514 3463
rect 1514 3411 1524 3463
rect 1548 3411 1578 3463
rect 1578 3411 1590 3463
rect 1590 3411 1604 3463
rect 1628 3411 1642 3463
rect 1642 3411 1654 3463
rect 1654 3411 1684 3463
rect 1708 3411 1718 3463
rect 1718 3411 1764 3463
rect 1788 3411 1834 3463
rect 1834 3411 1844 3463
rect 1388 3409 1444 3411
rect 1468 3409 1524 3411
rect 1548 3409 1604 3411
rect 1628 3409 1684 3411
rect 1708 3409 1764 3411
rect 1788 3409 1844 3411
rect 1932 3157 1988 3158
rect 1932 3105 1935 3157
rect 1935 3105 1987 3157
rect 1987 3105 1988 3157
rect 1932 3102 1988 3105
rect 3766 3462 3822 3464
rect 3846 3462 3902 3464
rect 3926 3462 3982 3464
rect 4006 3462 4062 3464
rect 4086 3462 4142 3464
rect 4166 3462 4222 3464
rect 3766 3410 3776 3462
rect 3776 3410 3822 3462
rect 3846 3410 3892 3462
rect 3892 3410 3902 3462
rect 3926 3410 3956 3462
rect 3956 3410 3968 3462
rect 3968 3410 3982 3462
rect 4006 3410 4020 3462
rect 4020 3410 4032 3462
rect 4032 3410 4062 3462
rect 4086 3410 4096 3462
rect 4096 3410 4142 3462
rect 4166 3410 4212 3462
rect 4212 3410 4222 3462
rect 3766 3408 3822 3410
rect 3846 3408 3902 3410
rect 3926 3408 3982 3410
rect 4006 3408 4062 3410
rect 4086 3408 4142 3410
rect 4166 3408 4222 3410
rect 2520 2944 2576 2946
rect 2520 2892 2522 2944
rect 2522 2892 2574 2944
rect 2574 2892 2576 2944
rect 2520 2890 2576 2892
rect 5704 4000 5760 4002
rect 5784 4000 5840 4002
rect 5864 4000 5920 4002
rect 5944 4000 6000 4002
rect 6024 4000 6080 4002
rect 6104 4000 6160 4002
rect 5704 3948 5714 4000
rect 5714 3948 5760 4000
rect 5784 3948 5830 4000
rect 5830 3948 5840 4000
rect 5864 3948 5894 4000
rect 5894 3948 5906 4000
rect 5906 3948 5920 4000
rect 5944 3948 5958 4000
rect 5958 3948 5970 4000
rect 5970 3948 6000 4000
rect 6024 3948 6034 4000
rect 6034 3948 6080 4000
rect 6104 3948 6150 4000
rect 6150 3948 6160 4000
rect 5704 3946 5760 3948
rect 5784 3946 5840 3948
rect 5864 3946 5920 3948
rect 5944 3946 6000 3948
rect 6024 3946 6080 3948
rect 6104 3946 6160 3948
rect 5724 3462 5780 3464
rect 5804 3462 5860 3464
rect 5884 3462 5940 3464
rect 5964 3462 6020 3464
rect 6044 3462 6100 3464
rect 6124 3462 6180 3464
rect 5724 3410 5734 3462
rect 5734 3410 5780 3462
rect 5804 3410 5850 3462
rect 5850 3410 5860 3462
rect 5884 3410 5914 3462
rect 5914 3410 5926 3462
rect 5926 3410 5940 3462
rect 5964 3410 5978 3462
rect 5978 3410 5990 3462
rect 5990 3410 6020 3462
rect 6044 3410 6054 3462
rect 6054 3410 6100 3462
rect 6124 3410 6170 3462
rect 6170 3410 6180 3462
rect 5724 3408 5780 3410
rect 5804 3408 5860 3410
rect 5884 3408 5940 3410
rect 5964 3408 6020 3410
rect 6044 3408 6100 3410
rect 6124 3408 6180 3410
rect 144 2710 212 2778
rect 1374 2761 1430 2763
rect 1454 2761 1510 2763
rect 1534 2761 1590 2763
rect 1614 2761 1670 2763
rect 1694 2761 1750 2763
rect 1774 2761 1830 2763
rect 1854 2761 1910 2763
rect 1374 2709 1412 2761
rect 1412 2709 1424 2761
rect 1424 2709 1430 2761
rect 1454 2709 1476 2761
rect 1476 2709 1488 2761
rect 1488 2709 1510 2761
rect 1534 2709 1540 2761
rect 1540 2709 1552 2761
rect 1552 2709 1590 2761
rect 1614 2709 1616 2761
rect 1616 2709 1668 2761
rect 1668 2709 1670 2761
rect 1694 2709 1732 2761
rect 1732 2709 1744 2761
rect 1744 2709 1750 2761
rect 1774 2709 1796 2761
rect 1796 2709 1808 2761
rect 1808 2709 1830 2761
rect 1854 2709 1860 2761
rect 1860 2709 1872 2761
rect 1872 2709 1910 2761
rect 1374 2707 1430 2709
rect 1454 2707 1510 2709
rect 1534 2707 1590 2709
rect 1614 2707 1670 2709
rect 1694 2707 1750 2709
rect 1774 2707 1830 2709
rect 1854 2707 1910 2709
rect 3746 2772 3802 2774
rect 3826 2772 3882 2774
rect 3906 2772 3962 2774
rect 3986 2772 4042 2774
rect 4066 2772 4122 2774
rect 4146 2772 4202 2774
rect 3746 2720 3756 2772
rect 3756 2720 3802 2772
rect 3826 2720 3872 2772
rect 3872 2720 3882 2772
rect 3906 2720 3936 2772
rect 3936 2720 3948 2772
rect 3948 2720 3962 2772
rect 3986 2720 4000 2772
rect 4000 2720 4012 2772
rect 4012 2720 4042 2772
rect 4066 2720 4076 2772
rect 4076 2720 4122 2772
rect 4146 2720 4192 2772
rect 4192 2720 4202 2772
rect 3746 2718 3802 2720
rect 3826 2718 3882 2720
rect 3906 2718 3962 2720
rect 3986 2718 4042 2720
rect 4066 2718 4122 2720
rect 4146 2718 4202 2720
rect 1388 2235 1444 2237
rect 1468 2235 1524 2237
rect 1548 2235 1604 2237
rect 1628 2235 1684 2237
rect 1708 2235 1764 2237
rect 1788 2235 1844 2237
rect 1388 2183 1398 2235
rect 1398 2183 1444 2235
rect 1468 2183 1514 2235
rect 1514 2183 1524 2235
rect 1548 2183 1578 2235
rect 1578 2183 1590 2235
rect 1590 2183 1604 2235
rect 1628 2183 1642 2235
rect 1642 2183 1654 2235
rect 1654 2183 1684 2235
rect 1708 2183 1718 2235
rect 1718 2183 1764 2235
rect 1788 2183 1834 2235
rect 1834 2183 1844 2235
rect 1388 2181 1444 2183
rect 1468 2181 1524 2183
rect 1548 2181 1604 2183
rect 1628 2181 1684 2183
rect 1708 2181 1764 2183
rect 1788 2181 1844 2183
rect 1932 1929 1988 1930
rect 1932 1877 1935 1929
rect 1935 1877 1987 1929
rect 1987 1877 1988 1929
rect 1932 1874 1988 1877
rect 3766 2234 3822 2236
rect 3846 2234 3902 2236
rect 3926 2234 3982 2236
rect 4006 2234 4062 2236
rect 4086 2234 4142 2236
rect 4166 2234 4222 2236
rect 3766 2182 3776 2234
rect 3776 2182 3822 2234
rect 3846 2182 3892 2234
rect 3892 2182 3902 2234
rect 3926 2182 3956 2234
rect 3956 2182 3968 2234
rect 3968 2182 3982 2234
rect 4006 2182 4020 2234
rect 4020 2182 4032 2234
rect 4032 2182 4062 2234
rect 4086 2182 4096 2234
rect 4096 2182 4142 2234
rect 4166 2182 4212 2234
rect 4212 2182 4222 2234
rect 3766 2180 3822 2182
rect 3846 2180 3902 2182
rect 3926 2180 3982 2182
rect 4006 2180 4062 2182
rect 4086 2180 4142 2182
rect 4166 2180 4222 2182
rect 2520 1716 2576 1718
rect 2520 1664 2522 1716
rect 2522 1664 2574 1716
rect 2574 1664 2576 1716
rect 2520 1662 2576 1664
rect 5704 2772 5760 2774
rect 5784 2772 5840 2774
rect 5864 2772 5920 2774
rect 5944 2772 6000 2774
rect 6024 2772 6080 2774
rect 6104 2772 6160 2774
rect 5704 2720 5714 2772
rect 5714 2720 5760 2772
rect 5784 2720 5830 2772
rect 5830 2720 5840 2772
rect 5864 2720 5894 2772
rect 5894 2720 5906 2772
rect 5906 2720 5920 2772
rect 5944 2720 5958 2772
rect 5958 2720 5970 2772
rect 5970 2720 6000 2772
rect 6024 2720 6034 2772
rect 6034 2720 6080 2772
rect 6104 2720 6150 2772
rect 6150 2720 6160 2772
rect 5704 2718 5760 2720
rect 5784 2718 5840 2720
rect 5864 2718 5920 2720
rect 5944 2718 6000 2720
rect 6024 2718 6080 2720
rect 6104 2718 6160 2720
rect 5724 2234 5780 2236
rect 5804 2234 5860 2236
rect 5884 2234 5940 2236
rect 5964 2234 6020 2236
rect 6044 2234 6100 2236
rect 6124 2234 6180 2236
rect 5724 2182 5734 2234
rect 5734 2182 5780 2234
rect 5804 2182 5850 2234
rect 5850 2182 5860 2234
rect 5884 2182 5914 2234
rect 5914 2182 5926 2234
rect 5926 2182 5940 2234
rect 5964 2182 5978 2234
rect 5978 2182 5990 2234
rect 5990 2182 6020 2234
rect 6044 2182 6054 2234
rect 6054 2182 6100 2234
rect 6124 2182 6170 2234
rect 6170 2182 6180 2234
rect 5724 2180 5780 2182
rect 5804 2180 5860 2182
rect 5884 2180 5940 2182
rect 5964 2180 6020 2182
rect 6044 2180 6100 2182
rect 6124 2180 6180 2182
rect 144 1490 212 1558
rect 1374 1533 1430 1535
rect 1454 1533 1510 1535
rect 1534 1533 1590 1535
rect 1614 1533 1670 1535
rect 1694 1533 1750 1535
rect 1774 1533 1830 1535
rect 1854 1533 1910 1535
rect 1374 1481 1412 1533
rect 1412 1481 1424 1533
rect 1424 1481 1430 1533
rect 1454 1481 1476 1533
rect 1476 1481 1488 1533
rect 1488 1481 1510 1533
rect 1534 1481 1540 1533
rect 1540 1481 1552 1533
rect 1552 1481 1590 1533
rect 1614 1481 1616 1533
rect 1616 1481 1668 1533
rect 1668 1481 1670 1533
rect 1694 1481 1732 1533
rect 1732 1481 1744 1533
rect 1744 1481 1750 1533
rect 1774 1481 1796 1533
rect 1796 1481 1808 1533
rect 1808 1481 1830 1533
rect 1854 1481 1860 1533
rect 1860 1481 1872 1533
rect 1872 1481 1910 1533
rect 1374 1479 1430 1481
rect 1454 1479 1510 1481
rect 1534 1479 1590 1481
rect 1614 1479 1670 1481
rect 1694 1479 1750 1481
rect 1774 1479 1830 1481
rect 1854 1479 1910 1481
rect 3746 1544 3802 1546
rect 3826 1544 3882 1546
rect 3906 1544 3962 1546
rect 3986 1544 4042 1546
rect 4066 1544 4122 1546
rect 4146 1544 4202 1546
rect 3746 1492 3756 1544
rect 3756 1492 3802 1544
rect 3826 1492 3872 1544
rect 3872 1492 3882 1544
rect 3906 1492 3936 1544
rect 3936 1492 3948 1544
rect 3948 1492 3962 1544
rect 3986 1492 4000 1544
rect 4000 1492 4012 1544
rect 4012 1492 4042 1544
rect 4066 1492 4076 1544
rect 4076 1492 4122 1544
rect 4146 1492 4192 1544
rect 4192 1492 4202 1544
rect 3746 1490 3802 1492
rect 3826 1490 3882 1492
rect 3906 1490 3962 1492
rect 3986 1490 4042 1492
rect 4066 1490 4122 1492
rect 4146 1490 4202 1492
rect 1388 1007 1444 1009
rect 1468 1007 1524 1009
rect 1548 1007 1604 1009
rect 1628 1007 1684 1009
rect 1708 1007 1764 1009
rect 1788 1007 1844 1009
rect 1388 955 1398 1007
rect 1398 955 1444 1007
rect 1468 955 1514 1007
rect 1514 955 1524 1007
rect 1548 955 1578 1007
rect 1578 955 1590 1007
rect 1590 955 1604 1007
rect 1628 955 1642 1007
rect 1642 955 1654 1007
rect 1654 955 1684 1007
rect 1708 955 1718 1007
rect 1718 955 1764 1007
rect 1788 955 1834 1007
rect 1834 955 1844 1007
rect 1388 953 1444 955
rect 1468 953 1524 955
rect 1548 953 1604 955
rect 1628 953 1684 955
rect 1708 953 1764 955
rect 1788 953 1844 955
rect 1932 701 1988 702
rect 1932 649 1935 701
rect 1935 649 1987 701
rect 1987 649 1988 701
rect 1932 646 1988 649
rect 5704 1544 5760 1546
rect 5784 1544 5840 1546
rect 5864 1544 5920 1546
rect 5944 1544 6000 1546
rect 6024 1544 6080 1546
rect 6104 1544 6160 1546
rect 5704 1492 5714 1544
rect 5714 1492 5760 1544
rect 5784 1492 5830 1544
rect 5830 1492 5840 1544
rect 5864 1492 5894 1544
rect 5894 1492 5906 1544
rect 5906 1492 5920 1544
rect 5944 1492 5958 1544
rect 5958 1492 5970 1544
rect 5970 1492 6000 1544
rect 6024 1492 6034 1544
rect 6034 1492 6080 1544
rect 6104 1492 6150 1544
rect 6150 1492 6160 1544
rect 5704 1490 5760 1492
rect 5784 1490 5840 1492
rect 5864 1490 5920 1492
rect 5944 1490 6000 1492
rect 6024 1490 6080 1492
rect 6104 1490 6160 1492
rect 3766 1006 3822 1008
rect 3846 1006 3902 1008
rect 3926 1006 3982 1008
rect 4006 1006 4062 1008
rect 4086 1006 4142 1008
rect 4166 1006 4222 1008
rect 3766 954 3776 1006
rect 3776 954 3822 1006
rect 3846 954 3892 1006
rect 3892 954 3902 1006
rect 3926 954 3956 1006
rect 3956 954 3968 1006
rect 3968 954 3982 1006
rect 4006 954 4020 1006
rect 4020 954 4032 1006
rect 4032 954 4062 1006
rect 4086 954 4096 1006
rect 4096 954 4142 1006
rect 4166 954 4212 1006
rect 4212 954 4222 1006
rect 3766 952 3822 954
rect 3846 952 3902 954
rect 3926 952 3982 954
rect 4006 952 4062 954
rect 4086 952 4142 954
rect 4166 952 4222 954
rect 2520 488 2576 490
rect 2520 436 2522 488
rect 2522 436 2574 488
rect 2574 436 2576 488
rect 2520 434 2576 436
rect 144 254 212 322
rect 1374 305 1430 307
rect 1454 305 1510 307
rect 1534 305 1590 307
rect 1614 305 1670 307
rect 1694 305 1750 307
rect 1774 305 1830 307
rect 1854 305 1910 307
rect 1374 253 1412 305
rect 1412 253 1424 305
rect 1424 253 1430 305
rect 1454 253 1476 305
rect 1476 253 1488 305
rect 1488 253 1510 305
rect 1534 253 1540 305
rect 1540 253 1552 305
rect 1552 253 1590 305
rect 1614 253 1616 305
rect 1616 253 1668 305
rect 1668 253 1670 305
rect 1694 253 1732 305
rect 1732 253 1744 305
rect 1744 253 1750 305
rect 1774 253 1796 305
rect 1796 253 1808 305
rect 1808 253 1830 305
rect 1854 253 1860 305
rect 1860 253 1872 305
rect 1872 253 1910 305
rect 1374 251 1430 253
rect 1454 251 1510 253
rect 1534 251 1590 253
rect 1614 251 1670 253
rect 1694 251 1750 253
rect 1774 251 1830 253
rect 1854 251 1910 253
rect 3746 316 3802 318
rect 3826 316 3882 318
rect 3906 316 3962 318
rect 3986 316 4042 318
rect 4066 316 4122 318
rect 4146 316 4202 318
rect 3746 264 3756 316
rect 3756 264 3802 316
rect 3826 264 3872 316
rect 3872 264 3882 316
rect 3906 264 3936 316
rect 3936 264 3948 316
rect 3948 264 3962 316
rect 3986 264 4000 316
rect 4000 264 4012 316
rect 4012 264 4042 316
rect 4066 264 4076 316
rect 4076 264 4122 316
rect 4146 264 4192 316
rect 4192 264 4202 316
rect 3746 262 3802 264
rect 3826 262 3882 264
rect 3906 262 3962 264
rect 3986 262 4042 264
rect 4066 262 4122 264
rect 4146 262 4202 264
<< metal3 >>
rect -2 4693 7724 4734
rect -2 4690 1388 4693
rect -2 4622 42 4690
rect 110 4637 1388 4690
rect 1444 4637 1468 4693
rect 1524 4637 1548 4693
rect 1604 4637 1628 4693
rect 1684 4637 1708 4693
rect 1764 4637 1788 4693
rect 1844 4692 7724 4693
rect 1844 4637 3766 4692
rect 110 4636 3766 4637
rect 3822 4636 3846 4692
rect 3902 4636 3926 4692
rect 3982 4636 4006 4692
rect 4062 4636 4086 4692
rect 4142 4636 4166 4692
rect 4222 4636 5724 4692
rect 5780 4636 5804 4692
rect 5860 4636 5884 4692
rect 5940 4636 5964 4692
rect 6020 4636 6044 4692
rect 6100 4636 6124 4692
rect 6180 4636 7724 4692
rect 110 4622 7724 4636
rect -2 4594 7724 4622
rect 1925 4386 1995 4393
rect 1925 4330 1932 4386
rect 1988 4330 1995 4386
rect 1925 4323 1995 4330
rect 1930 4176 1990 4323
rect 2513 4176 2583 4181
rect 1930 4174 2583 4176
rect 1930 4118 2520 4174
rect 2576 4118 2583 4174
rect 1930 4116 2583 4118
rect 2513 4111 2583 4116
rect -2 4014 7724 4044
rect -2 3946 144 4014
rect 212 4002 7724 4014
rect 212 3991 3746 4002
rect 212 3946 1374 3991
rect -2 3935 1374 3946
rect 1430 3935 1454 3991
rect 1510 3935 1534 3991
rect 1590 3935 1614 3991
rect 1670 3935 1694 3991
rect 1750 3935 1774 3991
rect 1830 3935 1854 3991
rect 1910 3946 3746 3991
rect 3802 3946 3826 4002
rect 3882 3946 3906 4002
rect 3962 3946 3986 4002
rect 4042 3946 4066 4002
rect 4122 3946 4146 4002
rect 4202 3946 5704 4002
rect 5760 3946 5784 4002
rect 5840 3946 5864 4002
rect 5920 3946 5944 4002
rect 6000 3946 6024 4002
rect 6080 3946 6104 4002
rect 6160 3946 7724 4002
rect 1910 3935 7724 3946
rect -2 3904 7724 3935
rect -2 3484 7724 3506
rect -2 3416 42 3484
rect 110 3465 7724 3484
rect 110 3416 1388 3465
rect -2 3409 1388 3416
rect 1444 3409 1468 3465
rect 1524 3409 1548 3465
rect 1604 3409 1628 3465
rect 1684 3409 1708 3465
rect 1764 3409 1788 3465
rect 1844 3464 7724 3465
rect 1844 3409 3766 3464
rect -2 3408 3766 3409
rect 3822 3408 3846 3464
rect 3902 3408 3926 3464
rect 3982 3408 4006 3464
rect 4062 3408 4086 3464
rect 4142 3408 4166 3464
rect 4222 3408 5724 3464
rect 5780 3408 5804 3464
rect 5860 3408 5884 3464
rect 5940 3408 5964 3464
rect 6020 3408 6044 3464
rect 6100 3408 6124 3464
rect 6180 3408 7724 3464
rect -2 3366 7724 3408
rect 1925 3158 1995 3165
rect 1925 3102 1932 3158
rect 1988 3102 1995 3158
rect 1925 3095 1995 3102
rect 1930 2948 1990 3095
rect 2513 2948 2583 2953
rect 1930 2946 2583 2948
rect 1930 2890 2520 2946
rect 2576 2890 2583 2946
rect 1930 2888 2583 2890
rect 2513 2883 2583 2888
rect -2 2778 7724 2816
rect -2 2710 144 2778
rect 212 2774 7724 2778
rect 212 2763 3746 2774
rect 212 2710 1374 2763
rect -2 2707 1374 2710
rect 1430 2707 1454 2763
rect 1510 2707 1534 2763
rect 1590 2707 1614 2763
rect 1670 2707 1694 2763
rect 1750 2707 1774 2763
rect 1830 2707 1854 2763
rect 1910 2718 3746 2763
rect 3802 2718 3826 2774
rect 3882 2718 3906 2774
rect 3962 2718 3986 2774
rect 4042 2718 4066 2774
rect 4122 2718 4146 2774
rect 4202 2718 5704 2774
rect 5760 2718 5784 2774
rect 5840 2718 5864 2774
rect 5920 2718 5944 2774
rect 6000 2718 6024 2774
rect 6080 2718 6104 2774
rect 6160 2718 7724 2774
rect 1910 2707 7724 2718
rect -2 2676 7724 2707
rect -2 2237 7724 2278
rect -2 2234 1388 2237
rect -2 2166 42 2234
rect 110 2181 1388 2234
rect 1444 2181 1468 2237
rect 1524 2181 1548 2237
rect 1604 2181 1628 2237
rect 1684 2181 1708 2237
rect 1764 2181 1788 2237
rect 1844 2236 7724 2237
rect 1844 2181 3766 2236
rect 110 2180 3766 2181
rect 3822 2180 3846 2236
rect 3902 2180 3926 2236
rect 3982 2180 4006 2236
rect 4062 2180 4086 2236
rect 4142 2180 4166 2236
rect 4222 2180 5724 2236
rect 5780 2180 5804 2236
rect 5860 2180 5884 2236
rect 5940 2180 5964 2236
rect 6020 2180 6044 2236
rect 6100 2180 6124 2236
rect 6180 2180 7724 2236
rect 110 2166 7724 2180
rect -2 2138 7724 2166
rect 1925 1930 1995 1937
rect 1925 1874 1932 1930
rect 1988 1874 1995 1930
rect 1925 1867 1995 1874
rect 1930 1720 1990 1867
rect 2513 1720 2583 1725
rect 1930 1718 2583 1720
rect 1930 1662 2520 1718
rect 2576 1662 2583 1718
rect 1930 1660 2583 1662
rect 2513 1655 2583 1660
rect -2 1558 7724 1588
rect -2 1490 144 1558
rect 212 1546 7724 1558
rect 212 1535 3746 1546
rect 212 1490 1374 1535
rect -2 1479 1374 1490
rect 1430 1479 1454 1535
rect 1510 1479 1534 1535
rect 1590 1479 1614 1535
rect 1670 1479 1694 1535
rect 1750 1479 1774 1535
rect 1830 1479 1854 1535
rect 1910 1490 3746 1535
rect 3802 1490 3826 1546
rect 3882 1490 3906 1546
rect 3962 1490 3986 1546
rect 4042 1490 4066 1546
rect 4122 1490 4146 1546
rect 4202 1490 5704 1546
rect 5760 1490 5784 1546
rect 5840 1490 5864 1546
rect 5920 1490 5944 1546
rect 6000 1490 6024 1546
rect 6080 1490 6104 1546
rect 6160 1490 7724 1546
rect 1910 1479 7724 1490
rect -2 1448 7724 1479
rect -2 1028 7724 1050
rect -2 960 42 1028
rect 110 1009 7724 1028
rect 110 960 1388 1009
rect -2 953 1388 960
rect 1444 953 1468 1009
rect 1524 953 1548 1009
rect 1604 953 1628 1009
rect 1684 953 1708 1009
rect 1764 953 1788 1009
rect 1844 1008 7724 1009
rect 1844 953 3766 1008
rect -2 952 3766 953
rect 3822 952 3846 1008
rect 3902 952 3926 1008
rect 3982 952 4006 1008
rect 4062 952 4086 1008
rect 4142 952 4166 1008
rect 4222 952 7724 1008
rect -2 910 7724 952
rect 1925 702 1995 709
rect 1925 646 1932 702
rect 1988 646 1995 702
rect 1925 639 1995 646
rect 1930 492 1990 639
rect 2513 492 2583 497
rect 1930 490 2583 492
rect 1930 434 2520 490
rect 2576 434 2583 490
rect 1930 432 2583 434
rect 2513 427 2583 432
rect -2 322 7724 360
rect -2 254 144 322
rect 212 318 7724 322
rect 212 307 3746 318
rect 212 254 1374 307
rect -2 251 1374 254
rect 1430 251 1454 307
rect 1510 251 1534 307
rect 1590 251 1614 307
rect 1670 251 1694 307
rect 1750 251 1774 307
rect 1830 251 1854 307
rect 1910 262 3746 307
rect 3802 262 3826 318
rect 3882 262 3906 318
rect 3962 262 3986 318
rect 4042 262 4066 318
rect 4122 262 4146 318
rect 4202 262 7724 318
rect 1910 251 7724 262
rect -2 220 7724 251
<< labels >>
rlabel metal2 3574 8 3574 8 3 D1_BUF
rlabel metal2 5140 1282 5140 1282 3 D2_BUF
rlabel metal2 5212 1290 5212 1290 3 D3_BUF
flabel metal1 5562 3032 5582 3070 7 FreeSans 600 0 0 0 switch_n_3v3_0.DX
flabel metal1 5534 2578 5562 2616 7 FreeSans 600 0 0 0 switch_n_3v3_0.DX_BUF
flabel metal3 7052 3366 7082 3506 3 FreeSans 600 0 0 0 switch_n_3v3_0.VCC
flabel metal3 7052 2676 7082 2816 3 FreeSans 600 0 0 0 switch_n_3v3_0.VSS
flabel metal3 5072 2676 5102 2816 7 FreeSans 600 0 0 0 switch_n_3v3_0.VSS
flabel metal3 5072 3366 5102 3506 7 FreeSans 600 0 0 0 switch_n_3v3_0.VCC
flabel metal2 5142 3582 5142 3582 1 FreeSans 400 0 0 0 switch_n_3v3_0.D2
flabel metal2 5222 3586 5222 3586 1 FreeSans 400 0 0 0 switch_n_3v3_0.D3
flabel metal2 5304 3586 5304 3586 1 FreeSans 400 0 0 0 switch_n_3v3_0.D4
flabel metal2 5384 3588 5384 3588 1 FreeSans 400 0 0 0 switch_n_3v3_0.D5
flabel metal2 5462 3588 5462 3588 1 FreeSans 400 0 0 0 switch_n_3v3_0.D6
flabel metal2 5542 3586 5542 3586 1 FreeSans 400 0 0 0 switch_n_3v3_0.D7
flabel metal1 6516 3530 6556 3554 3 FreeSans 600 0 0 0 switch_n_3v3_0.VOUT
flabel metal2 6518 2608 6556 2632 7 FreeSans 600 0 0 0 switch_n_3v3_0.VOUT
flabel metal1 5872 3006 5872 3006 7 FreeSans 600 0 0 0 switch_n_3v3_0.DX_
flabel metal1 6908 2602 6936 2626 3 FreeSans 600 0 0 0 switch_n_3v3_0.VREFH
flabel metal1 6986 3526 7016 3546 3 FreeSans 600 0 0 0 switch_n_3v3_0.VREFL
rlabel metal3 18 2234 18 2234 7 3_bit_dac_0[0].VCC
rlabel metal3 26 1522 26 1522 7 3_bit_dac_0[0].VSS
rlabel metal2 302 2430 302 2430 7 3_bit_dac_0[0].D0
rlabel metal2 406 2432 406 2432 7 3_bit_dac_0[0].VREFL
rlabel metal2 304 20 304 20 7 3_bit_dac_0[0].D0_BUF
rlabel metal2 400 12 400 12 7 3_bit_dac_0[0].VREFH
rlabel metal2 3586 2450 3586 2450 7 3_bit_dac_0[0].D1
rlabel metal2 3586 12 3586 12 7 3_bit_dac_0[0].D1_BUF
rlabel metal2 5141 2436 5141 2436 7 3_bit_dac_0[0].D2
rlabel metal2 5141 1290 5141 1290 7 3_bit_dac_0[0].D2_BUF
rlabel metal2 7139 2310 7139 2310 7 3_bit_dac_0[0].VOUT
flabel metal1 5562 1804 5582 1842 7 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.DX
flabel metal1 5534 1350 5562 1388 7 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.DX_BUF
flabel metal3 7052 2138 7082 2278 3 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal3 7052 1448 7082 1588 3 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 1448 5102 1588 7 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 2138 5102 2278 7 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal2 5142 2354 5142 2354 1 FreeSans 400 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.D2
flabel metal2 5222 2358 5222 2358 1 FreeSans 400 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.D3
flabel metal2 5304 2358 5304 2358 1 FreeSans 400 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.D4
flabel metal2 5384 2360 5384 2360 1 FreeSans 400 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.D5
flabel metal2 5462 2360 5462 2360 1 FreeSans 400 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.D6
flabel metal2 5542 2358 5542 2358 1 FreeSans 400 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.D7
flabel metal1 6516 2302 6556 2326 3 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal2 6518 1380 6556 1404 7 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal1 5872 1778 5872 1778 7 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.DX_
flabel metal1 6908 1374 6936 1398 3 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VREFH
flabel metal1 6986 2298 7016 2318 3 FreeSans 600 0 0 0 3_bit_dac_0[0].switch_n_3v3_1.VREFL
rlabel metal3 148 991 148 991 7 3_bit_dac_0[0].2_bit_dac_0[0].VCC
rlabel metal3 166 286 166 286 7 3_bit_dac_0[0].2_bit_dac_0[0].VSS
rlabel metal2 295 1186 295 1186 7 3_bit_dac_0[0].2_bit_dac_0[0].D0
rlabel metal2 406 1186 406 1186 7 3_bit_dac_0[0].2_bit_dac_0[0].VREFL
rlabel metal2 301 36 301 36 7 3_bit_dac_0[0].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 19 409 19 7 3_bit_dac_0[0].2_bit_dac_0[0].VREFH
rlabel metal2 5056 1077 5056 1077 7 3_bit_dac_0[0].2_bit_dac_0[0].VOUT
rlabel metal2 3586 18 3586 18 7 3_bit_dac_0[0].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 1204 3584 1204 7 3_bit_dac_0[0].2_bit_dac_0[0].D1
flabel metal1 3492 966 3492 966 3 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 252 3478 252 3 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 662 1254 662 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 930 2662 930 3 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 756 1266 756 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 578 624 578 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 464 614 464 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 902 634 902 5 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 220 528 360 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 910 528 1050 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 575 3624 614 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 121 3603 160 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 910 5124 1050 3 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 220 5124 360 3 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 1074 4597 1099 3 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 151 4598 175 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 550 3914 550 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 220 3462 360 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 910 3462 1050 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 1107 4888 1107 1 FreeSans 480 0 0 40 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 141 5041 141 5 FreeSans 480 0 0 -40 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 2219 148 2219 7 3_bit_dac_0[0].2_bit_dac_0[1].VCC
rlabel metal3 166 1514 166 1514 7 3_bit_dac_0[0].2_bit_dac_0[1].VSS
rlabel metal2 295 2414 295 2414 7 3_bit_dac_0[0].2_bit_dac_0[1].D0
rlabel metal2 406 2414 406 2414 7 3_bit_dac_0[0].2_bit_dac_0[1].VREFL
rlabel metal2 301 1264 301 1264 7 3_bit_dac_0[0].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 1247 409 1247 7 3_bit_dac_0[0].2_bit_dac_0[1].VREFH
rlabel metal2 5056 2305 5056 2305 7 3_bit_dac_0[0].2_bit_dac_0[1].VOUT
rlabel metal2 3586 1246 3586 1246 7 3_bit_dac_0[0].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 2432 3584 2432 7 3_bit_dac_0[0].2_bit_dac_0[1].D1
flabel metal1 3492 2194 3492 2194 3 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 1480 3478 1480 3 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 1890 1254 1890 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 2158 2662 2158 3 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 1984 1266 1984 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 1806 624 1806 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 1692 614 1692 7 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 2130 634 2130 5 FreeSans 400 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 1448 528 1588 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 2138 528 2278 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 1803 3624 1842 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 1349 3603 1388 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 2138 5124 2278 3 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 1448 5124 1588 3 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 2302 4597 2327 3 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 1379 4598 1403 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 1778 3914 1778 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 1448 3462 1588 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 2138 3462 2278 7 FreeSans 600 0 0 0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 2335 4888 2335 1 FreeSans 480 0 0 40 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 1369 5041 1369 5 FreeSans 480 0 0 -40 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal3 18 4690 18 4690 7 3_bit_dac_0[1].VCC
rlabel metal3 26 3978 26 3978 7 3_bit_dac_0[1].VSS
rlabel metal2 302 4886 302 4886 7 3_bit_dac_0[1].D0
rlabel metal2 406 4888 406 4888 7 3_bit_dac_0[1].VREFL
rlabel metal2 304 2476 304 2476 7 3_bit_dac_0[1].D0_BUF
rlabel metal2 400 2468 400 2468 7 3_bit_dac_0[1].VREFH
rlabel metal2 3586 4906 3586 4906 7 3_bit_dac_0[1].D1
rlabel metal2 3586 2468 3586 2468 7 3_bit_dac_0[1].D1_BUF
rlabel metal2 5141 4892 5141 4892 7 3_bit_dac_0[1].D2
rlabel metal2 5141 3746 5141 3746 7 3_bit_dac_0[1].D2_BUF
rlabel metal2 7139 4766 7139 4766 7 3_bit_dac_0[1].VOUT
flabel metal1 5562 4260 5582 4298 7 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.DX
flabel metal1 5534 3806 5562 3844 7 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.DX_BUF
flabel metal3 7052 4594 7082 4734 3 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal3 7052 3904 7082 4044 3 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 3904 5102 4044 7 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 4594 5102 4734 7 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal2 5142 4810 5142 4810 1 FreeSans 400 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.D2
flabel metal2 5222 4814 5222 4814 1 FreeSans 400 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.D3
flabel metal2 5304 4814 5304 4814 1 FreeSans 400 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.D4
flabel metal2 5384 4816 5384 4816 1 FreeSans 400 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.D5
flabel metal2 5462 4816 5462 4816 1 FreeSans 400 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.D6
flabel metal2 5542 4814 5542 4814 1 FreeSans 400 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.D7
flabel metal1 6516 4758 6556 4782 3 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal2 6518 3836 6556 3860 7 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal1 5872 4234 5872 4234 7 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.DX_
flabel metal1 6908 3830 6936 3854 3 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VREFH
flabel metal1 6986 4754 7016 4774 3 FreeSans 600 0 0 0 3_bit_dac_0[1].switch_n_3v3_1.VREFL
rlabel metal3 148 3447 148 3447 7 3_bit_dac_0[1].2_bit_dac_0[0].VCC
rlabel metal3 166 2742 166 2742 7 3_bit_dac_0[1].2_bit_dac_0[0].VSS
rlabel metal2 295 3642 295 3642 7 3_bit_dac_0[1].2_bit_dac_0[0].D0
rlabel metal2 406 3642 406 3642 7 3_bit_dac_0[1].2_bit_dac_0[0].VREFL
rlabel metal2 301 2492 301 2492 7 3_bit_dac_0[1].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 2475 409 2475 7 3_bit_dac_0[1].2_bit_dac_0[0].VREFH
rlabel metal2 5056 3533 5056 3533 7 3_bit_dac_0[1].2_bit_dac_0[0].VOUT
rlabel metal2 3586 2474 3586 2474 7 3_bit_dac_0[1].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 3660 3584 3660 7 3_bit_dac_0[1].2_bit_dac_0[0].D1
flabel metal1 3492 3422 3492 3422 3 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 2708 3478 2708 3 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 3118 1254 3118 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 3386 2662 3386 3 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 3212 1266 3212 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 3034 624 3034 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 2920 614 2920 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 3358 634 3358 5 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 2676 528 2816 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 3366 528 3506 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 3031 3624 3070 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 2577 3603 2616 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 3366 5124 3506 3 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 2676 5124 2816 3 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 3530 4597 3555 3 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 2607 4598 2631 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 3006 3914 3006 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 2676 3462 2816 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 3366 3462 3506 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 3563 4888 3563 1 FreeSans 480 0 0 40 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 2597 5041 2597 5 FreeSans 480 0 0 -40 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 4675 148 4675 7 3_bit_dac_0[1].2_bit_dac_0[1].VCC
rlabel metal3 166 3970 166 3970 7 3_bit_dac_0[1].2_bit_dac_0[1].VSS
rlabel metal2 295 4870 295 4870 7 3_bit_dac_0[1].2_bit_dac_0[1].D0
rlabel metal2 406 4870 406 4870 7 3_bit_dac_0[1].2_bit_dac_0[1].VREFL
rlabel metal2 301 3720 301 3720 7 3_bit_dac_0[1].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 3703 409 3703 7 3_bit_dac_0[1].2_bit_dac_0[1].VREFH
rlabel metal2 5056 4761 5056 4761 7 3_bit_dac_0[1].2_bit_dac_0[1].VOUT
rlabel metal2 3586 3702 3586 3702 7 3_bit_dac_0[1].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 4888 3584 4888 7 3_bit_dac_0[1].2_bit_dac_0[1].D1
flabel metal1 3492 4650 3492 4650 3 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 3936 3478 3936 3 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 4346 1254 4346 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 4614 2662 4614 3 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 4440 1266 4440 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 4262 624 4262 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 4148 614 4148 7 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 4586 634 4586 5 FreeSans 400 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 3904 528 4044 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 4594 528 4734 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 4259 3624 4298 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 3805 3603 3844 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 4594 5124 4734 3 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 3904 5124 4044 3 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 4758 4597 4783 3 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 3835 4598 3859 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 4234 3914 4234 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 3904 3462 4044 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 4594 3462 4734 7 FreeSans 600 0 0 0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 4791 4888 4791 1 FreeSans 480 0 0 40 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 3825 5041 3825 5 FreeSans 480 0 0 -40 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
flabel metal2 s 294 4902 294 4902 0 FreeSans 1600 0 -1120 1120 D0
port 5 nsew signal input
flabel metal2 s 416 4906 416 4906 0 FreeSans 1600 0 3040 1120 VREFL
port 4 nsew signal input
flabel metal2 s 3580 4900 3580 4900 0 FreeSans 1600 0 0 1120 D1
port 6 nsew signal input
flabel metal2 s 5136 4908 5136 4908 0 FreeSans 1600 0 -1600 1120 D2
port 7 nsew signal input
flabel metal2 s 5234 4906 5234 4906 0 FreeSans 1600 0 800 1120 D3
port 8 nsew signal input
flabel metal2 s 74 4488 74 4488 0 FreeSans 1600 0 -3200 1280 VCC
port 1 nsew power bidirectional
flabel metal2 s 180 3756 180 3756 0 FreeSans 1600 0 -3200 0 VSS
port 2 nsew ground bidirectional
flabel metal2 s 416 10 416 10 5 FreeSans 1600 0 1920 -800 VREFH
port 3 s signal input
flabel metal2 6536 2662 6536 2662 5 FreeSans 1600 0 1920 -800 VOUT
port 9 s signal output
<< end >>
