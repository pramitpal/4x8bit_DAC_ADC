** sch_path: /foss/designs/Comparator/schematic/Edge_pursuit_comparator/EPC_testbench.sch
**.subckt EPC_testbench
x1 VCC VSS VINP VINN START OUT EPC
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice




V1 VSS 0 dc 0
V2 VCC 0 dc 3.3
V3 START 0 dc 3.3
V4 VINP 0 dc 1.65
V5 VINN 0 dc 1.9

.print tran format=raw file=EPC.raw  v(*)
.tran 1n 200n



**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Comparator/schematic/Edge_pursuit_comparator/EPC.sym # of
*+ pins=6
** sym_path: /foss/designs/Comparator/schematic/Edge_pursuit_comparator/EPC.sym
** sch_path: /foss/designs/Comparator/schematic/Edge_pursuit_comparator/EPC.sch
.subckt EPC VCC VSS VINP VINN START OUT
*.iopin VCC
*.opin OUT
*.ipin VINN
*.iopin VSS
*.ipin VINP
*.ipin START
x1 VCC VSS net8 VINP VINP net1 delay_cell
x2 VCC VSS net1 VINN VINN net2 delay_cell
x3 VCC VSS net2 VINP VINP net3 delay_cell
x4 VCC VSS net3 VINN VINN OUT delay_cell
x5 VCC VSS net4 VINP VINP net9 delay_cell
x6 VCC VSS net5 VINN VINN net4 delay_cell
x7 VCC VSS net6 VINP VINP net5 delay_cell
x8 VCC VSS net7 VINN VINN net6 delay_cell
x9 VCC VSS OUT START net7 nand
x10 VCC VSS START net9 net8 nand
.ends


* expanding   symbol:  /foss/designs/Comparator/schematic/Edge_pursuit_comparator/delay_cell.sym #
*+ of pins=6
** sym_path: /foss/designs/Comparator/schematic/Edge_pursuit_comparator/delay_cell.sym
** sch_path: /foss/designs/Comparator/schematic/Edge_pursuit_comparator/delay_cell.sch
.subckt delay_cell VCC VSS IN VINP VINN OUT
*.iopin VCC
*.opin OUT
*.ipin VINP
*.ipin VINN
*.iopin VSS
*.ipin IN
XM1 OUT IN net1 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM2 OUT IN net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM3 net2 VINN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM4 net1 VINP VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
.ends


* expanding   symbol:  /foss/designs/Comparator/schematic/Edge_pursuit_comparator/nand.sym # of
*+ pins=5
** sym_path: /foss/designs/Comparator/schematic/Edge_pursuit_comparator/nand.sym
** sch_path: /foss/designs/Comparator/schematic/Edge_pursuit_comparator/nand.sch
.subckt nand VCC VSS A B OUT
*.iopin VCC
*.opin OUT
*.ipin B
*.iopin VSS
*.ipin A
XM1 OUT B VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM2 OUT A net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM3 net1 B VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
XM4 OUT A VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1
.ends

.end
