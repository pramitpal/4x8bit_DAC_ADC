* SPICE3 file created from 4x8bit_tx_buffer.ext - technology: sky130A

.subckt x4x8bit_tx_buffer D00 D01 D02 D03 D04 D05 D06 D07 D10 D11 D12 D13 D14 D15
+ D16 D17 D20 D21 D22 D23 D24 D25 D26 D27 D30 D31 D32 D33 D34 D35 D36 D37 VCCD VDDA
+ VOUT0 VOUT1 VOUT2 VOUT3 VREFH VREFL VSSA VSSD
X0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X14 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X15 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X16 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X17 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X18 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X19 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X20 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X22 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X23 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X24 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X25 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X26 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X27 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X28 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X29 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X31 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X32 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X33 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=513 ps=4.48k w=1 l=0.5
X34 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X35 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X36 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=254 ps=2.65k w=0.5 l=0.5
X37 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X38 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X39 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X40 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X41 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X42 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X43 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X44 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X45 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X46 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X47 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X48 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X49 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X50 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X51 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X52 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X53 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X54 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X55 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X56 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X57 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X58 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X59 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X60 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X61 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X62 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X63 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X64 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X65 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X66 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X67 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X68 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X69 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X70 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X71 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X72 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X73 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X74 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X75 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X76 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X77 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X78 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X79 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X80 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X81 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X82 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X83 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X84 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X85 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X86 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X87 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X88 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X89 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X90 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X91 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X92 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X93 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X94 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X95 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X96 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X97 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X98 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X99 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X100 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X101 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X102 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X103 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X104 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X105 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X106 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X107 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X108 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X109 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X110 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X111 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X112 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X113 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X114 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X115 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X116 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X117 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X118 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X119 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X120 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X121 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X122 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X123 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X124 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X125 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X126 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X127 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X128 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X129 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X130 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X131 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X132 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X133 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X134 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X135 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X136 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X137 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X138 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X139 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X140 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X141 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X142 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X143 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X144 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X145 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X146 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X147 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X148 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X149 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X150 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X151 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X152 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X153 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X154 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X155 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X156 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X157 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X158 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X159 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X160 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X161 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X162 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X163 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X164 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X165 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X166 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X167 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X168 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X169 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X170 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X171 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X172 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X173 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X174 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X175 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X176 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X177 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X178 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X179 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X180 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X181 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X182 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X183 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X184 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X185 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X186 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X187 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X188 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X189 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X190 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X191 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X192 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X193 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X194 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X195 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X196 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X197 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X198 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X199 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X200 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X201 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X202 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X203 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X204 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X205 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X206 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X207 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X208 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X209 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X210 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X211 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X212 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X213 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X214 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X215 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X216 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X217 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X218 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X219 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X220 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X221 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X222 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X223 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X224 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X225 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X226 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X227 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X228 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X229 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X230 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X231 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X232 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X233 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X234 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X235 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X236 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X237 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X238 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X239 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X240 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X241 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X242 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X243 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X244 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X245 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X246 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X247 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X248 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X249 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X250 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X251 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X252 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X253 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X254 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X255 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X256 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X257 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X258 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X259 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X260 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X261 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X262 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X263 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X264 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X265 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X266 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X267 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X268 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X269 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X270 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X271 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X272 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X273 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X274 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X275 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X276 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X277 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X278 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X279 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X280 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X281 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X282 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X283 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X284 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X285 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X286 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X287 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X288 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X289 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X290 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X291 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X292 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X293 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X294 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X295 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X296 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X297 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X298 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X299 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X300 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X301 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X302 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X303 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X304 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X305 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X306 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X307 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X308 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X309 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X310 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X311 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X312 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X313 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X314 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X315 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X316 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X317 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X318 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X319 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X320 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X321 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X322 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X323 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X324 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X325 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X326 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X327 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X328 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X329 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X330 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X331 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X332 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X333 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X334 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X335 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X336 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X337 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X338 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X339 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X340 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X341 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X342 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X343 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X344 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X345 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X346 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X347 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X348 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X349 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X350 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X351 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X352 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X353 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X354 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X355 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X356 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X357 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X358 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X359 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X360 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X361 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X362 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X363 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X364 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X365 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X366 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X367 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X368 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X369 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X370 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X371 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X372 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X373 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X374 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X375 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X376 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X377 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X378 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X379 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X380 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X381 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X382 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X383 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X384 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X385 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X386 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X387 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X388 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X389 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X390 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X391 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X392 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X393 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X394 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X395 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X396 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X397 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X398 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X399 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X400 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X401 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X402 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X403 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X404 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X405 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X406 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X407 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X408 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X409 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X410 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X411 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X412 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X413 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X414 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X415 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X416 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X417 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X418 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X419 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X420 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X421 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X422 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X423 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X424 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X425 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X426 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X427 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X428 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X429 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X430 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X431 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X432 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X433 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X434 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X435 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X436 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X437 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X438 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X439 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X440 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X441 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X442 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X443 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X444 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X445 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X446 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X447 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X448 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X449 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X450 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X451 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X452 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X453 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X454 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X455 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X456 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X457 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X458 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X459 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X460 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X461 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X462 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X463 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X464 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X465 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X466 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X467 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X468 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X469 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X470 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X471 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X472 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X473 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X474 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X475 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X476 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X477 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X478 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X479 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X480 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X481 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X482 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X483 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X484 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X485 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X486 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X487 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X488 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X489 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X490 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X491 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X492 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X493 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X494 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X495 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X496 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X497 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X498 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X499 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X500 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X501 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X502 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X503 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X504 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X505 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X506 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X507 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X508 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X509 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X510 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X511 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X512 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X513 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X514 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X515 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X516 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X517 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X518 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X519 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X520 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X521 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X522 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X523 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X524 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X525 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X526 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X527 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X528 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X529 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X530 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X531 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X532 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X533 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X534 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X535 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X536 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X537 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X538 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X539 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X540 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X541 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X542 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X543 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X544 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X545 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X546 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X547 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X548 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X549 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X550 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X551 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X552 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X553 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X554 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X555 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X556 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X557 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X558 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X559 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X560 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X561 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X562 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X563 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X564 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X565 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X566 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X567 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X568 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X569 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X570 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X571 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X572 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X573 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X574 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X575 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X576 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X577 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X578 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X579 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X580 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X581 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X582 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X583 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X584 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X585 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X586 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X587 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X588 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X589 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X590 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X591 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X592 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X593 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X594 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X595 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X596 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X597 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X598 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X599 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X600 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X601 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X602 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X603 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X604 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X605 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X606 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X607 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X608 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X609 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X610 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X611 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X612 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X613 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X614 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X615 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X616 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X617 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X618 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X619 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X620 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X621 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X622 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X623 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X624 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X625 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X626 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X627 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X628 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X629 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X630 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X631 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X632 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X633 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X634 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X635 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X636 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X637 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X638 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X639 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X640 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X641 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X642 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X643 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X644 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X645 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X646 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X647 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X648 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X649 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X650 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X651 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X652 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X653 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X654 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X655 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X656 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X657 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X658 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X659 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X660 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X661 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X662 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X663 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X664 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X665 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X666 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X667 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X668 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X669 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X670 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X671 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X672 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X673 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X674 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X675 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X676 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X677 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X678 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X679 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X680 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X681 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X682 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X683 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X684 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X685 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X686 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X687 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X688 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X689 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X690 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X691 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X692 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X693 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X694 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X695 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X696 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X697 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X698 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X699 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X700 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X701 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X702 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X703 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X704 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X705 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X706 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X707 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X708 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X709 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X710 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X711 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X712 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X713 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X714 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X715 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X716 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X717 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X718 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X719 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X720 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X721 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X722 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X723 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X724 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X725 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X726 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X727 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X728 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X729 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X730 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X731 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X732 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X733 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X734 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X735 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X736 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X737 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X738 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X739 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X740 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X741 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X742 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X743 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X744 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X745 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X746 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X747 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X748 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X749 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X750 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X751 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X752 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X753 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X754 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X755 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X756 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X757 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X758 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X759 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X760 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X761 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X762 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X763 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X764 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X765 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X766 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X767 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X768 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X769 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X770 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X771 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X772 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X773 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X774 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X775 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X776 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X777 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X778 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X779 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X780 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X781 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X782 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X783 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X784 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X785 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X786 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X787 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X788 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X789 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X790 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X791 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X792 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X793 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X794 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X795 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X796 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X797 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X798 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X799 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X800 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X801 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X802 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X803 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X804 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X805 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X806 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X807 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X808 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X809 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X810 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X811 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X812 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X813 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X814 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X815 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X816 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X817 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X818 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X819 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X820 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X821 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X822 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X823 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X824 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X825 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X826 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X827 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X828 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X829 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X830 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X831 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X832 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X833 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X834 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X835 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X836 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X837 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X838 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X839 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X840 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X841 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X842 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X843 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X844 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X845 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X846 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X847 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X848 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X849 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X850 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X851 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X852 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X853 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X854 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X855 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X856 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X857 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X858 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X859 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X860 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X861 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X862 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X863 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X864 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X865 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X866 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X867 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X868 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X869 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X870 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X871 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X872 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X873 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X874 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X875 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X876 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X877 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X878 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X879 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X880 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X881 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X882 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X883 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X884 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X885 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X886 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X887 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X888 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X889 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X890 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X891 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X892 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X893 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X894 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X895 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X896 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X897 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X898 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X899 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X900 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X901 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X902 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X903 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X904 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X905 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X906 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X907 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X908 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X909 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X910 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X911 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X912 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X913 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X914 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X915 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X916 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X917 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X918 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X919 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X920 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X921 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X922 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X923 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X924 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X925 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X926 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X927 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X928 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X929 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X930 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X931 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X932 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X933 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X934 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X935 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X936 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X937 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X938 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X939 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X940 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X941 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X942 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X943 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X944 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X945 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X946 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X947 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X948 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X949 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X950 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X951 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X952 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X953 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X954 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X955 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X956 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X957 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X958 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X959 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X960 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X961 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X962 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X963 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X964 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X965 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X966 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X967 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X968 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X969 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X970 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X971 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X972 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X973 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X974 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X975 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X976 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X977 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X978 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X979 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X980 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X981 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X982 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X983 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X984 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X985 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X986 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X987 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X988 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X989 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X990 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X991 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X992 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X993 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X994 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X995 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X996 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X997 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X998 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X999 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1000 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1001 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1002 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1003 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1004 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1005 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1006 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1007 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1008 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1009 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1010 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1011 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1012 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1013 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1014 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1015 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1016 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1017 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1018 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1019 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1020 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1021 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1022 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1023 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1024 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1025 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1026 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1027 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1028 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1029 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1030 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1031 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1032 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1033 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1034 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1035 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1036 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1037 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1038 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1039 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1040 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1041 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1042 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1043 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1044 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1045 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1046 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1047 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1048 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1049 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1050 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1051 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1052 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1053 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1054 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1055 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1056 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1057 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1058 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1059 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1060 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1061 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1062 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1063 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1064 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1065 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1066 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1067 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1068 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1069 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1070 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1071 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1072 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1073 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1074 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1075 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1076 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1077 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1078 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1079 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1080 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1081 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1082 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1083 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1084 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1085 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1086 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1087 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1088 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1089 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1090 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1091 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1092 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1093 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1094 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1095 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1096 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1097 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1098 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1099 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1100 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1101 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1102 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1103 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1104 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1105 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1106 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1107 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1108 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1109 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1110 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1111 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1112 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1113 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1114 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1115 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1116 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1117 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1118 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1119 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1120 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1121 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1122 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1123 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1124 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1125 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1126 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1127 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1128 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1129 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1130 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1131 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1132 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1133 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1134 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1135 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1136 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1137 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1138 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1139 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1140 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1141 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1142 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1143 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1144 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1145 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1146 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1147 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1148 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1149 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1150 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1151 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1152 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1153 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1154 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1155 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1156 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1157 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1158 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1159 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1160 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1161 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1162 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1163 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1164 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1165 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1166 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1167 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1168 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1169 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1170 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1171 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1172 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1173 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1174 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1175 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1176 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1177 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1178 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1179 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1180 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1181 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1182 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1183 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1184 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1185 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1186 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1187 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1188 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1189 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1190 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1191 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1192 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1193 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1194 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1195 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1196 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1197 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1198 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1199 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1200 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1201 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1202 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1203 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1204 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1205 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1206 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1207 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1208 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1209 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1210 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1211 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1212 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1213 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1214 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1215 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1216 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1217 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1218 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1219 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1220 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1221 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1222 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1223 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1224 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1225 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1226 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1227 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1228 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1229 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1230 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1231 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1232 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1233 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1234 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1235 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1236 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1237 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1238 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1239 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1240 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1241 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1242 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1243 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1244 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1245 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1246 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1247 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1248 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1249 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1250 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1251 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1252 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1253 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1254 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1255 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1256 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1257 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1258 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1259 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1260 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1261 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1262 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1263 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1264 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1265 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1266 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1267 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1268 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1269 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1270 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1271 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1272 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1273 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1274 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1275 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1276 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1277 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1278 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1279 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1280 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1281 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1282 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1283 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1284 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1285 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1286 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1287 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1288 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1289 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1290 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1291 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1292 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1293 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1294 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1295 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1296 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1297 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1298 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1299 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1300 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1301 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1302 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1303 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1304 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1305 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1306 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1307 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1308 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1309 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1310 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1311 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1312 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1313 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1314 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1315 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1316 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1317 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1318 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1319 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1320 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1321 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1322 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1323 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1324 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1325 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1326 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1327 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1328 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1329 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1330 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1331 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1332 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1333 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1334 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1335 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1336 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1337 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1338 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1339 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1340 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1341 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1342 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1343 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1344 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1345 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1346 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1347 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1348 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1349 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1350 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1351 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1352 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1353 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1354 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1355 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1356 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1357 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1358 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1359 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1360 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1361 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1362 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1363 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1364 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1365 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1366 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1367 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1368 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1369 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1370 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1371 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1372 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1373 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1374 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1375 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1376 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1377 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1378 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1379 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1380 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1381 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1382 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1383 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1384 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1385 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1386 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1387 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1388 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1389 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1390 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1391 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1392 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1393 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1394 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1395 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1396 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1397 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1398 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1399 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1400 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1401 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1402 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1403 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1404 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1405 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1406 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1407 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1408 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1409 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1410 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1411 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1412 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1413 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1414 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1415 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1416 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1417 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1418 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1419 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1420 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1421 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1422 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1423 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1424 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1425 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1426 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1427 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1428 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1429 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1430 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1431 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1432 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1433 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1434 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1435 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1436 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1437 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1438 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1439 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1440 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1441 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1442 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1443 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1444 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1445 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1446 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1447 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1448 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1449 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1450 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1451 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1452 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1453 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1454 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1455 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1456 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1457 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1458 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1459 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1460 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1461 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1462 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1463 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1464 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1465 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1466 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1467 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1468 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1469 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1470 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1471 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1472 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1473 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1474 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1475 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1476 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1477 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1478 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1479 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1480 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1481 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1482 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1483 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1484 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1485 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1486 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1487 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1488 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1489 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1490 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1491 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1492 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1493 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1494 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1495 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1496 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1497 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1498 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1499 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1500 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1501 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1502 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1503 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1504 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1505 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1506 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1507 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1508 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1509 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1510 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1511 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1512 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1513 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1514 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1515 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1516 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1517 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1518 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1519 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1520 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1521 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1522 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1523 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1524 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1525 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1526 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1527 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1528 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1529 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1530 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1531 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1532 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1533 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1534 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1535 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1536 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1537 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1538 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1539 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1540 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1541 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1542 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1543 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1544 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1545 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1546 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1547 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1548 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1549 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1550 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1551 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1552 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1553 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1554 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1555 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1556 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1557 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1558 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1559 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1560 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1561 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1562 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1563 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1564 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1565 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1566 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1567 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1568 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1569 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1570 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1571 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1572 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1573 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1574 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1575 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1576 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1577 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1578 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1579 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1580 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1581 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1582 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1583 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1584 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1585 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1586 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1587 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1588 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1589 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1590 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1591 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1592 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1593 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1594 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1595 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1596 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1597 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1598 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1599 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1600 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1601 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1602 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1603 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1604 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1605 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1606 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1607 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1608 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1609 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1610 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1611 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1612 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1613 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1614 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1615 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1616 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1617 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1618 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1619 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1620 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1621 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1622 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1623 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1624 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1625 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1626 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1627 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1628 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1629 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1630 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1631 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1632 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1633 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1634 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1635 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1636 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1637 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1638 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1639 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1640 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1641 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1642 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1643 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1644 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1645 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1646 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1647 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1648 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1649 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1650 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1651 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1652 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1653 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1654 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1655 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1656 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1657 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1658 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1659 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1660 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1661 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1662 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1663 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1664 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1665 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1666 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1667 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1668 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1669 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1670 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1671 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1672 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1673 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1674 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1675 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1676 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1677 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1678 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1679 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1680 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1681 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1682 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1683 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1684 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1685 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1686 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1687 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1688 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1689 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1690 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1691 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1692 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1693 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1694 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1695 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1696 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1697 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1698 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1699 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1700 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1701 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1702 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1703 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1704 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1705 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1706 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1707 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1708 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1709 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1710 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1711 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1712 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1713 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1714 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1715 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1716 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1717 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1718 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1719 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1720 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1721 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1722 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1723 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1724 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1725 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1726 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1727 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1728 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1729 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1730 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1731 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1732 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1733 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1734 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1735 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1736 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1737 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1738 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1739 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1740 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1741 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1742 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1743 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1744 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1745 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1746 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1747 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1748 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1749 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1750 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1751 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1752 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1753 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1754 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1755 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1756 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1757 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1758 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1759 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1760 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1761 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1762 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1763 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1764 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1765 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1766 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1767 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1768 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1769 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1770 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1771 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1772 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1773 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1774 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1775 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1776 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1777 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1778 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1779 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1780 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1781 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1782 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1783 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1784 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1785 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1786 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1787 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1788 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1789 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1790 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1791 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1792 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1793 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1794 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1795 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1796 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1797 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1798 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1799 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1800 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1801 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1802 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1803 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1804 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1805 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1806 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1807 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1808 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1809 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1810 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1811 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1812 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1813 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1814 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1815 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1816 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1817 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1818 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1819 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1820 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1821 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1822 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1823 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1824 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1825 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1826 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1827 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1828 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1829 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1830 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1831 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1832 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1833 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1834 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1835 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1836 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1837 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1838 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1839 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1840 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1841 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1842 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1843 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1844 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1845 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1846 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1847 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1848 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1849 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1850 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1851 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1852 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1853 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1854 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1855 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1856 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1857 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1858 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1859 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1860 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1861 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1862 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1863 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1864 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1865 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1866 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1867 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1868 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1869 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1870 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1871 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1872 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1873 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1874 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1875 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1876 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1877 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1878 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1879 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1880 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1881 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1882 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1883 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1884 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1885 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1886 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1887 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1888 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1889 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1890 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1891 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1892 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1893 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1894 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1895 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1896 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1897 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1898 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1899 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1900 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1901 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1902 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1903 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1904 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1905 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1906 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1907 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1908 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1909 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1910 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1911 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1912 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1913 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1914 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1915 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1916 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1917 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1918 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1919 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1920 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1921 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1922 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1923 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1924 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1925 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1926 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1927 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1928 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1929 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1930 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1931 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1932 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1933 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1934 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1935 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1936 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1937 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1938 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1939 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1940 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1941 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1942 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1943 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1944 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1945 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1946 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1947 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1948 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1949 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1950 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1951 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1952 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1953 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1954 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1955 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1956 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1957 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1958 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1959 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1960 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1961 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1962 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1963 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1964 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1965 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1966 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1967 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1968 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1969 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1970 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1971 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1972 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1973 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1974 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1975 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1976 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1977 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1978 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1979 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1980 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1981 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1982 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1983 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1984 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1985 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1986 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1987 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1988 VREFL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=10.3 as=0 ps=0 w=1 l=0.5
X1989 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1990 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1991 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VREFL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.45 ps=13.8 w=0.5 l=0.5
X1992 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1993 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1994 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1995 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VREFL VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1996 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1997 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1998 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1999 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2000 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2001 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2002 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2003 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2004 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2005 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2006 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2007 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2008 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2009 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2010 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2011 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2012 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2013 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2014 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2015 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2016 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2017 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2018 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2019 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2020 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2021 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2022 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2023 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2024 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2025 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2026 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2027 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2028 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2029 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2030 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2031 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2032 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X2033 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2034 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2035 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X2036 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2037 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2038 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2039 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2040 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X2041 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2042 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2043 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2044 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2045 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D00 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X2046 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2047 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D00 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X2048 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=37.1 pd=275 as=1.16 ps=8.58 w=4 l=0.5
X2049 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X2050 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=15.6 ps=145 w=0.84 l=0.15
X2051 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2052 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2053 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D01 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2054 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=7.8 ps=90.9 w=0.42 l=0.15
X2055 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D01 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2056 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X2057 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X2058 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2059 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2060 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2061 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D02 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2062 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2063 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D02 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2064 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X2065 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X2066 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2067 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2068 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2069 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D03 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2070 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2071 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D03 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2072 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X2073 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X2074 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2075 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2076 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2077 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D04 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2078 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2079 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D04 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2080 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X2081 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X2082 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2083 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2084 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2085 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D05 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2086 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2087 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D05 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2088 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X2089 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X2090 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2091 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2092 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2093 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D06 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2094 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2095 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D06 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2096 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X2097 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X2098 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2099 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2100 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2101 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D07 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X2102 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2103 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D07 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X2104 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1549_3140# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2105 VOUT0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.5
X2106 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VOUT0 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=0.87 ps=6.29 w=6 l=0.5
X2107 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2108 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1095_1321# VOUT0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_937_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X2109 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VOUT0 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.5
X2110 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2111 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
R0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VSSA sky130_fd_pr__res_generic_po w=0.33 l=65.2
X2112 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2113 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1549_3140# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2114 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VOUT0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X2115 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1549_3140# VOUT0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1392_2207# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X2116 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1095_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2117 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1095_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X2118 VOUT0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.6 w=6 l=0.5
X2119 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2120 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X2121 VOUT0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X2122 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
R1 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# sky130_fd_pr__res_generic_po w=0.33 l=38.5
X2123 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X2124 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X2125 VOUT0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=0.5
X2126 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VOUT0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=0.5
X2127 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2128 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X2129 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2130 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
R2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# VSSA sky130_fd_pr__res_generic_po w=0.33 l=23.6
X2131 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2132 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2133 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2134 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2135 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2136 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2137 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2138 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2139 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2140 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2141 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2142 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2143 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2144 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2145 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2146 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2147 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2148 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2149 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2150 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2151 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2152 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2153 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2154 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2155 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2156 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2157 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2158 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2159 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2160 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2161 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2162 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2163 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2164 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2165 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2166 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2167 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2168 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2169 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2170 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2171 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2172 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2173 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2174 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2175 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2176 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2177 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2178 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2179 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2180 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2181 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2182 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2183 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2184 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2185 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2186 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2187 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2188 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2189 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2190 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2191 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2192 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2193 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2194 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2195 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2196 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2197 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2198 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2199 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2200 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2201 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2202 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2203 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2204 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2205 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2206 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2207 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2208 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2209 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2210 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2211 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2212 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2213 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2214 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2215 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2216 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2217 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2218 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2219 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2220 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2221 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2222 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2223 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2224 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2225 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2226 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2227 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2228 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2229 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2230 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2231 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2232 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2233 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2234 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2235 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2236 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2237 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2238 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2239 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2240 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2241 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2242 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2243 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2244 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2245 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2246 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2247 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2248 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2249 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2250 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2251 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2252 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2253 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2254 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2255 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2256 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2257 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2258 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2259 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2260 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2261 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2262 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2263 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2264 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2265 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2266 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2267 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2268 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2269 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2270 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2271 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2272 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2273 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2274 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2275 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2276 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2277 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2278 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2279 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2280 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2281 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2282 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2283 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2284 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2285 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2286 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2287 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2288 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2289 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2290 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2291 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2292 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2293 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2294 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2295 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2296 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2297 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2298 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2299 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2300 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2301 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2302 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2303 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2304 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2305 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2306 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2307 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2308 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2309 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2310 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2311 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2312 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2313 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2314 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2315 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2316 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2317 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2318 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2319 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2320 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2321 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2322 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2323 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2324 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2325 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2326 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2327 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2328 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2329 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2330 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2331 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2332 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2333 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2334 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2335 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2336 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2337 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2338 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2339 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2340 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2341 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2342 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2343 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2344 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2345 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2346 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2347 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2348 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2349 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2350 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2351 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2352 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2353 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2354 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2355 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2356 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2357 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2358 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2359 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2360 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2361 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2362 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2363 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2364 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2365 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2366 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2367 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2368 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2369 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2370 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2371 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2372 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2373 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2374 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2375 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2376 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2377 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2378 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2379 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2380 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2381 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2382 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2383 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2384 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2385 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2386 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2387 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2388 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2389 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2390 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2391 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2392 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2393 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2394 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2395 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2396 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2397 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2398 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2399 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2400 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2401 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2402 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2403 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2404 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2405 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2406 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2407 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2408 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2409 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2410 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2411 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2412 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2413 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2414 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2415 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2416 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2417 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2418 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2419 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2420 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2421 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2422 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2423 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2424 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2425 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2426 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2427 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2428 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2429 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2430 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2431 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2432 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2433 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2434 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2435 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2436 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2437 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2438 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2439 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2440 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2441 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2442 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2443 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2444 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2445 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2446 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2447 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2448 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2449 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2450 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2451 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2452 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2453 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2454 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2455 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2456 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2457 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2458 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2459 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2460 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2461 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2462 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2463 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2464 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2465 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2466 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2467 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2468 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2469 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2470 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2471 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2472 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2473 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2474 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2475 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2476 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2477 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2478 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2479 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2480 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2481 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2482 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2483 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2484 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2485 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2486 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2487 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2488 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2489 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2490 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2491 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2492 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2493 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2494 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2495 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2496 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2497 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2498 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2499 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2500 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2501 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2502 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2503 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2504 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2505 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2506 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2507 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2508 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2509 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2510 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2511 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2512 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2513 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2514 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2515 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2516 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2517 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2518 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2519 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2520 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2521 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2522 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2523 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2524 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2525 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2526 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2527 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2528 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2529 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2530 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2531 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2532 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2533 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2534 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2535 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2536 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2537 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2538 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2539 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2540 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2541 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2542 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2543 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2544 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2545 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2546 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2547 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2548 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2549 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2550 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2551 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2552 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2553 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2554 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2555 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2556 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2557 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2558 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2559 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2560 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2561 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2562 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2563 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2564 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2565 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2566 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2567 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2568 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2569 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2570 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2571 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2572 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2573 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2574 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2575 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2576 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2577 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2578 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2579 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2580 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2581 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2582 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2583 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2584 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2585 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2586 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2587 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2588 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2589 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2590 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2591 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2592 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2593 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2594 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2595 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2596 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2597 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2598 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2599 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2600 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2601 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2602 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2603 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2604 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2605 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2606 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2607 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2608 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2609 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2610 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2611 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2612 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2613 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2614 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2615 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2616 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2617 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2618 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2619 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2620 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2621 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2622 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2623 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2624 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2625 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2626 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2627 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2628 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2629 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2630 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2631 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2632 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2633 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2634 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2635 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2636 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2637 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2638 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2639 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2640 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2641 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2642 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2643 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2644 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2645 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2646 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2647 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2648 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2649 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2650 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2651 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2652 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2653 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2654 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2655 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2656 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2657 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2658 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2659 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2660 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2661 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2662 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2663 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2664 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2665 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2666 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2667 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2668 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2669 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2670 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2671 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2672 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2673 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2674 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2675 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2676 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2677 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2678 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2679 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2680 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2681 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2682 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2683 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2684 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2685 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2686 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2687 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2688 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2689 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2690 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2691 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2692 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2693 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2694 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2695 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2696 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2697 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2698 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2699 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2700 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2701 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2702 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2703 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2704 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2705 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2706 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2707 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2708 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2709 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2710 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2711 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2712 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2713 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2714 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2715 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2716 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2717 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2718 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2719 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2720 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2721 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2722 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2723 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2724 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2725 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2726 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2727 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2728 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2729 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2730 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2731 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2732 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2733 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2734 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2735 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2736 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2737 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2738 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2739 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2740 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2741 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2742 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2743 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2744 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2745 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2746 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2747 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2748 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2749 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2750 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2751 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2752 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2753 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2754 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2755 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2756 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2757 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2758 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2759 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2760 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2761 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2762 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2763 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2764 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2765 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2766 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2767 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2768 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2769 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2770 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2771 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2772 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2773 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2774 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2775 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2776 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2777 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2778 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2779 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2780 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2781 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2782 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2783 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2784 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2785 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2786 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2787 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2788 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2789 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2790 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2791 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2792 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2793 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2794 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2795 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2796 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2797 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2798 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2799 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2800 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2801 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2802 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2803 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2804 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2805 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2806 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2807 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2808 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2809 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2810 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2811 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2812 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2813 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2814 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2815 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2816 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2817 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2818 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2819 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2820 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2821 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2822 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2823 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2824 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2825 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2826 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2827 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2828 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2829 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2830 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2831 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2832 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2833 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2834 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2835 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2836 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2837 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2838 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2839 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2840 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2841 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2842 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2843 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2844 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2845 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2846 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2847 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2848 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2849 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2850 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2851 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2852 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2853 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2854 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2855 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2856 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2857 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2858 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2859 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2860 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2861 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2862 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2863 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2864 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2865 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2866 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2867 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2868 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2869 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2870 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2871 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2872 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2873 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2874 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2875 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2876 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2877 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2878 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2879 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2880 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2881 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2882 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2883 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2884 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2885 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2886 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2887 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2888 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2889 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2890 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2891 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2892 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2893 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2894 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2895 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2896 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2897 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2898 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2899 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2900 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2901 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2902 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2903 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2904 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2905 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2906 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2907 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2908 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2909 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2910 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2911 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2912 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2913 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2914 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2915 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2916 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2917 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2918 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2919 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2920 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2921 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2922 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2923 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2924 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2925 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2926 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2927 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2928 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2929 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2930 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2931 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2932 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2933 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2934 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2935 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2936 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2937 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2938 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2939 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2940 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2941 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2942 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2943 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2944 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2945 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2946 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2947 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2948 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2949 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2950 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2951 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2952 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2953 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2954 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2955 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2956 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2957 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2958 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2959 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2960 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2961 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2962 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2963 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2964 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2965 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2966 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2967 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2968 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2969 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2970 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2971 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2972 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2973 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2974 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2975 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2976 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2977 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2978 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2979 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2980 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2981 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2982 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2983 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2984 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2985 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2986 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2987 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2988 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2989 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2990 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2991 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2992 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2993 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2994 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2995 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2996 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2997 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2998 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2999 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3000 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3001 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3002 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3003 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3004 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3005 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3006 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3007 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3008 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3009 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3010 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3011 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3012 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3013 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3014 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3015 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3016 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3017 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3018 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3019 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3020 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3021 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3022 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3023 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3024 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3025 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3026 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3027 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3028 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3029 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3030 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3031 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3032 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3033 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3034 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3035 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3036 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3037 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3038 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3039 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3040 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3041 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3042 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3043 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3044 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3045 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3046 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3047 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3048 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3049 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3050 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3051 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3052 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3053 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3054 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3055 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3056 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3057 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3058 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3059 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3060 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3061 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3062 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3063 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3064 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3065 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3066 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3067 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3068 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3069 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3070 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3071 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3072 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3073 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3074 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3075 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3076 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3077 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3078 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3079 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3080 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3081 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3082 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3083 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3084 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3085 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3086 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3087 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3088 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3089 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3090 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3091 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3092 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3093 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3094 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3095 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3096 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3097 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3098 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3099 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3100 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3101 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3102 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3103 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3104 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3105 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3106 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3107 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3108 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3109 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3110 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3111 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3112 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3113 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3114 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3115 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3116 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3117 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3118 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3119 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3120 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3121 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3122 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3123 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3124 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3125 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3126 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3127 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3128 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3129 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3130 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3131 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3132 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3133 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3134 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3135 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3136 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3137 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3138 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3139 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3140 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3141 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3142 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3143 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3144 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3145 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3146 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3147 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3148 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3149 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3150 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3151 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3152 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3153 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3154 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3155 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3156 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3157 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3158 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3159 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3160 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3161 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3162 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3163 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3164 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3165 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3166 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3167 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3168 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3169 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3170 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3171 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3172 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3173 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3174 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3175 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3176 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3177 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3178 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3179 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3180 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3181 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3182 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3183 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3184 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3185 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3186 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3187 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3188 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3189 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3190 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3191 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3192 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3193 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3194 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3195 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3196 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3197 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3198 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3199 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3200 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3201 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3202 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3203 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3204 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3205 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3206 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3207 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3208 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3209 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3210 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3211 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3212 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3213 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3214 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3215 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3216 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3217 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3218 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3219 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3220 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3221 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3222 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3223 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3224 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3225 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3226 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3227 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3228 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3229 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3230 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3231 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3232 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3233 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3234 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3235 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3236 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3237 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3238 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3239 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3240 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3241 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3242 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3243 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3244 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3245 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3246 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3247 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3248 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3249 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3250 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3251 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3252 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3253 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3254 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3255 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3256 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3257 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3258 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3259 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3260 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3261 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3262 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3263 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3264 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3265 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3266 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3267 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3268 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3269 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3270 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3271 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3272 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3273 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3274 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3275 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3276 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3277 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3278 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3279 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3280 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3281 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3282 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3283 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3284 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3285 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3286 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3287 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3288 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3289 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3290 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3291 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3292 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3293 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3294 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3295 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3296 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3297 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3298 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3299 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3300 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3301 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3302 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3303 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3304 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3305 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3306 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3307 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3308 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3309 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3310 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3311 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3312 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3313 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3314 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3315 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3316 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3317 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3318 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3319 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3320 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3321 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3322 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3323 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3324 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3325 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3326 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3327 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3328 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3329 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3330 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3331 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3332 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3333 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3334 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3335 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3336 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3337 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3338 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3339 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3340 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3341 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3342 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3343 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3344 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3345 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3346 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3347 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3348 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3349 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3350 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3351 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3352 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3353 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3354 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3355 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3356 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3357 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3358 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3359 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3360 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3361 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3362 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3363 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3364 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3365 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3366 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3367 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3368 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3369 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3370 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3371 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3372 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3373 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3374 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3375 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3376 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3377 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3378 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3379 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3380 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3381 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3382 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3383 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3384 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3385 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3386 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3387 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3388 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3389 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3390 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3391 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3392 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3393 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3394 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3395 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3396 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3397 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3398 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3399 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3400 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3401 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3402 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3403 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3404 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3405 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3406 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3407 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3408 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3409 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3410 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3411 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3412 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3413 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3414 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3415 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3416 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3417 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3418 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3419 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3420 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3421 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3422 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3423 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3424 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3425 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3426 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3427 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3428 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3429 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3430 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3431 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3432 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3433 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3434 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3435 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3436 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3437 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3438 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3439 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3440 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3441 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3442 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3443 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3444 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3445 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3446 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3447 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3448 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3449 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3450 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3451 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3452 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3453 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3454 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3455 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3456 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3457 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3458 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3459 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3460 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3461 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3462 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3463 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3464 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3465 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3466 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3467 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3468 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3469 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3470 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3471 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3472 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3473 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3474 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3475 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3476 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3477 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3478 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3479 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3480 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3481 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3482 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3483 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3484 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3485 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3486 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3487 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3488 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3489 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3490 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3491 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3492 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3493 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3494 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3495 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3496 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3497 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3498 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3499 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3500 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3501 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3502 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3503 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3504 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3505 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3506 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3507 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3508 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3509 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3510 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3511 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3512 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3513 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3514 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3515 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3516 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3517 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3518 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3519 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3520 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3521 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3522 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3523 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3524 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3525 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3526 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3527 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3528 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3529 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3530 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3531 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3532 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3533 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3534 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3535 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3536 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3537 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3538 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3539 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3540 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3541 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3542 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3543 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3544 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3545 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3546 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3547 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3548 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3549 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3550 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3551 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3552 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3553 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3554 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3555 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3556 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3557 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3558 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3559 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3560 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3561 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3562 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3563 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3564 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3565 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3566 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3567 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3568 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3569 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3570 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3571 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3572 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3573 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3574 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3575 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3576 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3577 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3578 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3579 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3580 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3581 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3582 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3583 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3584 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3585 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3586 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3587 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3588 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3589 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3590 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3591 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3592 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3593 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3594 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3595 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3596 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3597 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3598 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3599 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3600 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3601 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3602 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3603 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3604 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3605 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3606 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3607 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3608 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3609 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3610 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3611 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3612 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3613 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3614 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3615 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3616 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3617 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3618 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3619 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3620 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3621 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3622 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3623 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3624 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3625 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3626 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3627 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3628 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3629 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3630 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3631 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3632 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3633 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3634 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3635 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3636 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3637 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3638 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3639 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3640 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3641 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3642 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3643 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3644 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3645 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3646 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3647 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3648 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3649 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3650 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3651 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3652 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3653 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3654 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3655 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3656 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3657 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3658 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3659 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3660 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3661 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3662 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3663 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3664 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3665 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3666 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3667 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3668 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3669 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3670 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3671 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3672 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3673 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3674 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3675 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3676 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3677 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3678 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3679 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3680 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3681 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3682 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3683 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3684 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3685 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3686 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3687 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3688 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3689 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3690 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3691 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3692 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3693 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3694 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3695 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3696 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3697 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3698 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3699 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3700 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3701 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3702 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3703 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3704 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3705 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3706 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3707 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3708 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3709 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3710 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3711 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3712 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3713 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3714 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3715 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3716 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3717 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3718 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3719 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3720 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3721 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3722 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3723 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3724 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3725 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3726 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3727 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3728 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3729 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3730 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3731 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3732 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3733 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3734 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3735 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3736 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3737 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3738 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3739 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3740 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3741 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3742 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3743 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3744 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3745 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3746 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3747 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3748 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3749 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3750 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3751 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3752 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3753 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3754 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3755 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3756 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3757 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3758 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3759 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3760 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3761 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3762 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3763 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3764 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3765 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3766 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3767 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3768 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3769 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3770 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3771 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3772 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3773 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3774 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3775 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3776 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3777 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3778 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3779 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3780 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3781 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3782 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3783 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3784 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3785 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3786 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3787 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3788 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3789 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3790 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3791 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3792 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3793 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3794 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3795 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3796 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3797 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3798 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3799 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3800 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3801 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3802 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3803 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3804 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3805 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3806 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3807 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3808 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3809 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3810 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3811 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3812 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3813 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3814 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3815 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3816 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3817 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3818 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3819 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3820 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3821 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3822 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3823 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3824 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3825 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3826 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3827 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3828 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3829 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3830 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3831 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3832 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3833 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3834 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3835 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3836 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3837 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3838 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3839 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3840 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3841 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3842 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3843 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3844 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3845 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3846 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3847 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3848 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3849 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3850 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3851 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3852 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3853 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3854 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3855 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3856 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3857 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3858 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3859 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3860 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3861 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3862 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3863 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3864 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3865 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3866 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3867 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3868 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3869 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3870 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3871 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3872 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3873 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3874 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3875 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3876 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3877 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3878 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3879 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3880 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3881 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3882 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3883 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3884 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3885 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3886 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3887 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3888 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3889 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3890 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3891 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3892 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3893 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3894 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3895 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3896 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3897 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3898 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3899 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3900 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3901 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3902 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3903 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3904 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3905 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3906 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3907 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3908 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3909 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3910 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3911 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3912 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3913 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3914 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3915 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3916 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3917 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3918 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3919 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3920 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3921 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3922 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3923 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3924 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3925 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3926 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3927 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3928 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3929 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3930 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3931 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3932 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3933 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3934 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3935 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3936 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3937 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3938 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3939 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3940 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3941 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3942 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3943 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3944 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3945 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3946 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3947 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3948 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3949 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3950 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3951 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3952 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3953 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3954 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3955 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3956 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3957 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3958 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3959 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3960 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3961 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3962 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3963 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3964 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3965 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3966 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3967 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3968 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3969 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3970 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3971 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3972 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3973 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3974 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3975 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3976 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3977 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3978 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3979 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3980 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3981 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3982 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3983 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3984 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3985 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3986 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3987 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3988 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3989 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3990 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3991 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3992 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3993 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3994 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3995 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3996 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3997 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3998 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3999 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4000 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4001 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4002 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4003 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4004 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4005 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4006 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4007 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4008 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4009 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4010 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4011 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4012 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4013 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4014 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4015 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4016 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4017 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4018 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4019 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4020 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4021 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4022 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4023 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4024 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4025 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4026 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4027 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4028 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4029 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4030 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4031 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4032 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4033 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4034 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4035 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4036 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4037 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4038 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4039 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4040 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4041 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4042 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4043 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4044 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4045 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4046 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4047 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4048 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4049 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4050 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4051 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4052 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4053 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4054 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4055 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4056 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4057 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4058 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4059 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4060 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4061 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4062 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4063 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4064 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4065 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4066 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4067 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4068 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4069 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4070 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4071 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4072 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4073 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4074 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4075 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4076 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4077 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4078 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4079 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4080 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4081 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4082 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4083 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4084 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4085 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4086 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4087 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4088 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4089 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4090 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4091 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4092 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4093 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4094 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4095 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4096 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4097 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4098 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4099 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4100 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4101 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4102 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4103 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4104 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4105 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4106 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4107 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4108 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4109 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4110 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4111 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4112 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4113 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4114 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4115 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4116 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4117 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4118 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4119 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4120 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4121 VREFL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4122 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4123 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4124 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VREFL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4125 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4126 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4127 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4128 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VREFL VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4129 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4130 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4131 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4132 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4133 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4134 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4135 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4136 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4137 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4138 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4139 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4140 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4141 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4142 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4143 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4144 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4145 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4146 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4147 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4148 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4149 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4150 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4151 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4152 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4153 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4154 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4155 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4156 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4157 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4158 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4159 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4160 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4161 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4162 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4163 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4164 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4165 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X4166 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4167 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4168 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X4169 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4170 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4171 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4172 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4173 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4174 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4175 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4176 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4177 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4178 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D10 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4179 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4180 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D10 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4181 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4182 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4183 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4184 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4185 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4186 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D11 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4187 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4188 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D11 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4189 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4190 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4191 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4192 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4193 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4194 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D12 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4195 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4196 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D12 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4197 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4198 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4199 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4200 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4201 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4202 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D13 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4203 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4204 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D13 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4205 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4206 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4207 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4208 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4209 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4210 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D14 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4211 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4212 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D14 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4213 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4214 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4215 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4216 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4217 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4218 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D15 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4219 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4220 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D15 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4221 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4222 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4223 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4224 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4225 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4226 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D16 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4227 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4228 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D16 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4229 VSSD 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4230 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4231 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4232 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4233 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4234 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D17 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X4235 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4236 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D17 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X4237 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1549_3140# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0 ps=0 w=2 l=0.5
X4238 VOUT1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=3.48 pd=25.2 as=0 ps=0 w=6 l=0.5
X4239 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VOUT1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X4240 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X4241 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1095_1321# VOUT1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_937_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=13.2 as=0.58 ps=4.58 w=2 l=0.5
X4242 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VOUT1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X4243 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4244 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=9.16 w=2 l=0.5
R3 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VSSA sky130_fd_pr__res_generic_po w=0.33 l=65.2
X4245 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0.58 ps=4.58 w=2 l=0.5
X4246 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1549_3140# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4247 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VOUT1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=5.8 ps=41.2 w=10 l=0.5
X4248 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1549_3140# VOUT1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1392_2207# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4249 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1095_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X4250 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1095_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
X4251 VOUT1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X4252 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=1.74 ps=13.2 w=2 l=0.5
X4253 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4254 VOUT1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X4255 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
R4 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# sky130_fd_pr__res_generic_po w=0.33 l=38.5
X4256 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
X4257 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4258 VOUT1 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X4259 VDDA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VOUT1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X4260 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=9.16 as=0 ps=0 w=2 l=0.5
X4261 VSSA 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X4262 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X4263 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
R5 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# VSSA sky130_fd_pr__res_generic_po w=0.33 l=23.6
X4264 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X4265 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# 2x8bit_tx_buffer_0[0]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X4266 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4267 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4268 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4269 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4270 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4271 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4272 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4273 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4274 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4275 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4276 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4277 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4278 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4279 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4280 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4281 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4282 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4283 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4284 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4285 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4286 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4287 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4288 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4289 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4290 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4291 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4292 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4293 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4294 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4295 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4296 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4297 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4298 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4299 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4300 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4301 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4302 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4303 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4304 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4305 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4306 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4307 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4308 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4309 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4310 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4311 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4312 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4313 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4314 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4315 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4316 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4317 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4318 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4319 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4320 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4321 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4322 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4323 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4324 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4325 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4326 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4327 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4328 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4329 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4330 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4331 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4332 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4333 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4334 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4335 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4336 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4337 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4338 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4339 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4340 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4341 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4342 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4343 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4344 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4345 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4346 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4347 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4348 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4349 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4350 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4351 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4352 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4353 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4354 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4355 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4356 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4357 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4358 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4359 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4360 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4361 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4362 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4363 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4364 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4365 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4366 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4367 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4368 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4369 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4370 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4371 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4372 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4373 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4374 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4375 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4376 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4377 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4378 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4379 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4380 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4381 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4382 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4383 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4384 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4385 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4386 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4387 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4388 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4389 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4390 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4391 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4392 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4393 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4394 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4395 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4396 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4397 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4398 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4399 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4400 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4401 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4402 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4403 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4404 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4405 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4406 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4407 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4408 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4409 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4410 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4411 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4412 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4413 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4414 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4415 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4416 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4417 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4418 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4419 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4420 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4421 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4422 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4423 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4424 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4425 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4426 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4427 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4428 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4429 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4430 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4431 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4432 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4433 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4434 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4435 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4436 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4437 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4438 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4439 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4440 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4441 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4442 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4443 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4444 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4445 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4446 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4447 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4448 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4449 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4450 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4451 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4452 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4453 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4454 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4455 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4456 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4457 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4458 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4459 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4460 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4461 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4462 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4463 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4464 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4465 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4466 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4467 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4468 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4469 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4470 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4471 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4472 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4473 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4474 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4475 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4476 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4477 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4478 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4479 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4480 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4481 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4482 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4483 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4484 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4485 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4486 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4487 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4488 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4489 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4490 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4491 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4492 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4493 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4494 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4495 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4496 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4497 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4498 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4499 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4500 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4501 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4502 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4503 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4504 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4505 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4506 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4507 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4508 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4509 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4510 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4511 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4512 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4513 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4514 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4515 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4516 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4517 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4518 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4519 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4520 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4521 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4522 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4523 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4524 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4525 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4526 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4527 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4528 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4529 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4530 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4531 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4532 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4533 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4534 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4535 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4536 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4537 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4538 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4539 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4540 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4541 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4542 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4543 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4544 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4545 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4546 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4547 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4548 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4549 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4550 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4551 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4552 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4553 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4554 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4555 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4556 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4557 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4558 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4559 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4560 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4561 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4562 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4563 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4564 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4565 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4566 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4567 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4568 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4569 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4570 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4571 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4572 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4573 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4574 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4575 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4576 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4577 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4578 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4579 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4580 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4581 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4582 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4583 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4584 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4585 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4586 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4587 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4588 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4589 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4590 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4591 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4592 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4593 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4594 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4595 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4596 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4597 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4598 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4599 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4600 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4601 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4602 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4603 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4604 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4605 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4606 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4607 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4608 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4609 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4610 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4611 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4612 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4613 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4614 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4615 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4616 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4617 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4618 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4619 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4620 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4621 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4622 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4623 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4624 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4625 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4626 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4627 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4628 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4629 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4630 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4631 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4632 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4633 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4634 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4635 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4636 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4637 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4638 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4639 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4640 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4641 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4642 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4643 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4644 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4645 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4646 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4647 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4648 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4649 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4650 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4651 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4652 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4653 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4654 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4655 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4656 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4657 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4658 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4659 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4660 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4661 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4662 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4663 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4664 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4665 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4666 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4667 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4668 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4669 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4670 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4671 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4672 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4673 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4674 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4675 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4676 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4677 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4678 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4679 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4680 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4681 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4682 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4683 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4684 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4685 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4686 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4687 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4688 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4689 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4690 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4691 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4692 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4693 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4694 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4695 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4696 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4697 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4698 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4699 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4700 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4701 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4702 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4703 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4704 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4705 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4706 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4707 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4708 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4709 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4710 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4711 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4712 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4713 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4714 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4715 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4716 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4717 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4718 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4719 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4720 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4721 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4722 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4723 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4724 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4725 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4726 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4727 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4728 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4729 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4730 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4731 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4732 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4733 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4734 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4735 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4736 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4737 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4738 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4739 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4740 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4741 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4742 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4743 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4744 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4745 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4746 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4747 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4748 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4749 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4750 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4751 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4752 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4753 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4754 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4755 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4756 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4757 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4758 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4759 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4760 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4761 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4762 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4763 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4764 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4765 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4766 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4767 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4768 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4769 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4770 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4771 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4772 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4773 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4774 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4775 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4776 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4777 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4778 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4779 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4780 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4781 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4782 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4783 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4784 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4785 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4786 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4787 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4788 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4789 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4790 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4791 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4792 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4793 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4794 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4795 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4796 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4797 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4798 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4799 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4800 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4801 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4802 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4803 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4804 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4805 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4806 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4807 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4808 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4809 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4810 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4811 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4812 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4813 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4814 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4815 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4816 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4817 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4818 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4819 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4820 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4821 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4822 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4823 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4824 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4825 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4826 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4827 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4828 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4829 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4830 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4831 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4832 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4833 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4834 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4835 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4836 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4837 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4838 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4839 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4840 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4841 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4842 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4843 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4844 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4845 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4846 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4847 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4848 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4849 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4850 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4851 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4852 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4853 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4854 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4855 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4856 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4857 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4858 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4859 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4860 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4861 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4862 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4863 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4864 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4865 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4866 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4867 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4868 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4869 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4870 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4871 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4872 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4873 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4874 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4875 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4876 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4877 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4878 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4879 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4880 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4881 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4882 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4883 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4884 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4885 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4886 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4887 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4888 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4889 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4890 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4891 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4892 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4893 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4894 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4895 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4896 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4897 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4898 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4899 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4900 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4901 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4902 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4903 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4904 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4905 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4906 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4907 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4908 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4909 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4910 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4911 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4912 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4913 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4914 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4915 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4916 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4917 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4918 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4919 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4920 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4921 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4922 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4923 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4924 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4925 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4926 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4927 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4928 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4929 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4930 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4931 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4932 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4933 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4934 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4935 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4936 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4937 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4938 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4939 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4940 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4941 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4942 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4943 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4944 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4945 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4946 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4947 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4948 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4949 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4950 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4951 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4952 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4953 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4954 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4955 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4956 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4957 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4958 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4959 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4960 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4961 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4962 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4963 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4964 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4965 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4966 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4967 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4968 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4969 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4970 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4971 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4972 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4973 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4974 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4975 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4976 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4977 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4978 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4979 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4980 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4981 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4982 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4983 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4984 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4985 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4986 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4987 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4988 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4989 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4990 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4991 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4992 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4993 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4994 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4995 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4996 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4997 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4998 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4999 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5000 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5001 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5002 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5003 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5004 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5005 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5006 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5007 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5008 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5009 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5010 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5011 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5012 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5013 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5014 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5015 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5016 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5017 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5018 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5019 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5020 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5021 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5022 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5023 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5024 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5025 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5026 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5027 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5028 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5029 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5030 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5031 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5032 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5033 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5034 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5035 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5036 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5037 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5038 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5039 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5040 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5041 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5042 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5043 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5044 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5045 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5046 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5047 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5048 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5049 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5050 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5051 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5052 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5053 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5054 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5055 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5056 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5057 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5058 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5059 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5060 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5061 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5062 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5063 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5064 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5065 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5066 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5067 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5068 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5069 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5070 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5071 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5072 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5073 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5074 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5075 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5076 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5077 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5078 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5079 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5080 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5081 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5082 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5083 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5084 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5085 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5086 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5087 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5088 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5089 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5090 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5091 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5092 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5093 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5094 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5095 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5096 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5097 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5098 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5099 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5100 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5101 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5102 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5103 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5104 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5105 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5106 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5107 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5108 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5109 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5110 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5111 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5112 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5113 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5114 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5115 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5116 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5117 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5118 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5119 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5120 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5121 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5122 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5123 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5124 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5125 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5126 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5127 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5128 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5129 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5130 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5131 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5132 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5133 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5134 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5135 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5136 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5137 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5138 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5139 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5140 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5141 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5142 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5143 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5144 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5145 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5146 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5147 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5148 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5149 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5150 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5151 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5152 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5153 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5154 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5155 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5156 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5157 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5158 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5159 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5160 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5161 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5162 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5163 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5164 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5165 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5166 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5167 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5168 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5169 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5170 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5171 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5172 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5173 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5174 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5175 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5176 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5177 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5178 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5179 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5180 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5181 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5182 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5183 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5184 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5185 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5186 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5187 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5188 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5189 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5190 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5191 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5192 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5193 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5194 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5195 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5196 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5197 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5198 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5199 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5200 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5201 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5202 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5203 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5204 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5205 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5206 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5207 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5208 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5209 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5210 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5211 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5212 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5213 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5214 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5215 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5216 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5217 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5218 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5219 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5220 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5221 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5222 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5223 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5224 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5225 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5226 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5227 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5228 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5229 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5230 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5231 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5232 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5233 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5234 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5235 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5236 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5237 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5238 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5239 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5240 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5241 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5242 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5243 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5244 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5245 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5246 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5247 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5248 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5249 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5250 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5251 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5252 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5253 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5254 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5255 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5256 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5257 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5258 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5259 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5260 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5261 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5262 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5263 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5264 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5265 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5266 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5267 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5268 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5269 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5270 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5271 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5272 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5273 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5274 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5275 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5276 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5277 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5278 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5279 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5280 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5281 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5282 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5283 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5284 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5285 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5286 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5287 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5288 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5289 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5290 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5291 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5292 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5293 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5294 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5295 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5296 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5297 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5298 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5299 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5300 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5301 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5302 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5303 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5304 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5305 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5306 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5307 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5308 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5309 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5310 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5311 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5312 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5313 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5314 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5315 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5316 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5317 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5318 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5319 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5320 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5321 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5322 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5323 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5324 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5325 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5326 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5327 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5328 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5329 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5330 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5331 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5332 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5333 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5334 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5335 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5336 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5337 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5338 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5339 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5340 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5341 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5342 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5343 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5344 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5345 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5346 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5347 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5348 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5349 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5350 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5351 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5352 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5353 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5354 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5355 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5356 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5357 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5358 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5359 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5360 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5361 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5362 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5363 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5364 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5365 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5366 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5367 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5368 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5369 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5370 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5371 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5372 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5373 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5374 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5375 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5376 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5377 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5378 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5379 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5380 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5381 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5382 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5383 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5384 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5385 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5386 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5387 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5388 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5389 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5390 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5391 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5392 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5393 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5394 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5395 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5396 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5397 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5398 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5399 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5400 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5401 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5402 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5403 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5404 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5405 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5406 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5407 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5408 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5409 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5410 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5411 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5412 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5413 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5414 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5415 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5416 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5417 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5418 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5419 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5420 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5421 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5422 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5423 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5424 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5425 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5426 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5427 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5428 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5429 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5430 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5431 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5432 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5433 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5434 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5435 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5436 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5437 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5438 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5439 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5440 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5441 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5442 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5443 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5444 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5445 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5446 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5447 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5448 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5449 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5450 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5451 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5452 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5453 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5454 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5455 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5456 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5457 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5458 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5459 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5460 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5461 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5462 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5463 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5464 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5465 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5466 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5467 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5468 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5469 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5470 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5471 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5472 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5473 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5474 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5475 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5476 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5477 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5478 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5479 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5480 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5481 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5482 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5483 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5484 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5485 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5486 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5487 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5488 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5489 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5490 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5491 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5492 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5493 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5494 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5495 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5496 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5497 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5498 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5499 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5500 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5501 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5502 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5503 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5504 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5505 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5506 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5507 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5508 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5509 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5510 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5511 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5512 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5513 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5514 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5515 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5516 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5517 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5518 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5519 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5520 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5521 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5522 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5523 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5524 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5525 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5526 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5527 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5528 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5529 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5530 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5531 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5532 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5533 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5534 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5535 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5536 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5537 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5538 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5539 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5540 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5541 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5542 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5543 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5544 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5545 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5546 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5547 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5548 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5549 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5550 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5551 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5552 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5553 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5554 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5555 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5556 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5557 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5558 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5559 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5560 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5561 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5562 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5563 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5564 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5565 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5566 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5567 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5568 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5569 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5570 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5571 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5572 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5573 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5574 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5575 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5576 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5577 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5578 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5579 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5580 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5581 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5582 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5583 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5584 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5585 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5586 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5587 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5588 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5589 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5590 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5591 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5592 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5593 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5594 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5595 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5596 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5597 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5598 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5599 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5600 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5601 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5602 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5603 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5604 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5605 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5606 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5607 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5608 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5609 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5610 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5611 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5612 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5613 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5614 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5615 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5616 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5617 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5618 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5619 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5620 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5621 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5622 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5623 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5624 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5625 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5626 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5627 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5628 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5629 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5630 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5631 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5632 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5633 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5634 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5635 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5636 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5637 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5638 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5639 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5640 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5641 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5642 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5643 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5644 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5645 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5646 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5647 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5648 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5649 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5650 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5651 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5652 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5653 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5654 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5655 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5656 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5657 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5658 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5659 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5660 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5661 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5662 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5663 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5664 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5665 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5666 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5667 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5668 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5669 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5670 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5671 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5672 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5673 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5674 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5675 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5676 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5677 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5678 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5679 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5680 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5681 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5682 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5683 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5684 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5685 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5686 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5687 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5688 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5689 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5690 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5691 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5692 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5693 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5694 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5695 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5696 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5697 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5698 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5699 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5700 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5701 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5702 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5703 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5704 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5705 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5706 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5707 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5708 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5709 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5710 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5711 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5712 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5713 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5714 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5715 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5716 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5717 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5718 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5719 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5720 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5721 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5722 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5723 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5724 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5725 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5726 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5727 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5728 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5729 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5730 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5731 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5732 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5733 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5734 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5735 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5736 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5737 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5738 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5739 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5740 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5741 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5742 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5743 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5744 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5745 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5746 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5747 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5748 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5749 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5750 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5751 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5752 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5753 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5754 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5755 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5756 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5757 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5758 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5759 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5760 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5761 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5762 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5763 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5764 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5765 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5766 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5767 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5768 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5769 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5770 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5771 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5772 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5773 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5774 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5775 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5776 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5777 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5778 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5779 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5780 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5781 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5782 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5783 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5784 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5785 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5786 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5787 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5788 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5789 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5790 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5791 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5792 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5793 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5794 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5795 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5796 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5797 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5798 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5799 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5800 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5801 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5802 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5803 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5804 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5805 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5806 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5807 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5808 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5809 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5810 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5811 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5812 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5813 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5814 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5815 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5816 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5817 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5818 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5819 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5820 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5821 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5822 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5823 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5824 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5825 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5826 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5827 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5828 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5829 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5830 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5831 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5832 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5833 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5834 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5835 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5836 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5837 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5838 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5839 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5840 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5841 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5842 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5843 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5844 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5845 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5846 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5847 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5848 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5849 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5850 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5851 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5852 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5853 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5854 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5855 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5856 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5857 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5858 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5859 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5860 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5861 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5862 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5863 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5864 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5865 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5866 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5867 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5868 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5869 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5870 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5871 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5872 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5873 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5874 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5875 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5876 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5877 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5878 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5879 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5880 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5881 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5882 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5883 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5884 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5885 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5886 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5887 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5888 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5889 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5890 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5891 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5892 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5893 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5894 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5895 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5896 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5897 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5898 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5899 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5900 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5901 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5902 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5903 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5904 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5905 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5906 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5907 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5908 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5909 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5910 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5911 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5912 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5913 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5914 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5915 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5916 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5917 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5918 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5919 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5920 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5921 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5922 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5923 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5924 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5925 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5926 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5927 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5928 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5929 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5930 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5931 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5932 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5933 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5934 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5935 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5936 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5937 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5938 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5939 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5940 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5941 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5942 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5943 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5944 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5945 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5946 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5947 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5948 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5949 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5950 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5951 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5952 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5953 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5954 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5955 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5956 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5957 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5958 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5959 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5960 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5961 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5962 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5963 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5964 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5965 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5966 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5967 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5968 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5969 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5970 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5971 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5972 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5973 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5974 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5975 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5976 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5977 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5978 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5979 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5980 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5981 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5982 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5983 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5984 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5985 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5986 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5987 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5988 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5989 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5990 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5991 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5992 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5993 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5994 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5995 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5996 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5997 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5998 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5999 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6000 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6001 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6002 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6003 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6004 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6005 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6006 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6007 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6008 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6009 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6010 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6011 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6012 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6013 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6014 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6015 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6016 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6017 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6018 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6019 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6020 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6021 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6022 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6023 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6024 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6025 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6026 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6027 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6028 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6029 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6030 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6031 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6032 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6033 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6034 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6035 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6036 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6037 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6038 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6039 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6040 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6041 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6042 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6043 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6044 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6045 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6046 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6047 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6048 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6049 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6050 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6051 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6052 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6053 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6054 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6055 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6056 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6057 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6058 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6059 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6060 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6061 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6062 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6063 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6064 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6065 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6066 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6067 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6068 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6069 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6070 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6071 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6072 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6073 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6074 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6075 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6076 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6077 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6078 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6079 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6080 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6081 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6082 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6083 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6084 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6085 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6086 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6087 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6088 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6089 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6090 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6091 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6092 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6093 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6094 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6095 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6096 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6097 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6098 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6099 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6100 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6101 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6102 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6103 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6104 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6105 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6106 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6107 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6108 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6109 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6110 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6111 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6112 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6113 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6114 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6115 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6116 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6117 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6118 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6119 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6120 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6121 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6122 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6123 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6124 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6125 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6126 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6127 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6128 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6129 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6130 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6131 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6132 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6133 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6134 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6135 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6136 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6137 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6138 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6139 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6140 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6141 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6142 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6143 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6144 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6145 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6146 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6147 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6148 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6149 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6150 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6151 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6152 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6153 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6154 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6155 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6156 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6157 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6158 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6159 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6160 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6161 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6162 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6163 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6164 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6165 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6166 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6167 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6168 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6169 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6170 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6171 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6172 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6173 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6174 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6175 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6176 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6177 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6178 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6179 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6180 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6181 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6182 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6183 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6184 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6185 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6186 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6187 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6188 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6189 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6190 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6191 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6192 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6193 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6194 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6195 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6196 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6197 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6198 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6199 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6200 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6201 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6202 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6203 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6204 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6205 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6206 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6207 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6208 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6209 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6210 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6211 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6212 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6213 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6214 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6215 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6216 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6217 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6218 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6219 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6220 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6221 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6222 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6223 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6224 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6225 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6226 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6227 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6228 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6229 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6230 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6231 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6232 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6233 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6234 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6235 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6236 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6237 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6238 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6239 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6240 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6241 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6242 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6243 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6244 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6245 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6246 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6247 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6248 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6249 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6250 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6251 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6252 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6253 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6254 VREFL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6255 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6256 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6257 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VREFL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6258 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6259 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6260 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6261 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VREFL VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6262 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6263 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6264 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6265 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6266 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6267 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6268 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6269 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6270 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6271 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6272 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6273 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6274 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6275 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6276 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6277 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6278 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6279 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6280 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6281 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6282 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6283 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6284 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6285 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6286 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6287 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6288 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6289 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6290 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6291 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6292 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6293 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6294 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6295 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6296 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6297 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6298 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X6299 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6300 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6301 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X6302 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6303 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6304 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6305 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6306 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6307 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6308 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6309 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6310 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6311 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D20 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6312 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6313 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D20 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6314 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6315 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6316 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6317 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6318 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6319 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D21 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6320 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6321 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D21 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6322 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6323 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6324 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6325 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6326 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6327 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D22 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6328 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6329 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D22 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6330 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6331 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6332 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6333 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6334 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6335 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D23 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6336 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6337 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D23 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6338 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6339 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6340 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6341 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6342 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6343 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D24 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6344 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6345 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D24 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6346 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6347 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6348 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6349 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6350 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6351 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D25 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6352 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6353 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D25 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6354 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6355 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6356 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6357 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6358 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6359 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D26 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6360 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6361 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D26 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6362 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6363 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6364 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6365 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6366 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6367 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D27 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X6368 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6369 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D27 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X6370 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1549_3140# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0 ps=0 w=2 l=0.5
X6371 VOUT2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=3.48 pd=25.2 as=0 ps=0 w=6 l=0.5
X6372 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VOUT2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X6373 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X6374 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1095_1321# VOUT2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_937_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=13.2 as=0.58 ps=4.58 w=2 l=0.5
X6375 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VOUT2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X6376 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6377 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=9.16 w=2 l=0.5
R6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VSSA sky130_fd_pr__res_generic_po w=0.33 l=65.2
X6378 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0.58 ps=4.58 w=2 l=0.5
X6379 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1549_3140# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6380 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VOUT2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=5.8 ps=41.2 w=10 l=0.5
X6381 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1549_3140# VOUT2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1392_2207# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6382 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1095_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X6383 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1095_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
X6384 VOUT2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X6385 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=1.74 ps=13.2 w=2 l=0.5
X6386 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6387 VOUT2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X6388 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
R7 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# sky130_fd_pr__res_generic_po w=0.33 l=38.5
X6389 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
X6390 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_550_1291# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6391 VOUT2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X6392 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VOUT2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X6393 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=9.16 as=0 ps=0 w=2 l=0.5
X6394 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X6395 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X6396 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
R8 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_n804_1718# VSSA sky130_fd_pr__res_generic_po w=0.33 l=23.6
X6397 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_1473_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X6398 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2388_2094# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[0]/opamp_0/a_2168_2788# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X6399 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6400 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6401 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6402 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6403 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6404 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6405 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6406 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6407 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6408 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6409 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6410 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6411 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6412 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6413 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6414 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6415 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6416 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6417 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6418 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6419 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6420 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6421 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6422 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6423 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6424 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6425 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6426 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6427 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6428 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6429 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6430 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6431 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6432 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6433 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6434 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6435 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6436 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6437 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6438 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6439 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6440 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6441 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6442 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6443 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6444 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6445 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6446 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6447 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6448 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6449 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6450 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6451 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6452 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6453 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6454 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6455 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6456 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6457 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6458 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6459 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6460 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6461 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6462 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6463 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6464 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6465 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6466 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6467 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6468 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6469 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6470 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6471 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6472 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6473 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6474 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6475 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6476 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6477 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6478 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6479 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6480 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6481 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6482 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6483 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6484 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6485 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6486 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6487 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6488 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6489 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6490 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6491 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6492 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6493 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6494 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6495 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6496 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6497 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6498 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6499 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6500 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6501 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6502 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6503 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6504 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6505 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6506 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6507 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6508 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6509 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6510 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6511 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6512 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6513 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6514 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6515 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6516 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6517 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6518 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6519 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6520 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6521 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6522 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6523 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6524 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6525 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6526 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6527 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6528 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6529 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6530 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6531 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6532 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6533 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6534 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6535 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6536 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6537 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6538 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6539 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6540 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6541 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6542 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6543 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6544 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6545 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6546 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6547 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6548 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6549 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6550 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6551 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6552 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6553 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6554 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6555 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6556 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6557 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6558 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6559 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6560 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6561 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6562 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6563 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6564 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6565 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6566 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6567 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6568 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6569 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6570 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6571 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6572 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6573 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6574 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6575 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6576 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6577 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6578 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6579 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6580 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6581 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6582 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6583 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6584 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6585 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6586 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6587 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6588 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6589 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6590 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6591 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6592 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6593 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6594 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6595 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6596 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6597 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6598 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6599 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6600 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6601 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6602 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6603 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6604 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6605 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6606 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6607 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6608 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6609 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6610 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6611 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6612 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6613 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6614 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6615 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6616 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6617 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6618 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6619 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6620 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6621 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6622 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6623 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6624 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6625 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6626 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6627 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6628 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6629 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6630 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6631 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6632 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6633 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6634 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6635 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6636 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6637 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6638 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6639 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6640 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6641 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6642 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6643 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6644 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6645 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6646 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6647 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6648 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6649 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6650 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6651 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6652 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6653 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6654 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6655 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6656 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6657 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6658 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6659 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6660 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6661 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6662 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6663 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6664 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6665 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6666 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6667 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6668 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6669 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6670 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6671 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6672 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6673 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6674 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6675 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6676 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6677 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6678 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6679 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6680 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6681 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6682 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6683 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6684 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6685 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6686 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6687 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6688 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6689 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6690 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6691 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6692 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6693 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6694 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6695 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6696 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6697 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6698 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6699 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6700 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6701 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6702 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6703 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6704 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6705 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6706 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6707 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6708 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6709 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6710 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6711 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6712 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6713 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6714 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6715 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6716 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6717 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6718 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6719 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6720 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6721 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6722 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6723 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6724 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6725 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6726 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6727 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6728 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6729 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6730 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6731 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6732 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6733 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6734 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6735 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6736 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6737 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6738 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6739 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6740 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6741 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6742 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6743 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6744 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6745 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6746 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6747 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6748 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6749 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6750 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6751 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6752 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6753 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6754 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6755 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6756 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6757 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6758 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6759 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6760 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6761 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6762 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6763 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6764 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6765 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6766 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6767 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6768 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6769 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6770 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6771 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6772 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6773 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6774 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6775 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6776 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6777 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6778 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6779 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6780 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6781 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6782 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6783 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6784 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6785 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6786 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6787 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6788 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6789 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6790 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6791 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6792 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6793 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6794 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6795 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6796 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6797 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6798 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6799 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6800 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6801 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6802 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6803 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6804 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6805 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6806 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6807 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6808 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6809 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6810 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6811 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6812 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6813 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6814 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6815 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6816 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6817 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6818 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6819 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6820 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6821 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6822 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6823 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6824 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6825 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6826 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6827 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6828 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6829 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6830 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6831 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6832 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6833 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6834 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6835 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6836 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6837 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6838 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6839 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6840 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6841 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6842 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6843 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6844 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6845 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6846 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6847 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6848 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6849 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6850 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6851 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6852 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6853 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6854 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6855 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6856 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6857 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6858 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6859 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6860 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6861 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6862 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6863 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6864 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6865 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6866 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6867 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6868 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6869 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6870 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6871 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6872 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6873 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6874 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6875 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6876 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6877 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6878 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6879 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6880 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6881 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6882 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6883 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6884 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6885 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6886 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6887 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6888 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6889 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6890 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6891 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6892 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6893 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6894 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6895 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6896 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6897 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6898 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6899 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6900 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6901 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6902 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6903 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6904 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6905 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6906 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6907 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6908 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6909 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6910 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6911 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6912 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6913 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6914 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6915 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6916 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6917 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6918 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6919 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6920 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6921 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6922 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6923 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6924 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6925 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6926 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6927 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6928 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6929 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6930 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6931 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6932 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6933 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6934 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6935 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6936 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6937 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6938 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6939 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6940 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6941 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6942 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6943 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6944 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6945 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6946 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6947 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6948 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6949 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6950 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6951 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6952 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6953 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6954 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6955 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6956 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6957 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6958 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6959 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6960 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6961 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6962 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6963 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6964 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6965 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6966 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6967 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6968 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6969 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6970 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6971 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6972 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6973 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6974 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6975 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6976 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6977 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6978 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6979 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6980 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6981 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6982 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6983 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6984 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6985 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6986 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6987 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6988 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6989 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6990 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6991 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6992 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6993 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6994 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6995 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6996 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6997 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6998 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6999 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7000 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7001 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7002 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7003 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7004 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7005 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7006 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7007 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7008 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7009 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7010 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7011 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7012 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7013 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7014 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7015 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7016 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7017 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7018 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7019 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7020 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7021 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7022 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7023 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7024 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7025 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7026 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7027 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7028 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7029 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7030 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7031 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7032 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7033 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7034 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7035 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7036 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7037 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7038 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7039 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7040 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7041 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7042 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7043 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7044 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7045 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7046 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7047 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7048 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7049 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7050 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7051 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7052 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7053 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7054 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7055 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7056 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7057 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7058 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7059 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7060 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7061 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7062 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7063 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7064 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7065 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7066 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7067 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7068 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7069 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7070 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7071 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7072 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7073 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7074 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7075 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7076 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7077 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7078 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7079 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7080 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7081 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7082 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7083 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7084 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7085 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7086 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7087 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7088 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7089 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7090 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7091 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7092 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7093 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7094 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7095 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7096 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7097 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7098 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7099 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7100 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7101 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7102 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7103 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7104 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7105 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7106 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7107 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7108 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7109 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7110 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7111 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7112 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7113 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7114 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7115 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7116 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7117 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7118 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7119 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7120 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7121 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7122 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7123 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7124 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7125 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7126 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7127 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7128 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7129 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7130 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7131 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7132 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7133 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7134 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7135 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7136 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7137 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7138 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7139 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7140 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7141 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7142 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7143 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7144 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7145 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7146 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7147 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7148 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7149 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7150 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7151 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7152 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7153 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7154 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7155 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7156 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7157 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7158 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7159 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7160 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7161 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7162 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7163 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7164 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7165 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7166 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7167 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7168 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7169 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7170 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7171 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7172 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7173 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7174 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7175 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7176 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7177 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7178 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7179 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7180 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7181 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7182 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7183 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7184 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7185 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7186 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7187 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7188 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7189 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7190 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7191 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7192 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7193 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7194 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7195 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7196 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7197 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7198 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7199 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7200 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7201 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7202 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7203 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7204 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7205 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7206 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7207 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7208 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7209 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7210 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7211 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7212 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7213 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7214 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7215 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7216 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7217 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7218 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7219 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7220 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7221 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7222 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7223 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7224 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7225 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7226 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7227 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7228 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7229 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7230 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7231 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7232 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7233 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7234 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7235 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7236 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7237 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7238 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7239 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7240 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7241 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7242 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7243 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7244 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7245 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7246 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7247 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7248 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7249 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7250 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7251 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7252 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7253 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7254 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7255 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7256 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7257 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7258 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7259 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7260 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7261 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7262 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7263 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7264 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7265 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7266 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7267 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7268 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7269 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7270 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7271 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7272 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7273 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7274 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7275 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7276 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7277 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7278 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7279 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7280 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7281 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7282 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7283 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7284 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7285 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7286 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7287 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7288 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7289 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7290 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7291 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7292 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7293 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7294 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7295 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7296 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7297 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7298 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7299 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7300 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7301 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7302 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7303 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7304 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7305 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7306 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7307 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7308 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7309 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7310 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7311 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7312 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7313 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7314 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7315 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7316 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7317 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7318 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7319 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7320 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7321 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7322 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7323 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7324 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7325 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7326 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7327 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7328 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7329 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7330 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7331 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7332 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7333 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7334 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7335 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7336 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7337 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7338 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7339 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7340 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7341 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7342 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7343 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7344 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7345 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7346 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7347 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7348 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7349 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7350 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7351 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7352 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7353 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7354 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7355 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7356 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7357 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7358 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7359 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7360 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7361 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7362 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7363 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7364 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7365 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7366 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7367 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7368 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7369 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7370 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7371 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7372 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7373 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7374 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7375 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7376 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7377 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7378 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7379 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7380 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7381 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7382 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7383 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7384 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7385 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7386 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7387 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7388 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7389 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7390 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7391 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7392 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7393 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7394 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7395 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7396 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7397 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7398 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7399 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7400 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7401 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7402 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7403 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7404 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7405 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7406 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7407 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7408 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7409 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7410 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7411 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7412 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7413 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7414 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7415 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7416 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7417 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7418 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7419 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7420 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7421 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7422 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7423 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7424 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7425 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7426 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7427 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7428 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7429 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7430 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7431 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7432 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7433 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7434 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7435 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7436 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7437 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7438 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7439 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7440 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7441 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7442 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7443 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7444 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7445 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7446 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7447 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7448 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7449 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7450 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7451 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7452 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7453 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7454 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7455 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7456 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7457 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7458 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7459 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7460 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7461 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7462 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7463 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7464 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7465 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7466 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7467 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7468 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7469 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7470 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7471 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7472 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7473 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7474 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7475 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7476 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7477 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7478 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7479 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7480 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7481 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7482 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7483 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7484 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7485 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7486 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7487 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7488 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7489 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7490 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7491 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7492 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7493 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7494 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7495 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7496 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7497 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7498 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7499 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7500 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7501 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7502 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7503 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7504 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7505 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7506 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7507 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7508 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7509 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7510 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7511 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7512 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7513 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7514 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7515 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7516 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7517 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7518 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7519 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7520 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7521 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7522 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7523 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7524 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7525 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7526 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7527 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7528 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7529 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7530 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7531 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7532 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7533 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7534 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7535 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7536 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7537 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7538 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7539 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7540 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7541 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7542 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7543 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7544 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7545 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7546 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7547 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7548 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7549 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7550 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7551 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7552 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7553 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7554 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7555 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7556 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7557 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7558 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7559 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7560 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7561 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7562 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7563 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7564 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7565 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7566 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7567 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7568 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7569 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7570 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7571 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7572 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7573 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7574 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7575 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7576 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7577 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7578 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7579 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7580 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7581 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7582 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7583 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7584 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7585 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7586 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7587 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7588 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7589 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7590 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7591 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7592 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7593 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7594 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7595 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7596 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7597 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7598 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7599 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7600 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7601 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7602 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7603 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7604 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7605 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7606 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7607 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7608 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7609 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7610 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7611 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7612 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7613 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7614 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7615 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7616 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7617 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7618 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7619 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7620 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7621 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7622 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7623 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7624 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7625 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7626 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7627 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7628 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7629 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7630 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7631 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7632 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7633 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7634 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7635 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7636 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7637 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7638 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7639 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7640 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7641 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7642 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7643 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7644 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7645 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7646 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7647 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7648 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7649 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7650 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7651 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7652 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7653 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7654 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7655 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7656 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7657 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7658 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7659 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7660 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7661 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7662 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7663 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7664 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7665 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7666 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7667 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7668 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7669 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7670 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7671 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7672 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7673 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7674 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7675 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7676 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7677 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7678 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7679 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7680 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7681 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7682 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7683 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7684 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7685 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7686 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7687 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7688 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7689 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7690 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7691 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7692 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7693 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7694 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7695 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7696 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7697 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7698 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7699 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7700 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7701 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7702 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7703 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7704 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7705 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7706 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7707 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7708 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7709 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7710 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7711 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7712 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7713 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7714 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7715 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7716 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7717 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7718 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7719 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7720 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7721 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7722 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7723 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7724 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7725 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7726 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7727 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7728 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7729 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7730 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7731 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7732 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7733 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7734 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7735 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7736 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7737 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7738 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7739 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7740 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7741 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7742 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7743 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7744 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7745 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7746 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7747 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7748 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7749 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7750 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7751 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7752 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7753 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7754 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7755 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7756 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7757 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7758 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7759 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7760 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7761 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7762 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7763 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7764 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7765 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7766 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7767 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7768 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7769 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7770 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7771 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7772 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7773 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7774 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7775 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7776 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7777 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7778 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7779 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7780 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7781 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7782 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7783 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7784 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7785 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7786 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7787 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7788 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7789 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7790 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7791 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7792 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7793 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7794 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7795 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7796 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7797 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7798 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7799 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7800 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7801 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7802 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7803 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7804 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7805 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7806 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7807 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7808 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7809 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7810 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7811 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7812 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7813 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7814 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7815 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7816 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7817 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7818 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7819 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7820 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7821 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7822 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7823 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7824 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7825 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7826 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7827 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7828 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7829 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7830 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7831 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7832 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7833 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7834 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7835 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7836 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7837 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7838 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7839 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7840 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7841 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7842 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7843 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7844 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7845 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7846 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7847 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7848 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7849 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7850 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7851 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7852 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7853 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7854 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7855 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7856 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7857 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7858 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7859 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7860 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7861 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7862 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7863 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7864 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7865 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7866 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7867 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7868 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7869 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7870 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7871 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7872 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7873 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7874 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7875 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7876 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7877 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7878 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7879 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7880 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7881 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7882 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7883 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7884 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7885 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7886 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7887 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7888 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7889 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7890 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7891 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7892 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7893 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7894 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7895 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7896 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7897 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7898 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7899 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7900 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7901 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7902 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7903 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7904 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7905 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7906 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7907 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7908 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7909 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7910 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7911 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7912 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7913 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7914 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7915 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7916 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7917 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7918 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7919 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7920 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7921 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7922 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7923 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7924 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7925 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7926 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7927 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7928 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7929 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7930 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7931 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7932 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7933 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7934 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7935 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7936 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7937 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7938 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7939 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7940 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7941 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7942 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7943 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7944 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7945 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7946 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7947 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7948 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7949 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7950 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7951 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7952 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7953 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7954 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7955 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7956 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7957 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7958 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7959 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7960 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7961 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7962 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7963 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7964 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7965 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7966 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7967 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7968 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7969 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7970 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7971 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7972 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7973 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7974 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7975 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7976 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7977 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7978 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7979 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7980 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7981 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7982 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7983 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7984 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7985 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7986 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7987 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7988 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7989 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7990 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7991 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7992 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7993 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7994 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7995 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7996 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7997 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7998 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7999 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8000 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8001 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8002 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8003 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8004 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8005 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8006 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8007 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8008 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8009 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8010 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8011 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8012 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8013 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8014 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8015 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8016 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8017 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8018 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8019 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8020 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8021 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8022 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8023 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8024 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8025 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8026 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8027 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8028 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8029 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8030 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8031 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8032 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8033 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8034 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8035 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8036 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8037 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8038 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8039 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8040 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8041 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8042 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8043 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8044 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8045 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8046 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8047 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8048 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8049 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8050 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8051 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8052 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8053 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8054 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8055 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8056 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8057 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8058 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8059 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8060 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8061 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8062 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8063 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8064 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8065 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8066 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8067 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8068 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8069 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8070 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8071 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8072 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8073 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8074 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8075 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8076 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8077 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8078 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8079 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8080 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8081 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8082 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8083 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8084 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8085 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8086 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8087 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8088 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8089 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8090 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8091 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8092 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8093 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8094 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8095 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8096 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8097 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8098 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8099 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8100 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8101 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8102 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8103 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8104 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8105 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8106 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8107 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8108 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8109 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8110 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8111 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8112 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8113 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8114 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8115 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8116 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8117 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8118 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8119 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8120 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8121 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8122 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8123 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8124 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8125 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8126 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8127 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8128 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8129 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8130 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8131 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8132 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8133 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8134 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8135 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8136 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8137 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8138 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8139 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8140 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8141 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8142 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8143 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8144 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8145 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8146 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8147 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8148 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8149 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8150 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8151 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8152 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8153 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8154 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8155 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8156 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8157 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8158 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8159 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8160 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8161 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8162 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8163 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8164 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8165 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8166 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8167 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8168 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8169 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8170 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8171 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8172 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8173 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8174 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8175 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8176 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8177 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8178 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8179 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8180 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8181 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8182 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8183 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8184 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8185 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8186 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8187 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8188 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8189 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8190 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8191 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8192 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8193 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8194 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8195 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8196 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8197 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8198 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8199 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8200 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8201 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8202 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8203 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8204 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8205 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8206 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8207 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8208 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8209 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8210 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8211 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8212 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8213 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8214 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8215 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8216 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8217 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8218 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8219 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8220 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8221 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8222 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8223 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8224 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8225 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8226 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8227 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8228 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8229 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8230 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8231 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8232 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8233 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8234 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8235 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8236 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8237 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8238 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8239 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8240 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8241 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8242 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8243 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8244 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8245 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8246 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8247 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8248 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8249 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8250 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8251 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8252 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8253 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8254 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8255 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8256 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8257 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8258 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8259 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8260 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8261 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8262 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8263 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8264 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8265 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8266 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8267 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8268 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8269 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8270 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8271 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8272 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8273 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8274 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8275 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8276 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8277 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8278 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8279 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8280 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8281 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8282 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8283 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8284 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8285 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8286 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8287 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8288 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8289 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8290 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8291 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8292 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8293 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8294 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8295 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8296 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8297 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8298 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8299 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8300 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8301 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8302 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8303 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8304 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8305 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8306 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8307 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8308 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8309 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8310 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8311 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8312 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8313 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8314 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8315 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8316 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8317 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8318 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8319 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8320 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8321 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8322 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8323 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8324 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8325 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8326 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8327 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8328 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8329 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8330 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8331 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8332 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8333 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8334 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8335 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8336 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8337 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8338 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8339 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8340 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8341 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8342 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8343 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8344 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8345 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8346 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8347 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8348 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8349 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8350 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8351 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8352 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8353 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8354 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8355 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8356 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8357 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8358 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8359 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8360 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8361 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8362 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8363 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8364 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8365 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8366 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8367 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8368 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8369 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8370 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8371 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8372 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8373 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8374 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8375 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8376 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8377 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8378 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8379 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8380 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8381 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8382 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8383 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8384 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8385 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8386 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8387 VREFL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8388 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8389 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8390 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VREFL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8391 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8392 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8393 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8394 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VREFL VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8395 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8396 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8397 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8398 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8399 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8400 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8401 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8402 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8403 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8404 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8405 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8406 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8407 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8408 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8409 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8410 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8411 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8412 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8413 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8414 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8415 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8416 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8417 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8418 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8419 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8420 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8421 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8422 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8423 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8424 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8425 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8426 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8427 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8428 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8429 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8430 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8431 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X8432 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8433 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8434 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X8435 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8436 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8437 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7_BUF 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8438 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8439 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8440 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8441 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8442 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8443 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8444 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D30 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8445 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8446 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1810_540# D30 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8447 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8448 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8449 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8450 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8451 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8452 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D31 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8453 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8454 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1810_540# D31 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8455 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8456 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8457 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8458 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8459 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8460 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D32 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8461 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8462 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1810_540# D32 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8463 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8464 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8465 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8466 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8467 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8468 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D33 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8469 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8470 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1810_540# D33 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8471 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8472 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8473 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8474 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8475 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8476 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D34 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8477 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8478 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1810_540# D34 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8479 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8480 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8481 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8482 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8483 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8484 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D35 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8485 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8486 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1810_540# D35 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8487 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8488 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8489 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8490 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8491 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8492 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D36 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8493 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8494 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1810_540# D36 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8495 VSSD 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8496 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8497 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8498 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8499 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1428_490# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8500 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D37 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0 ps=0 w=0.84 l=0.15
X8501 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1600_540# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8502 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1810_540# D37 VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0 ps=0 w=0.42 l=0.15
X8503 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1549_3140# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0 ps=0 w=2 l=0.5
X8504 VOUT3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=3.48 pd=25.2 as=0 ps=0 w=6 l=0.5
X8505 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VOUT3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X8506 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X8507 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1095_1321# VOUT3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_937_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=13.2 as=0.58 ps=4.58 w=2 l=0.5
X8508 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VOUT3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X8509 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8510 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=9.16 w=2 l=0.5
R9 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VSSA sky130_fd_pr__res_generic_po w=0.33 l=65.2
X8511 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0.58 ps=4.58 w=2 l=0.5
X8512 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1549_3140# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
X8513 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VOUT3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=5.8 ps=41.2 w=10 l=0.5
X8514 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1549_3140# VOUT3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1392_2207# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8515 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/VIN 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1095_1321# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X8516 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1095_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
X8517 VOUT3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=6 l=0.5
X8518 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=1.74 ps=13.2 w=2 l=0.5
X8519 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8520 VOUT3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X8521 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1253_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
R10 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# sky130_fd_pr__res_generic_po w=0.33 l=38.5
X8522 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_937_1321# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=0.5
X8523 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_550_1291# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8524 VOUT3 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X8525 VDDA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VOUT3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
X8526 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_925_2276# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=9.16 as=0 ps=0 w=2 l=0.5
X8527 VSSA 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X8528 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1392_2207# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X8529 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1708_2207# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
R11 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_n804_1718# VSSA sky130_fd_pr__res_generic_po w=0.33 l=23.6
X8530 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2027_304# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_1473_304# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X8531 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2388_2094# 2x8bit_tx_buffer_0[1]/8_bit_dac_tx_buffer_v2_0[1]/opamp_0/a_2168_2788# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.5
.ends
*******************************************************
X1 D00 D01 D02 D03 D04 D05 D06 D07 D10 D11 D12 D13 D14 D15
+ D16 D17 D20 D21 D22 D23 D24 D25 D26 D27 D30 D31 D32 D33 D34 D35 D36 D37 VCCD VDDA
+ VOUT0 VOUT1 VOUT2 VOUT3 VREFH VREFL VSSA VSSD x4x8bit_tx_buffer
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


V1 VDDA 0 dc 3.3
V2 VSSA 0 dc 0
V3 VCCD 0 dc 1.8
V4 VSSD 0 dc 0
V5 VREFL 0 dc 0
V6 VREFH 0 dc 3.3

V7 D00 0 pulse(0 1.8 0ns 0.1ns 0.1ns 1us 2us)
V8 D01 0 pulse(0 1.8 0ns 0.1ns 0.1ns 2us 4us)
V9 D02 0 pulse(0 1.8 0ns 0.1ns 0.1ns 4us 8us)
V10 D03 0 pulse(0 1.8 0ns 0.1ns 0.1ns 8us 16us)
V11 D04 0 pulse(0 1.8 0ns 0.1ns 0.1ns 16us 32us)
V12 D05 0 pulse(0 1.8 0ns 0.1ns 0.1ns 32us 64us)
V13 D06 0 pulse(0 1.8 0ns 0.1ns 0.1ns 64us 128us)
V14 D07 0 pulse(0 1.8 0ns 0.1ns 0.1ns 128us 256us)

V15 D10 0 pulse(0 1.8 1us 0.1ns 0.1ns 1us 2us)
V16 D11 0 pulse(0 1.8 2us 0.1ns 0.1ns 2us 4us)
V17 D12 0 pulse(0 1.8 4us 0.1ns 0.1ns 4us 8us)
V18 D13 0 pulse(0 1.8 8us 0.1ns 0.1ns 8us 16us)
V19 D14 0 pulse(0 1.8 16us 0.1ns 0.1ns 16us 32us)
V20 D15 0 pulse(0 1.8 32us 0.1ns 0.1ns 32us 64us)
V21 D16 0 pulse(0 1.8 64us 0.1ns 0.1ns 64us 128us)
V22 D17 0 pulse(0 1.8 128us 0.1ns 0.1ns 128us 256us)

V23 D20 0 pulse(0 1.8 0ns 0.1ns 0.1ns 1us 2us)
V24 D21 0 pulse(0 1.8 0ns 0.1ns 0.1ns 2us 4us)
V25 D22 0 pulse(0 1.8 0ns 0.1ns 0.1ns 4us 8us)
V26 D23 0 pulse(0 1.8 0ns 0.1ns 0.1ns 8us 16us)
V27 D24 0 pulse(0 1.8 0ns 0.1ns 0.1ns 16us 32us)
V28 D25 0 pulse(0 1.8 0ns 0.1ns 0.1ns 32us 64us)
V29 D26 0 pulse(0 1.8 0ns 0.1ns 0.1ns 64us 128us)
V30 D27 0 pulse(0 1.8 0ns 0.1ns 0.1ns 128us 256us)

V31 D30 0 pulse(0 1.8 1us 0.1ns 0.1ns 1us 2us)
V32 D31 0 pulse(0 1.8 2us 0.1ns 0.1ns 2us 4us)
V33 D32 0 pulse(0 1.8 4us 0.1ns 0.1ns 4us 8us)
V34 D33 0 pulse(0 1.8 8us 0.1ns 0.1ns 8us 16us)
V35 D34 0 pulse(0 1.8 16us 0.1ns 0.1ns 16us 32us)
V36 D35 0 pulse(0 1.8 32us 0.1ns 0.1ns 32us 64us)
V37 D36 0 pulse(0 1.8 64us 0.1ns 0.1ns 64us 128us)
V38 D37 0 pulse(0 1.8 128us 0.1ns 0.1ns 128us 256us)

.tran 5u 50u
.control
run
plot VOUT0 VOUT1 VOUT2 VOUT3
.endc
.end
