magic
tech sky130A
magscale 1 2
timestamp 1686560844
<< locali >>
rect 0 78948 506 79088
rect 0 0 652 140
<< metal2 >>
rect 745 85717 779 85823
rect 848 85699 882 85828
rect 946 85685 980 85828
rect 1050 85697 1084 85828
rect 1158 85683 1192 85828
rect 1258 85679 1292 85828
rect 1366 85675 1400 85828
rect 1478 85679 1512 85828
rect 9265 85552 9373 85828
rect 11346 85719 11380 85828
rect 11449 85729 11483 85828
rect 11547 85721 11581 85828
rect 11651 85731 11685 85828
rect 11759 85717 11793 85828
rect 11859 85711 11893 85828
rect 11967 85713 12001 85828
rect 12079 85721 12113 85828
rect 19866 85634 19974 85828
rect 21947 85739 21981 85828
rect 22050 85725 22084 85828
rect 22148 85717 22182 85828
rect 22252 85725 22286 85828
rect 22360 85709 22394 85828
rect 22460 85695 22494 85828
rect 22568 85705 22602 85828
rect 22680 85711 22714 85828
rect 30467 85636 30575 85828
rect 32548 85721 32582 85828
rect 32651 85719 32685 85828
rect 32749 85735 32783 85828
rect 32853 85737 32887 85828
rect 32961 85729 32995 85828
rect 33061 85711 33095 85828
rect 33169 85713 33203 85828
rect 33281 85699 33315 85828
rect 41068 85610 41176 85828
<< metal3 >>
rect 0 85389 314 85489
rect 0 81638 628 81738
rect 0 80127 260 80227
rect 2 79395 358 79495
rect 0 78454 42404 78594
rect 0 77764 42404 77904
rect 0 77226 42404 77366
rect 0 76536 42404 76676
rect 0 75998 42404 76138
rect 0 75308 42404 75448
rect 0 74770 42404 74910
rect 0 74080 42404 74220
rect 0 73542 42404 73682
rect 0 72852 42404 72992
rect 0 72314 42404 72454
rect 0 71624 42404 71764
rect 0 71086 42404 71226
rect 0 70396 42404 70536
rect 0 69858 42404 69998
rect 0 69168 42404 69308
rect 0 68630 42404 68770
rect 0 67940 42404 68080
rect 0 67402 42404 67542
rect 0 66712 42404 66852
rect 0 66174 42404 66314
rect 0 65484 42404 65624
rect 0 64946 42404 65086
rect 0 64256 42404 64396
rect 0 63718 42404 63858
rect 0 63028 42404 63168
rect 0 62490 42404 62630
rect 0 61800 42404 61940
rect 0 61262 42404 61402
rect 0 60572 42404 60712
rect 0 60034 42404 60174
rect 0 59344 42404 59484
rect 0 58806 42404 58946
rect 0 58116 42404 58256
rect 0 57578 42404 57718
rect 0 56888 42404 57028
rect 0 56350 42404 56490
rect 0 55660 42404 55800
rect 0 55122 42404 55262
rect 0 54432 42404 54572
rect 0 53894 42404 54034
rect 0 53204 42404 53344
rect 0 52666 42404 52806
rect 0 51976 42404 52116
rect 0 51438 42404 51578
rect 0 50748 42404 50888
rect 0 50210 42404 50350
rect 0 49520 42404 49660
rect 0 48982 42404 49122
rect 0 48292 42404 48432
rect 0 47754 42404 47894
rect 0 47064 42404 47204
rect 0 46526 42404 46666
rect 0 45836 42404 45976
rect 0 45298 42404 45438
rect 0 44608 42404 44748
rect 0 44070 42404 44210
rect 0 43380 42404 43520
rect 0 42842 42404 42982
rect 0 42152 42404 42292
rect 0 41614 42404 41754
rect 0 40924 42404 41064
rect 0 40386 42404 40526
rect 0 39696 42404 39836
rect 0 39158 42404 39298
rect 0 38468 42404 38608
rect 0 37930 42404 38070
rect 0 37240 42404 37380
rect 0 36702 42404 36842
rect 0 36012 42404 36152
rect 0 35474 42404 35614
rect 0 34784 42404 34924
rect 0 34246 42404 34386
rect 0 33556 42404 33696
rect 0 33018 42404 33158
rect 0 32328 42404 32468
rect 0 31790 42404 31930
rect 0 31100 42404 31240
rect 0 30562 42404 30702
rect 0 29872 42404 30012
rect 0 29334 42404 29474
rect 0 28644 42404 28784
rect 0 28106 42404 28246
rect 0 27416 42404 27556
rect 0 26878 42404 27018
rect 0 26188 42404 26328
rect 0 25650 42404 25790
rect 0 24960 42404 25100
rect 0 24422 42404 24562
rect 0 23732 42404 23872
rect 0 23194 42404 23334
rect 0 22504 42404 22644
rect 0 21966 42404 22106
rect 0 21276 42404 21416
rect 0 20738 42404 20878
rect 0 20048 42404 20188
rect 0 19510 42404 19650
rect 0 18820 42404 18960
rect 0 18282 42404 18422
rect 0 17592 42404 17732
rect 0 17054 42404 17194
rect 0 16364 42404 16504
rect 0 15826 42404 15966
rect 0 15136 42404 15276
rect 0 14598 42404 14738
rect 0 13908 42404 14048
rect 0 13370 42404 13510
rect 0 12680 42404 12820
rect 0 12142 42404 12282
rect 0 11452 42404 11592
rect 0 10914 42404 11054
rect 0 10224 42404 10364
rect 0 9686 42404 9826
rect 0 8996 42404 9136
rect 0 8458 42404 8598
rect 0 7768 42404 7908
rect 0 7230 42404 7370
rect 0 6540 42404 6680
rect 0 6002 42404 6142
rect 0 5312 42404 5452
rect 0 4774 42404 4914
rect 0 4084 42404 4224
rect 0 3546 42404 3686
rect 0 2856 42404 2996
rect 0 2318 42404 2458
rect 0 1628 42404 1768
rect 0 1090 42404 1230
rect 0 400 42404 540
use 2x8bit_tx_buffer  2x8bit_tx_buffer_0
array 0 1 21202 0 0 85828
timestamp 1686481404
transform 1 0 0 0 1 0
box 0 0 21202 85828
<< labels >>
flabel metal2 s 762 85778 762 85778 1 FreeSans 480 0 0 160 D00
flabel metal2 s 864 85792 864 85792 1 FreeSans 480 0 0 160 D01
flabel metal2 s 960 85794 960 85794 1 FreeSans 480 0 0 160 D02
flabel metal2 s 1064 85802 1064 85802 1 FreeSans 480 0 0 160 D03
flabel metal2 s 1180 85798 1180 85798 1 FreeSans 480 0 0 160 D04
flabel metal2 s 1270 85794 1270 85794 1 FreeSans 480 0 0 160 D05
flabel metal2 s 1380 85798 1380 85798 1 FreeSans 480 0 0 160 D06
flabel metal2 s 1502 85790 1502 85790 1 FreeSans 480 0 0 160 D07
flabel metal2 s 9316 85740 9316 85740 1 FreeSans 480 0 0 160 VOUT0
flabel metal2 s 11364 85794 11364 85794 1 FreeSans 480 0 0 160 D10
flabel metal2 s 11468 85798 11468 85798 1 FreeSans 480 0 0 160 D11
flabel metal2 s 11562 85800 11562 85800 1 FreeSans 480 0 0 160 D12
flabel metal2 s 11668 85806 11668 85806 1 FreeSans 480 0 0 160 D13
flabel metal2 s 11788 85816 11788 85816 1 FreeSans 480 0 0 160 D14
flabel metal2 s 11880 85800 11880 85800 1 FreeSans 480 0 0 160 D15
flabel metal2 s 11980 85794 11980 85794 1 FreeSans 480 0 0 160 D16
flabel metal2 s 12106 85810 12106 85810 1 FreeSans 480 0 0 160 D17
flabel metal2 s 19916 85762 19916 85762 1 FreeSans 480 0 0 160 VOUT1
flabel metal2 s 21960 85818 21960 85818 1 FreeSans 480 0 0 160 D20
flabel metal2 s 22078 85816 22078 85816 1 FreeSans 480 0 0 160 D21
flabel metal2 s 22166 85816 22166 85816 1 FreeSans 480 0 0 160 D22
flabel metal2 s 22282 85814 22282 85814 1 FreeSans 480 0 0 160 D23
flabel metal2 s 22380 85818 22380 85818 1 FreeSans 480 0 0 160 D24
flabel metal2 s 22486 85810 22486 85810 1 FreeSans 480 0 0 160 D25
flabel metal2 s 22586 85818 22586 85818 1 FreeSans 480 0 0 160 D26
flabel metal2 s 22702 85808 22702 85808 1 FreeSans 480 0 0 160 D27
flabel metal2 s 30536 85804 30536 85804 1 FreeSans 480 0 0 160 VOUT2
flabel metal2 s 32562 85818 32562 85818 1 FreeSans 480 0 0 160 D30
flabel metal2 s 32668 85802 32668 85802 1 FreeSans 480 0 0 160 D31
flabel metal2 s 32762 85812 32762 85812 1 FreeSans 480 0 0 160 D32
flabel metal2 s 32876 85814 32876 85814 1 FreeSans 480 0 0 160 D33
flabel metal2 s 32988 85812 32988 85812 1 FreeSans 480 0 0 160 D34
flabel metal2 s 33086 85818 33086 85818 1 FreeSans 480 0 0 160 D35
flabel metal2 s 33184 85804 33184 85804 1 FreeSans 480 0 0 160 D36
flabel metal2 s 33300 85810 33300 85810 1 FreeSans 480 0 0 160 D37
flabel metal2 s 41126 85804 41126 85804 1 FreeSans 480 0 0 160 VOUT3
flabel metal3 s 104 79440 104 79440 7 FreeSans 480 0 0 160 VSSD
flabel metal3 s 42 80194 42 80194 7 FreeSans 480 0 0 160 VCCD
flabel locali s 60 86 60 86 7 FreeSans 480 0 0 160 VREFH
flabel locali s 40 79054 40 79054 7 FreeSans 480 0 0 160 VREFL
flabel metal3 s 72 77844 72 77844 7 FreeSans 480 0 0 160 VSSA
flabel metal3 s 34 85442 34 85442 7 FreeSans 640 0 0 0 VDDA
flabel metal3 s 26 81682 26 81682 7 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 474 68 474 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 1702 68 1702 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 2930 68 2930 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 4158 68 4158 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 5386 68 5386 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 6614 68 6614 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 7842 68 7842 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 9070 68 9070 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 10298 68 10298 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 11526 68 11526 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 12754 68 12754 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 13982 68 13982 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 15210 68 15210 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 16438 68 16438 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 17666 68 17666 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 18894 68 18894 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 20122 68 20122 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 21350 68 21350 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 22578 68 22578 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 23806 68 23806 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 25034 68 25034 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 26262 68 26262 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 27490 68 27490 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 28718 68 28718 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 29946 68 29946 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 31174 68 31174 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 32402 68 32402 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 33630 68 33630 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 34858 68 34858 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 36086 68 36086 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 37314 68 37314 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 38542 68 38542 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 39770 68 39770 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 40998 68 40998 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 42226 68 42226 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 43454 68 43454 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 44682 68 44682 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 45910 68 45910 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 47138 68 47138 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 48366 68 48366 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 49594 68 49594 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 50822 68 50822 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 52050 68 52050 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 53278 68 53278 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 54506 68 54506 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 55734 68 55734 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 56962 68 56962 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 58190 68 58190 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 59418 68 59418 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 60646 68 60646 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 61874 68 61874 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 63102 68 63102 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 64330 68 64330 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 65558 68 65558 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 66786 68 66786 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 68014 68 68014 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 69242 68 69242 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 70470 68 70470 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 71698 68 71698 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 72926 68 72926 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 74154 68 74154 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 75382 68 75382 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 76610 68 76610 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 68 77838 68 77838 0 FreeSans 640 0 0 0 VSSA
flabel metal3 s 92 1162 92 1162 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 2390 92 2390 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 3618 92 3618 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 4846 92 4846 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 6074 92 6074 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 7302 92 7302 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 8530 92 8530 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 9758 92 9758 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 10986 92 10986 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 12214 92 12214 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 13442 92 13442 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 14670 92 14670 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 15898 92 15898 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 17126 92 17126 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 18354 92 18354 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 19582 92 19582 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 20810 92 20810 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 22038 92 22038 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 23266 92 23266 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 24494 92 24494 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 25722 92 25722 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 26950 92 26950 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 28178 92 28178 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 29406 92 29406 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 30634 92 30634 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 31862 92 31862 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 33090 92 33090 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 34318 92 34318 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 35546 92 35546 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 36774 92 36774 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 38002 92 38002 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 39230 92 39230 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 40458 92 40458 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 41686 92 41686 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 42914 92 42914 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 44142 92 44142 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 45370 92 45370 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 46598 92 46598 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 47826 92 47826 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 49054 92 49054 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 50282 92 50282 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 51510 92 51510 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 52738 92 52738 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 53966 92 53966 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 55194 92 55194 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 56422 92 56422 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 57650 92 57650 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 58878 92 58878 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 60106 92 60106 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 61334 92 61334 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 62562 92 62562 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 63790 92 63790 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 65018 92 65018 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 66246 92 66246 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 67474 92 67474 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 68702 92 68702 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 69930 92 69930 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 71158 92 71158 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 72386 92 72386 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 73614 92 73614 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 74842 92 74842 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 76070 92 76070 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 77298 92 77298 0 FreeSans 640 0 0 0 VDDA
flabel metal3 s 92 78526 92 78526 0 FreeSans 640 0 0 0 VDDA
<< end >>
