* NGSPICE file created from 7_bit_dac_flat.ext - technology: sky130A

.subckt 7_bit_dac D0 VREFL D1 D2 D3 D5 D6 D0_BUF VREFH D1_BUF D2_BUF D3_BUF
+ D5_BUF D6_BUF VOUT D4_BUF D4 VSS VCC
X0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H D0_BUF.t2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t450 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.D3.t2 VSS.t194 VSS.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_32334# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 a_1556_24966# VCC.t307 VCC.t306 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X6 6_bit_dac_0[1].5_bit_dac_1.D3.t0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t606 VSS.t605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.D4.t2 VCC.t597 VCC.t596 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].VOUT VCC.t603 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X9 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_37246# a_544_37677# VCC.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 a_544_32765# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X11 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_29878# a_544_30309# VCC.t317 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t388 VCC.t387 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X13 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t130 VSS.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X14 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_33562# a_544_33993# VCC.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X15 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.VOUT.t0 VCC.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X16 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_7774# VSS.t465 VSS.t464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X17 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t183 VCC.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t364 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X19 switch_n_3v3_1.D5.t1 6_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t552 VCC.t551 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X20 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t142 VCC.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 a_544_11889# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X22 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X23 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X24 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].VOUT VSS.t604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X25 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t385 VCC.t384 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X26 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X27 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 a_1556_5318# VCC.t559 VCC.t558 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X28 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t0 VCC.t139 VCC.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X29 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_2862# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t595 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_20054# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X31 a_544_18029# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X32 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_28650# 6_bit_dac_0[1].5_bit_dac_1.VREFL VSS.t540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X33 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X34 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_32334# VSS.t595 VSS.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X35 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t448 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X36 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X37 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X38 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 VSS.t471 VSS.t470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X39 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_26194# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X40 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_37246# VCC.t337 VCC.t336 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X41 6_bit_dac_0[1].5_bit_dac_1.D0 a_1556_29878# VCC.t316 VCC.t315 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X42 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ D3.t0 VCC.t21 VCC.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X43 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_33562# VCC.t291 VCC.t290 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X44 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_6546# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X45 6_bit_dac_0[1].switch_n_3v3_0.DX_ D5.t0 VCC.t366 VCC.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X46 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_1634# a_544_2065# VCC.t124 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X47 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 VCC.t433 VCC.t432 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X48 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_4090# a_544_4521# VCC.t490 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X49 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X50 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X51 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS.t47 VSS.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X52 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VCC.t623 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X53 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.VREFL VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X54 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 VCC.t284 VCC.t283 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X55 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VREFL.t2 VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X56 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X57 a_544_30309# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X58 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_33562# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X59 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X60 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X61 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t269 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X62 VOUT.t2 D6_BUF.t2 6_bit_dac_0[1].VOUT.t1 VCC.t491 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X63 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X64 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X65 a_544_15573# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X66 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X67 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X68 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t437 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X69 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_36018# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X70 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X71 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_31106# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t577 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X72 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X73 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_9002# VCC.t607 VCC.t606 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X74 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t358 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X75 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X76 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t359 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X77 a_1556_11458# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 VCC.t398 VCC.t397 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X78 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X79 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS.t207 VSS.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X80 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X81 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 VCC.t408 VCC.t407 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X82 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_4090# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X83 a_1556_17598# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t495 VCC.t494 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X84 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 VCC.t526 VCC.t525 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X85 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT D2_BUF.t2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X86 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VCC.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X87 a_544_25397# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X88 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X89 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_7774# a_544_8205# VCC.t464 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X90 6_bit_dac_0[0].5_bit_dac_0.VOUT.t4 6_bit_dac_0[0].5_bit_dac_1.D4.t2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].VOUT VSS.t322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X91 a_544_20485# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X92 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t483 VCC.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X93 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X94 a_544_10661# 6_bit_dac_0[0].5_bit_dac_1.D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X95 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t379 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X96 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t246 VCC.t245 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X97 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_11458# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X98 a_544_26625# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X99 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X100 a_1556_24966# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t260 VSS.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X101 6_bit_dac_0[0].5_bit_dac_1.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t263 VSS.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X102 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X103 a_1556_10230# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t270 VSS.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X104 a_544_11889# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X105 a_1556_22510# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t169 VCC.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X106 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t592 VSS.t591 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X107 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_12686# a_544_13117# VCC.t217 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X108 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t327 VSS.t326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X109 6_bit_dac_0[0].VOUT.t1 D5_BUF.t2 6_bit_dac_0[0].5_bit_dac_0.VOUT.t3 VCC.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X110 6_bit_dac_0[0].5_bit_dac_1.D3.t1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t506 VCC.t505 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X111 a_1556_15142# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t32 VCC.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X112 a_544_18029# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X113 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t341 VCC.t340 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X114 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t147 VSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X115 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t91 VCC.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X116 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X117 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X118 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t97 VCC.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X119 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.D3.t2 VCC.t115 VCC.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X120 6_bit_dac_0[0].5_bit_dac_1.D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t213 VSS.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X121 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_11458# VSS.t177 VSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X122 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t517 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X123 6_bit_dac_0[0].5_bit_dac_1.VOUT D4_BUF.t2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].VOUT VSS.t567 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X124 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X125 6_bit_dac_0[0].VOUT.t0 switch_n_3v3_1.DX_ VOUT.t1 VCC.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X126 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X127 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X128 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t220 VCC.t219 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X129 D3_BUF.t0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t423 VSS.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X130 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS.t192 VSS.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X131 a_544_38905# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X132 a_544_3293# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X133 a_544_31537# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X134 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t405 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X135 a_544_35221# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X136 a_544_29081# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X137 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_12686# VCC.t216 VCC.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X138 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X139 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X140 D4_BUF.t0 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.DX_ VSS.t54 VSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X141 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.VOUT VCC.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X142 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X143 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_29878# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X144 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_1.D3.t2 VSS.t201 VSS.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X145 a_544_5749# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X146 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 VCC.t152 VCC.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X147 switch_n_3v3_1.D5.t0 6_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t556 VSS.t555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X148 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X149 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t245 VSS.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X150 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_15142# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X151 a_544_30309# 6_bit_dac_0[1].5_bit_dac_1.VREFL VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X152 a_1556_20054# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t447 VCC.t446 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X153 a_1556_28650# 6_bit_dac_0[1].5_bit_dac_1.D0 VSS.t461 VSS.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X154 6_bit_dac_0[0].5_bit_dac_1.D4.t0 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.DX_ VSS.t25 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X155 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t620 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X156 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t76 VSS.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X157 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t516 VCC.t515 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X158 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X159 a_544_15573# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X160 a_544_8205# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X161 a_1556_26194# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 VCC.t441 VCC.t440 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X162 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X163 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_12686# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X164 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t79 VCC.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X165 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t11 VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X166 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X167 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X168 a_1556_1634# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 VCC.t566 VCC.t565 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X169 a_1556_6546# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS.t474 VSS.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X170 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X171 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X172 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.VOUT.t1 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X173 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X174 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X175 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X176 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t310 VCC.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X177 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_10230# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t514 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X178 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X179 6_bit_dac_0[1].5_bit_dac_1.D0 a_1556_29878# VSS.t317 VSS.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X180 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t447 VSS.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X181 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_18826# 6_bit_dac_0[1].VREFH VSS.t544 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X182 6_bit_dac_0[1].5_bit_dac_0.VOUT 6_bit_dac_0[1].5_bit_dac_1.D4.t3 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].VOUT VSS.t601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X183 a_1556_4090# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 VCC.t59 VCC.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X184 a_544_33993# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X185 a_544_6977# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X186 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t549 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X187 6_bit_dac_0[1].switch_n_3v3_0.DX_ D5.t1 VSS.t301 VSS.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X188 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t251 VCC.t250 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X189 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_16370# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X190 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 a_1556_15142# VSS.t619 VSS.t618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X191 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t223 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X192 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X193 a_544_36449# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X194 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X195 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X196 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X197 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.DX_ switch_n_3v3_1.D4.t2 VSS.t56 VSS.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X198 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_20054# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X199 a_1556_33562# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 VSS.t114 VSS.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X200 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t634 VSS.t633 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X201 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t630 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X202 6_bit_dac_0[0].5_bit_dac_1.VOUT 6_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].VOUT.t5 VCC.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X203 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_7774# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X204 a_544_9433# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X205 a_544_20485# 6_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X206 a_1556_36018# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS.t350 VSS.t349 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X207 a_1556_31106# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 VCC.t156 VCC.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X208 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_21282# a_544_21713# VCC.t281 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X209 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.D1 VSS.t44 VSS.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X210 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t627 VSS.t626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X211 switch_n_3v3_1.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t106 VCC.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X212 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VCC.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X213 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_5318# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t557 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X214 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.VREFL VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X215 a_544_26625# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X216 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X217 a_1556_4090# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 VSS.t63 VSS.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X218 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t481 VSS.t480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X219 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X220 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_23738# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X221 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X222 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 VCC.t222 VCC.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X223 6_bit_dac_0[1].5_bit_dac_1.VOUT.t1 switch_n_3v3_1.D4.t3 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT VCC.t615 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X224 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X225 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_16370# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X226 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t299 VSS.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X227 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_28650# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t536 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X228 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t625 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X229 6_bit_dac_0[0].D0 a_1556_20054# VSS.t36 VSS.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X230 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X231 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t162 VCC.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X232 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X233 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t585 VSS.t584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X234 6_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t493 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X235 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X236 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X237 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t573 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X238 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_13914# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X239 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t411 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X240 a_1556_7774# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t572 VCC.t571 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X241 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X242 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_21282# VCC.t280 VCC.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X243 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS.t624 VSS.t623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X244 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_38474# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X245 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_31106# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X246 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 VCC.t633 VCC.t632 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X247 a_544_837# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X248 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t233 VSS.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X249 6_bit_dac_0[1].5_bit_dac_1.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t8 VSS.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X250 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t414 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X251 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D1 VSS.t414 VSS.t413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X252 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_36018# a_544_36449# VCC.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X253 6_bit_dac_0[1].5_bit_dac_1.D4.t0 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.DX_ VSS.t22 VSS.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X254 a_544_38905# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X255 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X256 a_544_31537# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X257 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t470 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X258 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t486 VCC.t485 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X259 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS.t70 VSS.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X260 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X261 a_544_35221# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X262 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 VCC.t522 VCC.t521 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X263 6_bit_dac_0[1].VOUT.t4 switch_n_3v3_1.D5.t2 6_bit_dac_0[1].5_bit_dac_0.VOUT VCC.t259 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X264 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_1634# VCC.t123 VCC.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X265 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_6546# VSS.t79 VSS.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X266 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X267 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X268 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X269 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_21282# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X270 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X271 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X272 a_544_14345# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X273 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X274 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.VOUT VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X275 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X276 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_4090# VCC.t489 VCC.t488 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X277 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X278 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_9002# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t605 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X279 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_38474# VSS.t188 VSS.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X280 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t439 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X281 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_27422# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X282 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_31106# VSS.t581 VSS.t580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X283 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X284 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t510 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X285 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t477 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X286 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X287 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_406# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t201 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X288 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ D2.t0 VSS.t235 VSS.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X289 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_2862# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X290 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS.t404 VSS.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X291 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_36018# VCC.t287 VCC.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X292 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.DX_ D4.t0 VSS.t503 VSS.t502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X293 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_24966# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X294 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_5318# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X295 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 VCC.t467 VCC.t466 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X296 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t590 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X297 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X298 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t314 VSS.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X299 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_4090# VSS.t491 VSS.t490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X300 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X301 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X302 a_544_13117# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X303 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.VOUT.t2 VCC.t334 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X304 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X305 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t456 VCC.t455 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X306 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X307 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X308 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X309 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X310 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X311 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_32334# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X312 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X313 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t329 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X314 a_544_19257# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X315 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X316 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_37246# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X317 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X318 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].VOUT VSS.t421 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X319 a_1556_12686# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t506 VSS.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X320 VREFL.t0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X321 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t555 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X322 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_29878# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t314 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X323 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X324 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_7774# VCC.t463 VCC.t462 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X325 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t569 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X326 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_33562# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X327 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X328 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 VSS.t256 VSS.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X329 a_1556_10230# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t268 VCC.t267 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X330 a_1556_18826# 6_bit_dac_0[0].D0 VSS.t407 VSS.t406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X331 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.D4.t3 VSS.t324 VSS.t323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X332 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t564 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X333 a_1556_406# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t630 VSS.t629 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X334 D0_BUF.t1 a_1556_406# VSS.t199 VSS.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X335 a_1556_16370# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 VCC.t357 VCC.t356 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X336 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t92 VSS.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X337 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X338 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VOUT VCC.t386 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X339 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_9002# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t613 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X340 6_bit_dac_0[1].5_bit_dac_1.VOUT.t4 6_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].VOUT.t3 VCC.t550 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X341 6_bit_dac_0[0].5_bit_dac_1.D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t213 VCC.t212 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X342 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X343 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X344 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t275 VSS.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X345 a_544_24169# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X346 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X347 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X348 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D1 VSS.t144 VSS.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X349 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X350 a_544_22941# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X351 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X352 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t543 VCC.t542 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X353 a_544_16801# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X354 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X355 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X356 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X357 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_17598# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X358 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.D1 VCC.t295 VCC.t294 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X359 a_1556_23738# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 VSS.t59 VSS.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X360 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X361 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t550 VSS.t549 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X362 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_13914# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X363 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t503 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X364 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X365 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X366 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t230 VSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X367 a_1556_16370# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS.t362 VSS.t361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X368 a_1556_28650# 6_bit_dac_0[1].5_bit_dac_1.D0 VCC.t460 VCC.t459 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X369 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t348 VCC.t347 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X370 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t133 VSS.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X371 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X372 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t71 VCC.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X373 a_544_14345# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X374 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].D1 VSS.t86 VSS.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X375 6_bit_dac_0[0].5_bit_dac_1.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t262 VCC.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X376 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.D3.t3 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X377 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS.t632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X378 a_1556_13914# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 VCC.t15 VCC.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X379 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t9 VCC.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X380 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.D2 VSS.t265 VSS.t264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X381 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t204 VSS.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X382 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X383 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 VCC.t68 VCC.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X384 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t580 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X385 6_bit_dac_0[1].VOUT.t5 switch_n_3v3_1.D5.t3 6_bit_dac_0[1].5_bit_dac_1.VOUT.t5 VSS.t319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X386 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_17598# VSS.t500 VSS.t499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X387 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t547 VSS.t546 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X388 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t444 VCC.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X389 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].VOUT switch_n_3v3_1.D3.t3 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X390 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X391 a_544_21713# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X392 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X393 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X394 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_13914# VSS.t117 VSS.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X395 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VCC.t610 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X396 D2_BUF.t0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t616 VSS.t615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X397 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t453 VCC.t452 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X398 a_544_37677# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X399 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t417 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X400 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 VSS.t384 VSS.t383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X401 a_544_2065# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X402 a_544_27853# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X403 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X404 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t354 VCC.t353 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X405 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t527 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X406 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t529 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X407 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_23738# a_544_24169# VCC.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X408 a_1556_21282# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS.t379 VSS.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X409 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 VCC.t193 VCC.t192 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X410 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X411 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t236 VCC.t235 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X412 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF.t2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X413 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D1 VSS.t396 VSS.t395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X414 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t524 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X415 a_1556_27422# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t4 VSS.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X416 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS.t73 VSS.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X417 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.D1 VCC.t43 VCC.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X418 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_18826# a_544_19257# VCC.t540 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X419 a_1556_2862# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t174 VSS.t173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X420 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X421 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X422 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t125 VSS.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X423 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t423 VCC.t422 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X424 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t627 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X425 a_544_6977# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X426 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X427 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_11458# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X428 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X429 a_1556_24966# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t257 VCC.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X430 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t520 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X431 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D1 VCC.t416 VCC.t415 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X432 a_1556_5318# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t513 VSS.t512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X433 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X434 a_544_3293# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X435 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X436 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X437 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t587 VCC.t586 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X438 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t104 VSS.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X439 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X440 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t355 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X441 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VOUT VSS.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X442 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_23738# VCC.t226 VCC.t225 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X443 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t481 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X444 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_12686# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X445 a_544_32765# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X446 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X447 a_544_5749# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X448 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 VCC.t532 VCC.t531 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X449 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t243 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X450 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t149 VCC.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X451 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X452 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X453 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t458 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X454 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X455 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_26194# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X456 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_406# a_544_837# VCC.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X457 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t375 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X458 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_18826# VCC.t539 VCC.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X459 a_1556_32334# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t375 VSS.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X460 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_22510# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t589 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X461 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS.t101 VSS.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X462 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_1.D2 VCC.t109 VCC.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X463 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X464 D3_BUF.t1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t420 VCC.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X465 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT VCC.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X466 switch_n_3v3_1.D3.t0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t609 VSS.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X467 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_6546# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X468 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_27422# a_544_27853# VCC.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X469 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X470 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_1634# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t121 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X471 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].VOUT VCC.t504 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X472 a_1556_37246# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t186 VCC.t185 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X473 a_1556_29878# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t39 VCC.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X474 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t351 VCC.t350 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X475 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X476 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X477 a_544_22941# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X478 a_1556_33562# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 VCC.t112 VCC.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X479 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t169 VSS.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X480 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_1.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X481 a_544_4521# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X482 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L D0_BUF.t3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X483 D1_BUF.t0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t371 VSS.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X484 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_4090# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t487 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X485 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X486 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_29878# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X487 6_bit_dac_0[1].5_bit_dac_0.VOUT 6_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].VOUT.t2 VSS.t554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X488 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].VOUT D3_BUF.t2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X489 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X490 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t334 VSS.t333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X491 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X492 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X493 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t378 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X494 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].VOUT VSS.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X495 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t242 VCC.t241 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X496 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X497 VOUT.t3 D6_BUF.t3 6_bit_dac_0[0].VOUT.t3 VSS.t485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X498 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_26194# VSS.t28 VSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X499 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X500 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_15142# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X501 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t391 VCC.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X502 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X503 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X504 6_bit_dac_0[1].5_bit_dac_1.D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t159 VCC.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X505 a_1556_9002# 6_bit_dac_0[0].5_bit_dac_1.D0 VSS.t135 VSS.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X506 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t480 VCC.t479 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X507 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_22510# VSS.t588 VSS.t587 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X508 a_544_837# D0_BUF.t4 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X509 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t474 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X510 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X511 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 VSS.t304 VSS.t303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X512 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_34790# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t433 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X513 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_27422# VCC.t325 VCC.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X514 a_544_9433# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X515 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.D3.t3 VCC.t196 VCC.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X516 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_37246# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X517 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_32334# a_544_32765# VCC.t591 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X518 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t390 VSS.t389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X519 6_bit_dac_0[1].5_bit_dac_1.D3.t1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t600 VCC.t599 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X520 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_4090# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS.t489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X521 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t180 VSS.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X522 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_2862# VSS.t599 VSS.t598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X523 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_34790# a_544_35221# VCC.t430 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X524 a_544_37677# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X525 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_38474# a_544_38905# VCC.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X526 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t129 VCC.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X527 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t431 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X528 6_bit_dac_0[1].5_bit_dac_1.D4.t1 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.DX_ VCC.t19 VCC.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X529 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t164 VCC.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X530 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 a_1556_5318# VSS.t562 VSS.t561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X531 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t233 VCC.t232 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X532 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X533 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VOUT VSS.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X534 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D1 VCC.t410 VCC.t409 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X535 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t404 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X536 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_20054# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X537 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X538 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 a_1556_34790# VSS.t432 VSS.t431 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X539 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t472 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X540 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_7774# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t461 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X541 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X542 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t255 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X543 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_37246# VSS.t342 VSS.t341 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X544 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_32334# VCC.t590 VCC.t589 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X545 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X546 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_21282# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X547 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X548 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ D3.t1 VSS.t14 VSS.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X549 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 VCC.t469 VCC.t468 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X550 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_1634# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X551 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 a_1556_34790# VCC.t429 VCC.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X552 a_544_837# VREFH.t0 VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X553 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_38474# VCC.t190 VCC.t189 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X554 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_6546# a_544_6977# VCC.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X555 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X556 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.DX_ D4.t1 VCC.t368 VCC.t367 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X557 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ D2.t1 VCC.t11 VCC.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X558 D6_BUF.t0 switch_n_3v3_1.DX_ VSS.t89 VSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X559 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X560 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X561 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X562 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VCC.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X563 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 VCC.t46 VCC.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X564 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS.t285 VSS.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X565 a_544_25397# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X566 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X567 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X568 a_544_11889# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X569 6_bit_dac_0[1].VOUT.t0 switch_n_3v3_1.DX_ VOUT.t0 VSS.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X570 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D1 VCC.t145 VCC.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X571 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X572 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_38474# VREFL.t1 VSS.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X573 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X574 a_544_10661# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X575 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X576 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t439 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X577 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X578 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X579 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_31106# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X580 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X581 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_9002# VSS.t612 VSS.t611 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X582 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X583 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_36018# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X584 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X585 a_1556_11458# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS.t400 VSS.t399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X586 switch_n_3v3_1.DX_ D6.t0 VSS.t250 VSS.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X587 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X588 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS.t410 VSS.t409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X589 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 VCC.t207 VCC.t206 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X590 6_bit_dac_0[0].5_bit_dac_1.VREFL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t570 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X591 a_1556_12686# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t502 VCC.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X592 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF.t3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X593 6_bit_dac_0[1].5_bit_dac_1.VOUT.t0 switch_n_3v3_1.D4.t4 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].VOUT VSS.t621 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X594 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t553 VSS.t552 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X595 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X596 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VCC.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X597 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_2862# a_544_3293# VCC.t594 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X598 6_bit_dac_0[0].VOUT.t2 D5_BUF.t3 6_bit_dac_0[0].5_bit_dac_1.VOUT VSS.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X599 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t484 VSS.t483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X600 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t293 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X601 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t88 VCC.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X602 a_544_30309# 6_bit_dac_0[1].5_bit_dac_1.D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X603 a_544_29081# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X604 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X605 a_544_15573# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X606 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X607 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t312 VCC.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X608 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X609 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X610 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_11458# a_544_11889# VCC.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X611 a_1556_29878# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t40 VSS.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X612 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t524 VSS.t523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X613 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS.t365 VSS.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X614 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X615 a_1556_15142# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t32 VSS.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X616 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_17598# a_544_18029# VCC.t499 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X617 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.VOUT VSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X618 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t345 VSS.t344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X619 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X620 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t322 VCC.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X621 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t94 VSS.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X622 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t546 VCC.t545 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X623 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t265 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X624 6_bit_dac_0[1].5_bit_dac_1.D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t157 VSS.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X625 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 VCC.t254 VCC.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X626 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X627 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t220 VSS.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X628 a_544_33993# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X629 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X630 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_11458# VCC.t179 VCC.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X631 a_544_20485# 6_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X632 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t210 VSS.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X633 a_544_36449# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X634 a_544_8205# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X635 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X636 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_24966# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X637 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_17598# VCC.t498 VCC.t497 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X638 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X639 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X640 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X641 switch_n_3v3_1.D4.t0 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.DX_ VSS.t339 VSS.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X642 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X643 D4_BUF.t1 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.DX_ VCC.t51 VCC.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X644 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_1.D3.t4 VCC.t273 VCC.t272 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X645 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X646 a_1556_20054# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t450 VSS.t449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X647 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_10230# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t518 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X648 a_544_25397# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X649 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_22510# a_544_22941# VCC.t584 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X650 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t162 VSS.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X651 switch_n_3v3_1.D3.t1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t602 VCC.t601 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X652 D5_BUF.t0 6_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t566 VSS.t565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X653 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t631 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X654 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_15142# a_544_15573# VCC.t614 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X655 6_bit_dac_0[0].5_bit_dac_1.VOUT D4_BUF.t3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT VCC.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X656 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X657 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.VOUT.t3 VSS.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X658 6_bit_dac_0[0].5_bit_dac_1.D4.t1 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.DX_ VCC.t23 VCC.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X659 a_544_3293# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X660 a_544_10661# 6_bit_dac_0[0].5_bit_dac_1.VREFL VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X661 a_1556_21282# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 VCC.t377 VCC.t376 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X662 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t82 VSS.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X663 a_1556_1634# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS.t569 VSS.t568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X664 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_17598# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X665 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X666 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X667 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X668 6_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t478 VSS.t477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X669 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X670 a_544_5749# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X671 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t311 VSS.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X672 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X673 6_bit_dac_0[0].5_bit_dac_0.VOUT.t5 6_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].VOUT.t4 VSS.t564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X674 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X675 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X676 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X677 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X678 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_13914# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X679 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X680 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 a_1556_24966# VSS.t307 VSS.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X681 a_1556_6546# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 VCC.t473 VCC.t472 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X682 a_544_2065# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X683 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.D4.t4 VSS.t603 VSS.t602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X684 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t253 VSS.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X685 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X686 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_22510# VCC.t583 VCC.t582 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X687 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t126 VCC.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X688 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t541 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X689 6_bit_dac_0[0].5_bit_dac_1.D0 a_1556_10230# VSS.t517 VSS.t516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X690 a_544_38905# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X691 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X692 a_544_31537# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X693 6_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_1.D5.t4 VSS.t321 VSS.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X694 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X695 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 VCC.t301 VCC.t300 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X696 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 a_1556_15142# VCC.t613 VCC.t612 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X697 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X698 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t436 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X699 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.DX_ switch_n_3v3_1.D4.t5 VCC.t617 VCC.t616 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X700 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t533 VSS.t532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X701 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X702 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_20054# a_544_20485# VCC.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X703 a_1556_38474# D0.t0 VSS.t336 VSS.t335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X704 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_28650# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X705 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_2862# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X706 a_544_4521# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X707 a_1556_31106# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS.t153 VSS.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X708 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t417 VSS.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X709 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t66 VSS.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X710 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t629 VCC.t628 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X711 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_5318# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X712 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VCC.t260 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X713 a_1556_36018# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 VCC.t344 VCC.t343 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X714 a_544_29081# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X715 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_26194# a_544_26625# VCC.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X716 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X717 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X718 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t299 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X719 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t622 VCC.t621 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X720 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS.t222 VSS.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X721 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 VCC.t99 VCC.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X722 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X723 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t574 VSS.t573 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X724 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X725 6_bit_dac_0[1].5_bit_dac_1.VREFL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X726 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS.t415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X727 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X728 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t160 VSS.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X729 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X730 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_23738# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t224 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X731 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t559 VSS.t558 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X732 a_544_9433# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t577 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X733 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t500 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X734 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X735 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t297 VCC.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X736 6_bit_dac_0[0].D0 a_1556_20054# VCC.t34 VCC.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X737 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X738 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X739 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_28650# VSS.t538 VSS.t537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X740 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t579 VCC.t578 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X741 a_1556_2862# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t175 VCC.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X742 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X743 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X744 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_18826# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t537 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X745 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X746 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.D2 VSS.t368 VSS.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X747 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t557 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X748 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_33562# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X749 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_26194# VCC.t26 VCC.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X750 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t140 VSS.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X751 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 VCC.t619 VCC.t618 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X752 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X753 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_36018# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X754 a_544_33993# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X755 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_31106# a_544_31537# VCC.t576 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X756 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t1 VSS.t127 VSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X757 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t487 VSS.t486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X758 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X759 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.D3.t4 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t197 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X760 6_bit_dac_0[1].5_bit_dac_1.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t5 VCC.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X761 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS.t526 VSS.t525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X762 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_1634# VSS.t121 VSS.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X763 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t386 VSS.t385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X764 a_544_13117# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X765 a_544_36449# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X766 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X767 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X768 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X769 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t421 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X770 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 VCC.t65 VCC.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X771 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X772 6_bit_dac_0[1].5_bit_dac_0.VOUT 6_bit_dac_0[1].5_bit_dac_1.D4.t5 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VOUT VCC.t271 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X773 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_6546# VCC.t75 VCC.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X774 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t465 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X775 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_26194# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X776 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_9002# 6_bit_dac_0[0].5_bit_dac_1.VREFL VSS.t610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X777 a_544_19257# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X778 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X779 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_33562# VSS.t291 VSS.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X780 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_22510# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t586 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X781 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X782 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t626 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X783 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_406# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X784 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t548 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X785 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 VSS.t436 VSS.t435 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X786 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_27422# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t323 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X787 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X788 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_36018# VSS.t287 VSS.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X789 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_31106# VCC.t575 VCC.t574 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X790 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X791 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t173 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X792 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS.t467 VSS.t466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X793 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_7774# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X794 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 VCC.t400 VCC.t399 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X795 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_5318# a_544_5749# VCC.t556 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X796 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X797 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X798 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.D3.t4 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X799 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t248 VSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X800 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT VCC.t349 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X801 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X802 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t456 VSS.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X803 a_544_24169# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X804 a_544_18029# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X805 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_34790# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X806 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X807 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X808 D6_BUF.t1 switch_n_3v3_1.DX_ VCC.t84 VCC.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X809 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X810 a_544_16801# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X811 a_544_14345# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X812 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X813 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t342 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X814 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X815 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t389 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X816 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_37246# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X817 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_32334# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t588 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X818 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t457 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X819 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X820 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X821 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X822 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X823 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X824 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_2862# VCC.t593 VCC.t592 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X825 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X826 a_1556_17598# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t495 VSS.t494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X827 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_34790# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t427 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X828 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT VSS.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X829 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.D3.t5 VSS.t282 VSS.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X830 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_38474# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t188 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X831 a_1556_13914# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 VSS.t18 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X832 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X833 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t471 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X834 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.D4.t4 VCC.t93 VCC.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X835 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].VOUT D3_BUF.t3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X836 a_1556_406# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t625 VCC.t624 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X837 D0_BUF.t0 a_1556_406# VCC.t199 VCC.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X838 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].VOUT VCC.t598 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X839 switch_n_3v3_1.DX_ D6.t1 VCC.t248 VCC.t247 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X840 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_9002# a_544_9433# VCC.t604 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X841 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t454 VSS.t453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X842 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.VOUT VCC.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X843 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X844 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X845 a_544_21713# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X846 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t548 VCC.t547 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X847 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t361 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X848 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X849 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X850 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.D1 VSS.t295 VSS.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X851 a_544_27853# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X852 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_12686# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X853 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X854 6_bit_dac_0[0].5_bit_dac_1.D3.t0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t510 VSS.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X855 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X856 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X857 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_10230# a_544_10661# VCC.t513 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X858 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t492 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X859 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_18826# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t543 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X860 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X861 a_544_13117# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X862 a_1556_23738# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 VCC.t54 VCC.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X863 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t346 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X864 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t352 VSS.t351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X865 D5_BUF.t1 6_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t561 VCC.t560 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X866 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t426 VSS.t425 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X867 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D1 VSS.t419 VSS.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X868 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].VOUT VSS.t508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X869 a_544_19257# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X870 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_16370# a_544_16801# VCC.t239 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X871 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS.t531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X872 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X873 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t132 VCC.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X874 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 VSS.t529 VSS.t528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X875 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X876 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t48 VCC.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X877 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_1.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X878 a_1556_18826# 6_bit_dac_0[0].D0 VCC.t403 VCC.t402 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X879 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 VCC.t360 VCC.t359 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X880 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS.t424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X881 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t203 VCC.t202 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X882 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.D2 VCC.t264 VCC.t263 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X883 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_12686# VSS.t215 VSS.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X884 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t454 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X885 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 VSS.t149 VSS.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X886 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X887 a_544_32765# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X888 6_bit_dac_0[0].5_bit_dac_1.D0 a_1556_10230# VCC.t512 VCC.t511 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X889 a_544_26625# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X890 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_18826# VSS.t542 VSS.t541 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X891 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X892 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t358 VSS.t357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X893 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VCC.t352 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X894 a_544_22941# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X895 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t276 VCC.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X896 D2_BUF.t1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t609 VCC.t608 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X897 6_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_1.D5.t5 VCC.t319 VCC.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X898 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t551 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X899 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_1.D2 VSS.t109 VSS.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X900 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X901 a_544_6977# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X902 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_23738# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X903 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_16370# VCC.t238 VCC.t237 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X904 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X905 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t438 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X906 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t237 VSS.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X907 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t528 VCC.t527 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X908 a_1556_26194# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS.t442 VSS.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X909 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X910 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 VCC.t425 VCC.t424 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X911 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_16370# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X912 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_28650# a_544_29081# VCC.t535 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X913 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT D2_BUF.t3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t302 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X914 a_544_24169# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X915 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t50 VSS.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X916 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t413 VCC.t412 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X917 a_1556_22510# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t165 VSS.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X918 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D1 VCC.t393 VCC.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X919 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].VOUT switch_n_3v3_1.D3.t5 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X920 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_13914# a_544_14345# VCC.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X921 a_544_16801# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X922 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X923 a_1556_27422# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t1 VCC.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X924 a_544_2065# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X925 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X926 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X927 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t229 VCC.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X928 6_bit_dac_0[0].5_bit_dac_0.VOUT.t2 6_bit_dac_0[0].5_bit_dac_1.D4.t5 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VOUT VCC.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X929 a_1556_7774# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t576 VSS.t575 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X930 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X931 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X932 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.D3.t5 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X933 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].D1 VCC.t81 VCC.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X934 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t509 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X935 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t585 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X936 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_11458# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X937 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X938 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t519 VCC.t518 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X939 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X940 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_23738# VSS.t225 VSS.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X941 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t98 VSS.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X942 a_1556_5318# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t508 VCC.t507 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X943 a_544_8205# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X944 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X945 a_544_35221# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X946 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X947 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t102 VCC.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X948 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 VSS.t535 VSS.t534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X949 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_17598# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t496 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X950 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_16370# VSS.t240 VSS.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X951 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_28650# VCC.t534 VCC.t533 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X952 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X953 6_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t476 VCC.t475 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X954 a_544_37677# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t347 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X955 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS.t428 VSS.t427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X956 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X957 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X958 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X959 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.D2 VCC.t363 VCC.t362 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X960 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_406# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X961 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X962 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_21282# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X963 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_13914# VCC.t118 VCC.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X964 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X965 a_1556_34790# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t438 VSS.t437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X966 switch_n_3v3_1.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t107 VSS.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X967 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].VOUT VCC.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X968 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 VCC.t381 VCC.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X969 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t184 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X970 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_27422# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X971 a_544_21713# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X972 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_1634# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X973 a_1556_37246# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t183 VSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X974 a_1556_32334# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t373 VCC.t372 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X975 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t356 VSS.t355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X976 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t209 VCC.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X977 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t520 VSS.t519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X978 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VOUT VCC.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X979 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X980 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X981 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_6546# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X982 a_1556_34790# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t435 VCC.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X983 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X984 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.D0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X985 a_544_27853# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X986 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X987 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_24966# a_544_25397# VCC.t304 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X988 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_24966# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X989 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X990 a_1556_38474# D0.t1 VCC.t331 VCC.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X991 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t171 VCC.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X992 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t530 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X993 switch_n_3v3_1.D4.t1 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.DX_ VCC.t333 VCC.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X994 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t62 VCC.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X995 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH D0_BUF.t5 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t449 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X996 D1_BUF.t1 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t370 VCC.t369 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X997 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X998 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t51 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X999 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1000 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_10230# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1001 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t392 VSS.t391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1002 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t328 VCC.t327 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1003 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT VSS.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1004 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_22510# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t581 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1005 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_21282# VSS.t277 VSS.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1006 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS.t636 VSS.t635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1007 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].VOUT 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t434 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1008 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_15142# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t611 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1009 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t383 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1010 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t554 VCC.t553 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1011 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t563 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1012 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_27422# VSS.t329 VSS.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1013 a_1556_9002# 6_bit_dac_0[0].5_bit_dac_1.D0 VCC.t135 VCC.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1014 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t568 VCC.t567 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1015 a_544_4521# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
R0 VSS.n18877 VSS.n40 106073
R1 VSS.n1019 VSS.n40 54262.5
R2 VSS.n18877 VSS.n24 12274.8
R3 VSS.n18877 VSS.n25 12232.2
R4 VSS.n18877 VSS.n23 12232.2
R5 VSS.n18877 VSS.n32 12232.2
R6 VSS.n18877 VSS.n22 12232.2
R7 VSS.n18877 VSS.n26 12232.2
R8 VSS.n18877 VSS.n21 12232.2
R9 VSS.n18877 VSS.n27 12232.2
R10 VSS.n18877 VSS.n20 12232.2
R11 VSS.n18877 VSS.n28 12232.2
R12 VSS.n18877 VSS.n19 12232.2
R13 VSS.n18877 VSS.n29 12232.2
R14 VSS.n18878 VSS.n18877 12232.2
R15 VSS.n18877 VSS.n30 12232.2
R16 VSS.n18877 VSS.n18 12232.2
R17 VSS.n18877 VSS.n31 12232.2
R18 VSS.n18877 VSS.n17 12232.2
R19 VSS.n18877 VSS.n16 12232.2
R20 VSS.n18877 VSS.n33 12232.2
R21 VSS.n18877 VSS.n15 12232.2
R22 VSS.n18877 VSS.n34 12232.2
R23 VSS.n18877 VSS.n14 12232.2
R24 VSS.n18877 VSS.n35 12232.2
R25 VSS.n18877 VSS.n13 12232.2
R26 VSS.n18877 VSS.n36 12232.2
R27 VSS.n18877 VSS.n12 12232.2
R28 VSS.n18877 VSS.n37 12232.2
R29 VSS.n18877 VSS.n11 12232.2
R30 VSS.n18877 VSS.n38 12232.2
R31 VSS.n18877 VSS.n39 12232.2
R32 VSS.n18877 VSS.n10 12232.2
R33 VSS.n18877 VSS.n18876 12232.2
R34 VSS.n1020 VSS.n1019 6909.46
R35 VSS.n18072 VSS.n1020 6909.46
R36 VSS.n18072 VSS.n18071 6909.46
R37 VSS.n18071 VSS.n18070 6909.46
R38 VSS.n18070 VSS.n18069 6909.46
R39 VSS.n18069 VSS.n18068 6909.46
R40 VSS.n18068 VSS.n18067 6909.46
R41 VSS.n18067 VSS.n18066 6909.46
R42 VSS.n18066 VSS.n18065 6909.46
R43 VSS.n18065 VSS.n18064 6909.46
R44 VSS.n18064 VSS.n18063 6909.46
R45 VSS.n18063 VSS.n18062 6909.46
R46 VSS.n18062 VSS.n18061 6909.46
R47 VSS.n18061 VSS.n18060 6909.46
R48 VSS.n18060 VSS.n18059 6909.46
R49 VSS.n18059 VSS.n18058 6909.46
R50 VSS.n18058 VSS.n18057 6909.46
R51 VSS.n18057 VSS.n18056 6909.46
R52 VSS.n18056 VSS.n18055 6909.46
R53 VSS.n18055 VSS.n18054 6909.46
R54 VSS.n18054 VSS.n18053 6909.46
R55 VSS.n18053 VSS.n18052 6909.46
R56 VSS.n18052 VSS.n18051 6909.46
R57 VSS.n18051 VSS.n18050 6909.46
R58 VSS.n18050 VSS.n18049 6909.46
R59 VSS.n18049 VSS.n18048 6909.46
R60 VSS.n18048 VSS.n18047 6909.46
R61 VSS.n18047 VSS.n18046 6909.46
R62 VSS.n18046 VSS.n18045 6909.46
R63 VSS.n18045 VSS.t614 6273.77
R64 VSS.n15981 VSS.n15980 6000
R65 VSS.n15979 VSS.n15978 5972.41
R66 VSS.n17126 VSS.t570 4305.17
R67 VSS.n17718 VSS.t628 4305.17
R68 VSS.n9768 VSS.t405 4305.17
R69 VSS.n16711 VSS.t172 4305.17
R70 VSS.n16118 VSS.t61 4305.17
R71 VSS.n2303 VSS.t514 4305.17
R72 VSS.n3259 VSS.t475 4305.17
R73 VSS.n3851 VSS.t577 4305.17
R74 VSS.n4443 VSS.t137 4305.17
R75 VSS.n5035 VSS.t268 4305.17
R76 VSS.n5268 VSS.t401 4305.17
R77 VSS.n5841 VSS.t504 4305.17
R78 VSS.n6433 VSS.t19 4305.17
R79 VSS.n7992 VSS.t33 4305.17
R80 VSS.n8584 VSS.t360 4305.17
R81 VSS.n9176 VSS.t497 4305.17
R82 VSS.n10360 VSS.t451 4305.17
R83 VSS.n10952 VSS.t377 4305.17
R84 VSS.n11544 VSS.t167 4305.17
R85 VSS.n12136 VSS.t60 4305.17
R86 VSS.n12728 VSS.t257 4305.17
R87 VSS.n13320 VSS.t444 4305.17
R88 VSS.n13912 VSS.t5 4305.17
R89 VSS.n14504 VSS.t459 4305.17
R90 VSS.n15096 VSS.t38 4305.17
R91 VSS.n15688 VSS.t154 4305.17
R92 VSS.n15921 VSS.t376 4305.17
R93 VSS.n7400 VSS.t111 4305.17
R94 VSS.n18712 VSS.t347 4305.17
R95 VSS.n18538 VSS.t440 4305.17
R96 VSS.n835 VSS.t184 4305.17
R97 VSS.n17998 VSS.n1154 3531.03
R98 VSS.n15992 VSS.n1154 3531.03
R99 VSS.n15992 VSS.n15991 3531.03
R100 VSS.n15991 VSS.n15990 3531.03
R101 VSS.n15990 VSS.n15989 3531.03
R102 VSS.n15989 VSS.n15988 3531.03
R103 VSS.n15988 VSS.n15987 3531.03
R104 VSS.n15987 VSS.n15986 3531.03
R105 VSS.n15986 VSS.n15985 3531.03
R106 VSS.n15985 VSS.n15984 3531.03
R107 VSS.n15984 VSS.n15983 3531.03
R108 VSS.n15983 VSS.n15982 3531.03
R109 VSS.n15982 VSS.n15981 3531.03
R110 VSS.n15978 VSS.n15977 3531.03
R111 VSS.n15977 VSS.n15976 3531.03
R112 VSS.n15976 VSS.n15975 3531.03
R113 VSS.n15975 VSS.n15974 3531.03
R114 VSS.n15974 VSS.n15973 3531.03
R115 VSS.n15973 VSS.n15972 3531.03
R116 VSS.n15972 VSS.n15971 3531.03
R117 VSS.n15971 VSS.n15970 3531.03
R118 VSS.n15970 VSS.n15969 3531.03
R119 VSS.n15969 VSS.n15968 3531.03
R120 VSS.n15968 VSS.n207 3531.03
R121 VSS.n18586 VSS.n40 3531.03
R122 VSS.n18586 VSS.n18585 3531.03
R123 VSS.n18585 VSS.n207 3531.03
R124 VSS.n17998 VSS.n17997 3531.03
R125 VSS.t9 VSS.n1154 3054.19
R126 VSS.n15992 VSS.t346 3054.19
R127 VSS.n15991 VSS.t131 3054.19
R128 VSS.n15990 VSS.t590 3054.19
R129 VSS.n15989 VSS.t309 3054.19
R130 VSS.n15988 VSS.t211 3054.19
R131 VSS.n15987 VSS.t551 3054.19
R132 VSS.n15986 VSS.t90 3054.19
R133 VSS.n15985 VSS.t452 3054.19
R134 VSS.n15984 VSS.t218 3054.19
R135 VSS.n15983 VSS.t545 3054.19
R136 VSS.n15982 VSS.t482 3054.19
R137 VSS.n15981 VSS.t273 3054.19
R138 VSS.n15978 VSS.t123 3054.19
R139 VSS.n15977 VSS.t96 3054.19
R140 VSS.n15976 VSS.t202 3054.19
R141 VSS.n15975 VSS.t145 3054.19
R142 VSS.n15974 VSS.t251 3054.19
R143 VSS.n15973 VSS.t102 3054.19
R144 VSS.n15972 VSS.t445 3054.19
R145 VSS.n15971 VSS.t155 3054.19
R146 VSS.n15970 VSS.t158 3054.19
R147 VSS.n15969 VSS.t332 3054.19
R148 VSS.n15968 VSS.t479 3054.19
R149 VSS.t557 VSS.n207 3054.19
R150 VSS.n18586 VSS.t393 3054.19
R151 VSS.n18585 VSS.t297 3054.19
R152 VSS.t572 VSS.n40 3054.19
R153 VSS.n17998 VSS.t522 3054.19
R154 VSS.n17949 VSS.t493 2804.58
R155 VSS.n17948 VSS.t394 2770.93
R156 VSS.n17950 VSS.n17949 2671.38
R157 VSS.t394 VSS.t197 2603.46
R158 VSS.n15978 VSS.n6484 2588.91
R159 VSS.n18585 VSS.n208 2588.02
R160 VSS.n16586 VSS.n1154 2588.02
R161 VSS.n15993 VSS.n15992 2588.02
R162 VSS.n15991 VSS.n1758 2588.02
R163 VSS.n15990 VSS.n2350 2588.02
R164 VSS.n15989 VSS.n2351 2588.02
R165 VSS.n15988 VSS.n2352 2588.02
R166 VSS.n15987 VSS.n2353 2588.02
R167 VSS.n15986 VSS.n2354 2588.02
R168 VSS.n15985 VSS.n5315 2588.02
R169 VSS.n15984 VSS.n5888 2588.02
R170 VSS.n15983 VSS.n6480 2588.02
R171 VSS.n15982 VSS.n6481 2588.02
R172 VSS.n15981 VSS.n6482 2588.02
R173 VSS.n15977 VSS.n6485 2588.02
R174 VSS.n15976 VSS.n6486 2588.02
R175 VSS.n15975 VSS.n6487 2588.02
R176 VSS.n15974 VSS.n6488 2588.02
R177 VSS.n15973 VSS.n6489 2588.02
R178 VSS.n15972 VSS.n6490 2588.02
R179 VSS.n15971 VSS.n6491 2588.02
R180 VSS.n15970 VSS.n6492 2588.02
R181 VSS.n15969 VSS.n6493 2588.02
R182 VSS.n15968 VSS.n6494 2588.02
R183 VSS.n7275 VSS.n207 2588.02
R184 VSS.n18587 VSS.n18586 2588.02
R185 VSS.n973 VSS.n40 2588.02
R186 VSS.n17999 VSS.n17998 2588.02
R187 VSS.n17127 VSS.n17126 2406.66
R188 VSS.n17719 VSS.n17718 2406.66
R189 VSS.n9769 VSS.n9768 2406.66
R190 VSS.n16712 VSS.n16711 2406.66
R191 VSS.n16119 VSS.n16118 2406.66
R192 VSS.n2304 VSS.n2303 2406.66
R193 VSS.n3260 VSS.n3259 2406.66
R194 VSS.n3852 VSS.n3851 2406.66
R195 VSS.n4444 VSS.n4443 2406.66
R196 VSS.n5036 VSS.n5035 2406.66
R197 VSS.n5269 VSS.n5268 2406.66
R198 VSS.n5842 VSS.n5841 2406.66
R199 VSS.n6434 VSS.n6433 2406.66
R200 VSS.n7993 VSS.n7992 2406.66
R201 VSS.n8585 VSS.n8584 2406.66
R202 VSS.n9177 VSS.n9176 2406.66
R203 VSS.n10361 VSS.n10360 2406.66
R204 VSS.n10953 VSS.n10952 2406.66
R205 VSS.n11545 VSS.n11544 2406.66
R206 VSS.n12137 VSS.n12136 2406.66
R207 VSS.n12729 VSS.n12728 2406.66
R208 VSS.n13321 VSS.n13320 2406.66
R209 VSS.n13913 VSS.n13912 2406.66
R210 VSS.n14505 VSS.n14504 2406.66
R211 VSS.n15097 VSS.n15096 2406.66
R212 VSS.n15689 VSS.n15688 2406.66
R213 VSS.n15922 VSS.n15921 2406.66
R214 VSS.n7401 VSS.n7400 2406.66
R215 VSS.n18713 VSS.n18712 2406.66
R216 VSS.n18539 VSS.n18538 2406.66
R217 VSS.n836 VSS.n835 2406.66
R218 VSS.t15 VSS.n17995 2349.66
R219 VSS.t372 VSS.t15 2304.76
R220 VSS.n17001 VSS.t45 1937.11
R221 VSS.n17415 VSS.t583 1937.11
R222 VSS.n9465 VSS.t84 1937.11
R223 VSS.n16407 VSS.t246 1937.11
R224 VSS.t142 VSS.n1757 1937.11
R225 VSS.t457 VSS.n2349 1937.11
R226 VSS.n2956 VSS.t283 1937.11
R227 VSS.n3548 VSS.t312 1937.11
R228 VSS.n4140 VSS.t296 1937.11
R229 VSS.n4732 VSS.t74 1937.11
R230 VSS.t366 VSS.n5314 1937.11
R231 VSS.t548 VSS.n5887 1937.11
R232 VSS.t420 VSS.n6479 1937.11
R233 VSS.n7689 VSS.t83 1937.11
R234 VSS.n8281 VSS.t71 1937.11
R235 VSS.n8873 VSS.t95 1937.11
R236 VSS.n10057 VSS.t67 1937.11
R237 VSS.n10649 VSS.t99 1937.11
R238 VSS.n11241 VSS.t521 1937.11
R239 VSS.n11833 VSS.t397 1937.11
R240 VSS.n12425 VSS.t243 1937.11
R241 VSS.n13017 VSS.t223 1937.11
R242 VSS.n13609 VSS.t170 1937.11
R243 VSS.n14201 VSS.t42 1937.11
R244 VSS.n14793 VSS.t163 1937.11
R245 VSS.n15385 VSS.t527 1937.11
R246 VSS.t181 VSS.n15967 1937.11
R247 VSS.n7096 VSS.t412 1937.11
R248 VSS.t68 VSS.n206 1937.11
R249 VSS.t387 VSS.n18584 1937.11
R250 VSS.n560 VSS.t128 1937.11
R251 VSS.n10138 VSS.t110 1933.6
R252 VSS.n18073 VSS.t434 1930.89
R253 VSS.n16482 VSS.t411 1930.89
R254 VSS.n1647 VSS.t567 1930.89
R255 VSS.n1838 VSS.t530 1930.89
R256 VSS.n3037 VSS.t254 1930.89
R257 VSS.n3629 VSS.t205 1930.89
R258 VSS.n4221 VSS.t271 1930.89
R259 VSS.n4813 VSS.t266 1930.89
R260 VSS.n2434 VSS.t280 1930.89
R261 VSS.n5395 VSS.t190 1930.89
R262 VSS.n5968 VSS.t322 1930.89
R263 VSS.n7770 VSS.t382 1930.89
R264 VSS.n8362 VSS.t150 1930.89
R265 VSS.n8954 VSS.t429 1930.89
R266 VSS.n10730 VSS.t272 1930.89
R267 VSS.n11322 VSS.t637 1930.89
R268 VSS.n11914 VSS.t621 1930.89
R269 VSS.n12506 VSS.t536 1930.89
R270 VSS.n13098 VSS.t302 1930.89
R271 VSS.n13690 VSS.t622 1930.89
R272 VSS.n14282 VSS.t319 1930.89
R273 VSS.n14874 VSS.t369 1930.89
R274 VSS.n15466 VSS.t195 1930.89
R275 VSS.n6574 VSS.t402 1930.89
R276 VSS.n7171 VSS.t601 1930.89
R277 VSS.t469 VSS.n453 1930.89
R278 VSS.t468 VSS.n1018 1930.89
R279 VSS.t141 VSS.n18044 1930.89
R280 VSS.n9546 VSS.t485 1928.19
R281 VSS.n17126 VSS.n17125 1896.55
R282 VSS.n17718 VSS.n17717 1896.55
R283 VSS.n9768 VSS.n9767 1896.55
R284 VSS.n16711 VSS.n16710 1896.55
R285 VSS.n16118 VSS.n16117 1896.55
R286 VSS.n2303 VSS.n2302 1896.55
R287 VSS.n3259 VSS.n3258 1896.55
R288 VSS.n3851 VSS.n3850 1896.55
R289 VSS.n4443 VSS.n4442 1896.55
R290 VSS.n5035 VSS.n5034 1896.55
R291 VSS.n5268 VSS.n5267 1896.55
R292 VSS.n5841 VSS.n5840 1896.55
R293 VSS.n6433 VSS.n6432 1896.55
R294 VSS.n7992 VSS.n7991 1896.55
R295 VSS.n8584 VSS.n8583 1896.55
R296 VSS.n9176 VSS.n9175 1896.55
R297 VSS.n10360 VSS.n10359 1896.55
R298 VSS.n10952 VSS.n10951 1896.55
R299 VSS.n11544 VSS.n11543 1896.55
R300 VSS.n12136 VSS.n12135 1896.55
R301 VSS.n12728 VSS.n12727 1896.55
R302 VSS.n13320 VSS.n13319 1896.55
R303 VSS.n13912 VSS.n13911 1896.55
R304 VSS.n14504 VSS.n14503 1896.55
R305 VSS.n15096 VSS.n15095 1896.55
R306 VSS.n15688 VSS.n15687 1896.55
R307 VSS.n15921 VSS.n15920 1896.55
R308 VSS.n7400 VSS.n7399 1896.55
R309 VSS.n18712 VSS.n18711 1896.55
R310 VSS.n18538 VSS.n18537 1896.55
R311 VSS.n835 VSS.n834 1896.55
R312 VSS.t110 VSS.t105 1895.38
R313 VSS.t583 VSS.t353 1892.74
R314 VSS.t434 VSS.t488 1892.74
R315 VSS.t84 VSS.t476 1892.74
R316 VSS.t411 VSS.t531 1892.74
R317 VSS.t246 VSS.t9 1892.74
R318 VSS.t567 VSS.t52 1892.74
R319 VSS.t346 VSS.t142 1892.74
R320 VSS.t530 VSS.t359 1892.74
R321 VSS.t131 VSS.t457 1892.74
R322 VSS.t254 VSS.t208 1892.74
R323 VSS.t283 VSS.t590 1892.74
R324 VSS.t205 VSS.t632 1892.74
R325 VSS.t312 VSS.t309 1892.74
R326 VSS.t271 VSS.t564 1892.74
R327 VSS.t296 VSS.t211 1892.74
R328 VSS.t266 VSS.t261 1892.74
R329 VSS.t74 VSS.t551 1892.74
R330 VSS.t280 VSS.t508 1892.74
R331 VSS.t90 VSS.t366 1892.74
R332 VSS.t190 VSS.t228 1892.74
R333 VSS.t452 VSS.t548 1892.74
R334 VSS.t322 VSS.t23 1892.74
R335 VSS.t218 VSS.t420 1892.74
R336 VSS.t382 VSS.t48 1892.74
R337 VSS.t83 VSS.t545 1892.74
R338 VSS.t150 VSS.t325 1892.74
R339 VSS.t71 VSS.t482 1892.74
R340 VSS.t429 VSS.t424 1892.74
R341 VSS.t95 VSS.t273 1892.74
R342 VSS.t67 VSS.t123 1892.74
R343 VSS.t272 VSS.t607 1892.74
R344 VSS.t99 VSS.t96 1892.74
R345 VSS.t637 VSS.t238 1892.74
R346 VSS.t521 VSS.t202 1892.74
R347 VSS.t621 VSS.t337 1892.74
R348 VSS.t397 VSS.t145 1892.74
R349 VSS.t536 VSS.t625 1892.74
R350 VSS.t243 VSS.t251 1892.74
R351 VSS.t302 VSS.t354 1892.74
R352 VSS.t223 VSS.t102 1892.74
R353 VSS.t622 VSS.t415 1892.74
R354 VSS.t170 VSS.t445 1892.74
R355 VSS.t319 VSS.t554 1892.74
R356 VSS.t42 VSS.t155 1892.74
R357 VSS.t369 VSS.t6 1892.74
R358 VSS.t163 VSS.t158 1892.74
R359 VSS.t195 VSS.t604 1892.74
R360 VSS.t527 VSS.t332 1892.74
R361 VSS.t402 VSS.t138 1892.74
R362 VSS.t479 VSS.t181 1892.74
R363 VSS.t601 VSS.t20 1892.74
R364 VSS.t412 VSS.t557 1892.74
R365 VSS.t388 VSS.t469 1892.74
R366 VSS.t393 VSS.t68 1892.74
R367 VSS.t297 VSS.t387 1892.74
R368 VSS.t231 VSS.t468 1892.74
R369 VSS.t128 VSS.t572 1892.74
R370 VSS.t421 VSS.t141 1892.74
R371 VSS.t45 VSS.t522 1892.74
R372 VSS.t485 VSS.t87 1890.1
R373 VSS.n17125 VSS.t571 1791.5
R374 VSS.n17717 VSS.t631 1791.5
R375 VSS.n9767 VSS.t408 1791.5
R376 VSS.n16710 VSS.t171 1791.5
R377 VSS.n16117 VSS.t64 1791.5
R378 VSS.n2302 VSS.t511 1791.5
R379 VSS.n3258 VSS.t472 1791.5
R380 VSS.n3850 VSS.t578 1791.5
R381 VSS.n4442 VSS.t136 1791.5
R382 VSS.n5034 VSS.t267 1791.5
R383 VSS.n5267 VSS.t398 1791.5
R384 VSS.n5840 VSS.t507 1791.5
R385 VSS.n6432 VSS.t16 1791.5
R386 VSS.n7991 VSS.t30 1791.5
R387 VSS.n8583 VSS.t363 1791.5
R388 VSS.n9175 VSS.t496 1791.5
R389 VSS.n10359 VSS.t448 1791.5
R390 VSS.n10951 VSS.t380 1791.5
R391 VSS.n11543 VSS.t166 1791.5
R392 VSS.n12135 VSS.t57 1791.5
R393 VSS.n12727 VSS.t258 1791.5
R394 VSS.n13319 VSS.t443 1791.5
R395 VSS.n13911 VSS.t2 1791.5
R396 VSS.n14503 VSS.t458 1791.5
R397 VSS.n15095 VSS.t41 1791.5
R398 VSS.n15687 VSS.t151 1791.5
R399 VSS.n15920 VSS.t373 1791.5
R400 VSS.n7399 VSS.t112 1791.5
R401 VSS.n18711 VSS.t348 1791.5
R402 VSS.n18537 VSS.t439 1791.5
R403 VSS.n834 VSS.t185 1791.5
R404 VSS.t571 VSS.t597 1683.22
R405 VSS.t631 VSS.t119 1683.22
R406 VSS.t408 VSS.t34 1683.22
R407 VSS.t171 VSS.t489 1683.22
R408 VSS.t64 VSS.t560 1683.22
R409 VSS.t511 VSS.t77 1683.22
R410 VSS.t472 VSS.t463 1683.22
R411 VSS.t578 VSS.t610 1683.22
R412 VSS.t136 VSS.t515 1683.22
R413 VSS.t267 VSS.t175 1683.22
R414 VSS.t398 VSS.t217 1683.22
R415 VSS.t507 VSS.t115 1683.22
R416 VSS.t16 VSS.t617 1683.22
R417 VSS.t30 VSS.t242 1683.22
R418 VSS.t363 VSS.t498 1683.22
R419 VSS.t496 VSS.t544 1683.22
R420 VSS.t448 VSS.t279 1683.22
R421 VSS.t380 VSS.t586 1683.22
R422 VSS.t166 VSS.t227 1683.22
R423 VSS.t57 VSS.t305 1683.22
R424 VSS.t258 VSS.t26 1683.22
R425 VSS.t443 VSS.t331 1683.22
R426 VSS.t2 VSS.t540 1683.22
R427 VSS.t458 VSS.t315 1683.22
R428 VSS.t41 VSS.t579 1683.22
R429 VSS.t151 VSS.t593 1683.22
R430 VSS.t373 VSS.t293 1683.22
R431 VSS.t112 VSS.t430 1683.22
R432 VSS.t348 VSS.t340 1683.22
R433 VSS.t439 VSS.t289 1683.22
R434 VSS.t185 VSS.t186 1683.22
R435 VSS.t197 VSS.n17947 1560.55
R436 VSS.n17996 VSS.t372 1331.97
R437 VSS.n18060 VSS.t105 1095.38
R438 VSS.n17996 VSS.t353 1093.85
R439 VSS.t488 VSS.n18072 1093.85
R440 VSS.n15980 VSS.t476 1093.85
R441 VSS.n18046 VSS.t531 1093.85
R442 VSS.n18047 VSS.t52 1093.85
R443 VSS.n18048 VSS.t359 1093.85
R444 VSS.n18049 VSS.t208 1093.85
R445 VSS.n18050 VSS.t632 1093.85
R446 VSS.n18051 VSS.t564 1093.85
R447 VSS.n18052 VSS.t261 1093.85
R448 VSS.n18053 VSS.t508 1093.85
R449 VSS.n18054 VSS.t228 1093.85
R450 VSS.n18055 VSS.t23 1093.85
R451 VSS.n18056 VSS.t48 1093.85
R452 VSS.n18057 VSS.t325 1093.85
R453 VSS.n18058 VSS.t424 1093.85
R454 VSS.n18061 VSS.t607 1093.85
R455 VSS.n18062 VSS.t238 1093.85
R456 VSS.n18063 VSS.t337 1093.85
R457 VSS.n18064 VSS.t625 1093.85
R458 VSS.n18065 VSS.t354 1093.85
R459 VSS.n18066 VSS.t415 1093.85
R460 VSS.n18067 VSS.t554 1093.85
R461 VSS.n18068 VSS.t6 1093.85
R462 VSS.n18069 VSS.t604 1093.85
R463 VSS.n18070 VSS.t138 1093.85
R464 VSS.n18071 VSS.t20 1093.85
R465 VSS.n1020 VSS.t388 1093.85
R466 VSS.n1019 VSS.t231 1093.85
R467 VSS.n18045 VSS.t421 1093.85
R468 VSS.n18059 VSS.t87 1092.33
R469 VSS.t597 VSS.n17124 1045.79
R470 VSS.t119 VSS.n17716 1045.79
R471 VSS.t34 VSS.n9766 1045.79
R472 VSS.t489 VSS.n16709 1045.79
R473 VSS.t560 VSS.n16116 1045.79
R474 VSS.t77 VSS.n2301 1045.79
R475 VSS.t463 VSS.n3257 1045.79
R476 VSS.t610 VSS.n3849 1045.79
R477 VSS.t515 VSS.n4441 1045.79
R478 VSS.t175 VSS.n5033 1045.79
R479 VSS.t217 VSS.n5266 1045.79
R480 VSS.t115 VSS.n5839 1045.79
R481 VSS.t617 VSS.n6431 1045.79
R482 VSS.t242 VSS.n7990 1045.79
R483 VSS.t498 VSS.n8582 1045.79
R484 VSS.t544 VSS.n9174 1045.79
R485 VSS.t279 VSS.n10358 1045.79
R486 VSS.t586 VSS.n10950 1045.79
R487 VSS.t227 VSS.n11542 1045.79
R488 VSS.t305 VSS.n12134 1045.79
R489 VSS.t26 VSS.n12726 1045.79
R490 VSS.t331 VSS.n13318 1045.79
R491 VSS.t540 VSS.n13910 1045.79
R492 VSS.t315 VSS.n14502 1045.79
R493 VSS.t579 VSS.n15094 1045.79
R494 VSS.t593 VSS.n15686 1045.79
R495 VSS.t293 VSS.n15919 1045.79
R496 VSS.t430 VSS.n7398 1045.79
R497 VSS.t340 VSS.n18710 1045.79
R498 VSS.t289 VSS.n18536 1045.79
R499 VSS.t186 VSS.n833 1045.79
R500 VSS.n17997 VSS.n1155 1017.62
R501 VSS.n17997 VSS.n17996 772.908
R502 VSS.n17496 VSS.t381 758.37
R503 VSS.t381 VSS.t614 746.255
R504 VSS.n15979 VSS.n6483 626.798
R505 VSS.n17124 VSS.n17123 590.341
R506 VSS.n16865 VSS.n25 590.341
R507 VSS.n17716 VSS.n17715 590.341
R508 VSS.n17279 VSS.n23 590.341
R509 VSS.n18536 VSS.n18535 590.341
R510 VSS.n18436 VSS.n10 590.341
R511 VSS.n9766 VSS.n9765 590.341
R512 VSS.n9330 VSS.n32 590.341
R513 VSS.n16709 VSS.n16708 590.341
R514 VSS.n16272 VSS.n22 590.341
R515 VSS.n16116 VSS.n16115 590.341
R516 VSS.n1444 VSS.n26 590.341
R517 VSS.n2301 VSS.n2300 590.341
R518 VSS.n2205 VSS.n21 590.341
R519 VSS.n3257 VSS.n3256 590.341
R520 VSS.n2821 VSS.n27 590.341
R521 VSS.n3849 VSS.n3848 590.341
R522 VSS.n3413 VSS.n20 590.341
R523 VSS.n4441 VSS.n4440 590.341
R524 VSS.n4005 VSS.n28 590.341
R525 VSS.n5033 VSS.n5032 590.341
R526 VSS.n4597 VSS.n19 590.341
R527 VSS.n5266 VSS.n5265 590.341
R528 VSS.n2801 VSS.n29 590.341
R529 VSS.n5839 VSS.n5838 590.341
R530 VSS.n18878 VSS.n6 590.341
R531 VSS.n6431 VSS.n6430 590.341
R532 VSS.n6335 VSS.n30 590.341
R533 VSS.n7990 VSS.n7989 590.341
R534 VSS.n7554 VSS.n18 590.341
R535 VSS.n8582 VSS.n8581 590.341
R536 VSS.n8146 VSS.n31 590.341
R537 VSS.n9174 VSS.n9173 590.341
R538 VSS.n8738 VSS.n17 590.341
R539 VSS.n10358 VSS.n10357 590.341
R540 VSS.n9922 VSS.n16 590.341
R541 VSS.n10950 VSS.n10949 590.341
R542 VSS.n10514 VSS.n33 590.341
R543 VSS.n11542 VSS.n11541 590.341
R544 VSS.n11106 VSS.n15 590.341
R545 VSS.n12134 VSS.n12133 590.341
R546 VSS.n11698 VSS.n34 590.341
R547 VSS.n12726 VSS.n12725 590.341
R548 VSS.n12290 VSS.n14 590.341
R549 VSS.n13318 VSS.n13317 590.341
R550 VSS.n12882 VSS.n35 590.341
R551 VSS.n13910 VSS.n13909 590.341
R552 VSS.n13474 VSS.n13 590.341
R553 VSS.n14502 VSS.n14501 590.341
R554 VSS.n14066 VSS.n36 590.341
R555 VSS.n15094 VSS.n15093 590.341
R556 VSS.n14658 VSS.n12 590.341
R557 VSS.n15686 VSS.n15685 590.341
R558 VSS.n15250 VSS.n37 590.341
R559 VSS.n15919 VSS.n15918 590.341
R560 VSS.n6941 VSS.n11 590.341
R561 VSS.n7398 VSS.n7397 590.341
R562 VSS.n6961 VSS.n38 590.341
R563 VSS.n18710 VSS.n18709 590.341
R564 VSS.n59 VSS.n39 590.341
R565 VSS.n833 VSS.n832 590.341
R566 VSS.n18876 VSS.n18875 590.341
R567 VSS.n17947 VSS.n17946 590.341
R568 VSS.n1423 VSS.n24 590.341
R569 VSS.n17000 VSS.n16989 585
R570 VSS.n17002 VSS.n16989 585
R571 VSS.n16988 VSS.n16987 585
R572 VSS.n17029 VSS.n16988 585
R573 VSS.n17049 VSS.n17048 585
R574 VSS.n17050 VSS.n17049 585
R575 VSS.n16955 VSS.n16954 585
R576 VSS.n16954 VSS.n16953 585
R577 VSS.n17084 VSS.n17083 585
R578 VSS.n17083 VSS.t247 585
R579 VSS.n17102 VSS.n17101 585
R580 VSS.n17103 VSS.n17102 585
R581 VSS.n16973 VSS.n16971 585
R582 VSS.n17052 VSS.n16973 585
R583 VSS.n16972 VSS.n16970 585
R584 VSS.n17051 VSS.n16972 585
R585 VSS.n17032 VSS.n17031 585
R586 VSS.n17031 VSS.n17030 585
R587 VSS.n16952 VSS.n16951 585
R588 VSS.n17082 VSS.n16952 585
R589 VSS.n16937 VSS.n16936 585
R590 VSS.n17104 VSS.n16937 585
R591 VSS.n17005 VSS.n17004 585
R592 VSS.n17004 VSS.n17003 585
R593 VSS.n17115 VSS.n17111 585
R594 VSS.n17119 VSS.n17111 585
R595 VSS.n17163 VSS.n17162 585
R596 VSS.n17164 VSS.n17163 585
R597 VSS.n16914 VSS.n16912 585
R598 VSS.n17166 VSS.n16914 585
R599 VSS.n17219 VSS.n17218 585
R600 VSS.n17218 VSS.n17217 585
R601 VSS.n16880 VSS.n16879 585
R602 VSS.t173 VSS.n16880 585
R603 VSS.n17260 VSS.n17259 585
R604 VSS.n17261 VSS.n17260 585
R605 VSS.n17258 VSS.n16866 585
R606 VSS.n17262 VSS.n16866 585
R607 VSS.n17239 VSS.n17238 585
R608 VSS.n17238 VSS.n17237 585
R609 VSS.n17220 VSS.n16882 585
R610 VSS.n16882 VSS.n16881 585
R611 VSS.n16917 VSS.n16916 585
R612 VSS.n16916 VSS.n16915 585
R613 VSS.n17169 VSS.n17168 585
R614 VSS.n17168 VSS.n17167 585
R615 VSS.n17263 VSS.n16867 585
R616 VSS.n17106 VSS.n17105 585
R617 VSS.n17117 VSS.n17116 585
R618 VSS.n17118 VSS.n17117 585
R619 VSS.n17414 VSS.n17403 585
R620 VSS.n17416 VSS.n17403 585
R621 VSS.n17402 VSS.n17401 585
R622 VSS.n17621 VSS.n17402 585
R623 VSS.n17641 VSS.n17640 585
R624 VSS.n17642 VSS.n17641 585
R625 VSS.n17369 VSS.n17368 585
R626 VSS.n17368 VSS.n17367 585
R627 VSS.n17676 VSS.n17675 585
R628 VSS.n17675 VSS.t46 585
R629 VSS.n17694 VSS.n17693 585
R630 VSS.n17695 VSS.n17694 585
R631 VSS.n17387 VSS.n17385 585
R632 VSS.n17644 VSS.n17387 585
R633 VSS.n17386 VSS.n17384 585
R634 VSS.n17643 VSS.n17386 585
R635 VSS.n17624 VSS.n17623 585
R636 VSS.n17623 VSS.n17622 585
R637 VSS.n17366 VSS.n17365 585
R638 VSS.n17674 VSS.n17366 585
R639 VSS.n17351 VSS.n17350 585
R640 VSS.n17696 VSS.n17351 585
R641 VSS.n17419 VSS.n17418 585
R642 VSS.n17418 VSS.n17417 585
R643 VSS.n17707 VSS.n17703 585
R644 VSS.n17711 VSS.n17703 585
R645 VSS.n17755 VSS.n17754 585
R646 VSS.n17756 VSS.n17755 585
R647 VSS.n17328 VSS.n17326 585
R648 VSS.n17758 VSS.n17328 585
R649 VSS.n17811 VSS.n17810 585
R650 VSS.n17810 VSS.n17809 585
R651 VSS.n17294 VSS.n17293 585
R652 VSS.t568 VSS.n17294 585
R653 VSS.n17852 VSS.n17851 585
R654 VSS.n17853 VSS.n17852 585
R655 VSS.n17850 VSS.n17280 585
R656 VSS.n17854 VSS.n17280 585
R657 VSS.n17831 VSS.n17830 585
R658 VSS.n17830 VSS.n17829 585
R659 VSS.n17812 VSS.n17296 585
R660 VSS.n17296 VSS.n17295 585
R661 VSS.n17331 VSS.n17330 585
R662 VSS.n17330 VSS.n17329 585
R663 VSS.n17761 VSS.n17760 585
R664 VSS.n17760 VSS.n17759 585
R665 VSS.n17855 VSS.n17281 585
R666 VSS.n17698 VSS.n17697 585
R667 VSS.n17709 VSS.n17708 585
R668 VSS.n17710 VSS.n17709 585
R669 VSS.n287 VSS.n286 585
R670 VSS.n18074 VSS.n287 585
R671 VSS.n18100 VSS.n18099 585
R672 VSS.n18101 VSS.n18100 585
R673 VSS.n272 VSS.n270 585
R674 VSS.n18105 VSS.n272 585
R675 VSS.n242 VSS.n240 585
R676 VSS.n18136 VSS.n242 585
R677 VSS.n220 VSS.n219 585
R678 VSS.n18137 VSS.n219 585
R679 VSS.n228 VSS.n218 585
R680 VSS.n18168 VSS.n218 585
R681 VSS.n18134 VSS.n18133 585
R682 VSS.n18135 VSS.n18134 585
R683 VSS.n18103 VSS.n252 585
R684 VSS.n18104 VSS.n18103 585
R685 VSS.n18098 VSS.n271 585
R686 VSS.n18102 VSS.n271 585
R687 VSS.n249 VSS.n248 585
R688 VSS.n18138 VSS.n249 585
R689 VSS.n18170 VSS.n217 585
R690 VSS.n18170 VSS.n18169 585
R691 VSS.n18077 VSS.n18076 585
R692 VSS.n18076 VSS.n18075 585
R693 VSS.n9464 VSS.n9453 585
R694 VSS.n9466 VSS.n9453 585
R695 VSS.n9452 VSS.n9451 585
R696 VSS.n9671 VSS.n9452 585
R697 VSS.n9691 VSS.n9690 585
R698 VSS.n9692 VSS.n9691 585
R699 VSS.n9419 VSS.n9418 585
R700 VSS.n9418 VSS.n9417 585
R701 VSS.n9726 VSS.n9725 585
R702 VSS.n9725 VSS.t65 585
R703 VSS.n9744 VSS.n9743 585
R704 VSS.n9745 VSS.n9744 585
R705 VSS.n9437 VSS.n9435 585
R706 VSS.n9694 VSS.n9437 585
R707 VSS.n9436 VSS.n9434 585
R708 VSS.n9693 VSS.n9436 585
R709 VSS.n9674 VSS.n9673 585
R710 VSS.n9673 VSS.n9672 585
R711 VSS.n9416 VSS.n9415 585
R712 VSS.n9724 VSS.n9416 585
R713 VSS.n9401 VSS.n9400 585
R714 VSS.n9746 VSS.n9401 585
R715 VSS.n9469 VSS.n9468 585
R716 VSS.n9468 VSS.n9467 585
R717 VSS.n9757 VSS.n9753 585
R718 VSS.n9761 VSS.n9753 585
R719 VSS.n9805 VSS.n9804 585
R720 VSS.n9806 VSS.n9805 585
R721 VSS.n9378 VSS.n9376 585
R722 VSS.n9808 VSS.n9378 585
R723 VSS.n9861 VSS.n9860 585
R724 VSS.n9860 VSS.n9859 585
R725 VSS.n9344 VSS.n9343 585
R726 VSS.t449 VSS.n9344 585
R727 VSS.n9903 VSS.n9902 585
R728 VSS.n9904 VSS.n9903 585
R729 VSS.n9901 VSS.n9331 585
R730 VSS.n9905 VSS.n9331 585
R731 VSS.n9881 VSS.n9880 585
R732 VSS.n9880 VSS.n9879 585
R733 VSS.n9862 VSS.n9346 585
R734 VSS.n9346 VSS.n9345 585
R735 VSS.n9381 VSS.n9380 585
R736 VSS.n9380 VSS.n9379 585
R737 VSS.n9811 VSS.n9810 585
R738 VSS.n9810 VSS.n9809 585
R739 VSS.n9906 VSS.n9332 585
R740 VSS.n9748 VSS.n9747 585
R741 VSS.n9759 VSS.n9758 585
R742 VSS.n9760 VSS.n9759 585
R743 VSS.n9545 VSS.n9544 585
R744 VSS.n9547 VSS.n9545 585
R745 VSS.n9573 VSS.n9572 585
R746 VSS.n9574 VSS.n9573 585
R747 VSS.n9530 VSS.n9528 585
R748 VSS.n9578 VSS.n9530 585
R749 VSS.n9500 VSS.n9498 585
R750 VSS.n9609 VSS.n9500 585
R751 VSS.n9478 VSS.n9477 585
R752 VSS.n9610 VSS.n9477 585
R753 VSS.n9486 VSS.n9476 585
R754 VSS.n9641 VSS.n9476 585
R755 VSS.n9607 VSS.n9606 585
R756 VSS.n9608 VSS.n9607 585
R757 VSS.n9571 VSS.n9529 585
R758 VSS.n9575 VSS.n9529 585
R759 VSS.n9576 VSS.n9510 585
R760 VSS.n9577 VSS.n9576 585
R761 VSS.n9507 VSS.n9506 585
R762 VSS.n9611 VSS.n9507 585
R763 VSS.n9643 VSS.n9475 585
R764 VSS.n9643 VSS.n9642 585
R765 VSS.n9550 VSS.n9549 585
R766 VSS.n9549 VSS.n9548 585
R767 VSS.n16406 VSS.n16395 585
R768 VSS.n16408 VSS.n16395 585
R769 VSS.n16394 VSS.n16393 585
R770 VSS.n16614 VSS.n16394 585
R771 VSS.n16634 VSS.n16633 585
R772 VSS.n16635 VSS.n16634 585
R773 VSS.n16361 VSS.n16360 585
R774 VSS.n16360 VSS.n16359 585
R775 VSS.n16669 VSS.n16668 585
R776 VSS.n16668 VSS.t143 585
R777 VSS.n16687 VSS.n16686 585
R778 VSS.n16688 VSS.n16687 585
R779 VSS.n16379 VSS.n16377 585
R780 VSS.n16637 VSS.n16379 585
R781 VSS.n16378 VSS.n16376 585
R782 VSS.n16636 VSS.n16378 585
R783 VSS.n16617 VSS.n16616 585
R784 VSS.n16616 VSS.n16615 585
R785 VSS.n16358 VSS.n16357 585
R786 VSS.n16667 VSS.n16358 585
R787 VSS.n16343 VSS.n16342 585
R788 VSS.n16689 VSS.n16343 585
R789 VSS.n16411 VSS.n16410 585
R790 VSS.n16410 VSS.n16409 585
R791 VSS.n16700 VSS.n16696 585
R792 VSS.n16704 VSS.n16696 585
R793 VSS.n16748 VSS.n16747 585
R794 VSS.n16749 VSS.n16748 585
R795 VSS.n16320 VSS.n16318 585
R796 VSS.n16751 VSS.n16320 585
R797 VSS.n16804 VSS.n16803 585
R798 VSS.n16803 VSS.n16802 585
R799 VSS.n16286 VSS.n16285 585
R800 VSS.t62 VSS.n16286 585
R801 VSS.n16846 VSS.n16845 585
R802 VSS.n16847 VSS.n16846 585
R803 VSS.n16844 VSS.n16273 585
R804 VSS.n16848 VSS.n16273 585
R805 VSS.n16824 VSS.n16823 585
R806 VSS.n16823 VSS.n16822 585
R807 VSS.n16805 VSS.n16288 585
R808 VSS.n16288 VSS.n16287 585
R809 VSS.n16323 VSS.n16322 585
R810 VSS.n16322 VSS.n16321 585
R811 VSS.n16754 VSS.n16753 585
R812 VSS.n16753 VSS.n16752 585
R813 VSS.n16849 VSS.n16274 585
R814 VSS.n16691 VSS.n16690 585
R815 VSS.n16702 VSS.n16701 585
R816 VSS.n16703 VSS.n16702 585
R817 VSS.n16481 VSS.n16470 585
R818 VSS.n16483 VSS.n16470 585
R819 VSS.n16469 VSS.n16468 585
R820 VSS.n16509 VSS.n16469 585
R821 VSS.n16529 VSS.n16528 585
R822 VSS.n16530 VSS.n16529 585
R823 VSS.n16436 VSS.n16435 585
R824 VSS.n16435 VSS.n16434 585
R825 VSS.n16565 VSS.n16564 585
R826 VSS.n16564 VSS.n16563 585
R827 VSS.n16583 VSS.n16582 585
R828 VSS.n16584 VSS.n16583 585
R829 VSS.n16456 VSS.n16454 585
R830 VSS.n16532 VSS.n16456 585
R831 VSS.n16455 VSS.n16453 585
R832 VSS.n16531 VSS.n16455 585
R833 VSS.n16512 VSS.n16511 585
R834 VSS.n16511 VSS.n16510 585
R835 VSS.n16433 VSS.n16432 585
R836 VSS.n16562 VSS.n16433 585
R837 VSS.n16418 VSS.n16417 585
R838 VSS.n16585 VSS.n16418 585
R839 VSS.n16486 VSS.n16485 585
R840 VSS.n16485 VSS.n16484 585
R841 VSS.n1753 VSS.n1567 585
R842 VSS.n1751 VSS.n1567 585
R843 VSS.n1566 VSS.n1565 585
R844 VSS.n16021 VSS.n1566 585
R845 VSS.n16041 VSS.n16040 585
R846 VSS.n16042 VSS.n16041 585
R847 VSS.n1533 VSS.n1532 585
R848 VSS.n1532 VSS.n1531 585
R849 VSS.n16076 VSS.n16075 585
R850 VSS.n16075 VSS.t455 585
R851 VSS.n16094 VSS.n16093 585
R852 VSS.n16095 VSS.n16094 585
R853 VSS.n1551 VSS.n1549 585
R854 VSS.n16044 VSS.n1551 585
R855 VSS.n1550 VSS.n1548 585
R856 VSS.n16043 VSS.n1550 585
R857 VSS.n16024 VSS.n16023 585
R858 VSS.n16023 VSS.n16022 585
R859 VSS.n1530 VSS.n1529 585
R860 VSS.n16074 VSS.n1530 585
R861 VSS.n1515 VSS.n1514 585
R862 VSS.n16096 VSS.n1515 585
R863 VSS.n1755 VSS.n1754 585
R864 VSS.n1755 VSS.n1752 585
R865 VSS.n16107 VSS.n16103 585
R866 VSS.n16111 VSS.n16103 585
R867 VSS.n16155 VSS.n16154 585
R868 VSS.n16156 VSS.n16155 585
R869 VSS.n1492 VSS.n1490 585
R870 VSS.n16158 VSS.n1492 585
R871 VSS.n16211 VSS.n16210 585
R872 VSS.n16210 VSS.n16209 585
R873 VSS.n1458 VSS.n1457 585
R874 VSS.t512 VSS.n1458 585
R875 VSS.n16253 VSS.n16252 585
R876 VSS.n16254 VSS.n16253 585
R877 VSS.n16251 VSS.n1445 585
R878 VSS.n16255 VSS.n1445 585
R879 VSS.n16231 VSS.n16230 585
R880 VSS.n16230 VSS.n16229 585
R881 VSS.n16212 VSS.n1460 585
R882 VSS.n1460 VSS.n1459 585
R883 VSS.n1495 VSS.n1494 585
R884 VSS.n1494 VSS.n1493 585
R885 VSS.n16161 VSS.n16160 585
R886 VSS.n16160 VSS.n16159 585
R887 VSS.n16256 VSS.n1446 585
R888 VSS.n16098 VSS.n16097 585
R889 VSS.n16109 VSS.n16108 585
R890 VSS.n16110 VSS.n16109 585
R891 VSS.n1646 VSS.n1635 585
R892 VSS.n1648 VSS.n1635 585
R893 VSS.n1634 VSS.n1633 585
R894 VSS.n1674 VSS.n1634 585
R895 VSS.n1694 VSS.n1693 585
R896 VSS.n1695 VSS.n1694 585
R897 VSS.n1601 VSS.n1600 585
R898 VSS.n1600 VSS.n1599 585
R899 VSS.n1730 VSS.n1729 585
R900 VSS.n1729 VSS.n1728 585
R901 VSS.n1748 VSS.n1747 585
R902 VSS.n1749 VSS.n1748 585
R903 VSS.n1621 VSS.n1619 585
R904 VSS.n1697 VSS.n1621 585
R905 VSS.n1620 VSS.n1618 585
R906 VSS.n1696 VSS.n1620 585
R907 VSS.n1677 VSS.n1676 585
R908 VSS.n1676 VSS.n1675 585
R909 VSS.n1598 VSS.n1597 585
R910 VSS.n1727 VSS.n1598 585
R911 VSS.n1583 VSS.n1582 585
R912 VSS.n1750 VSS.n1583 585
R913 VSS.n1651 VSS.n1650 585
R914 VSS.n1650 VSS.n1649 585
R915 VSS.n2003 VSS.n2002 585
R916 VSS.n2002 VSS.n2001 585
R917 VSS.n2026 VSS.n2025 585
R918 VSS.n2027 VSS.n2026 585
R919 VSS.n2032 VSS.n1995 585
R920 VSS.n1995 VSS.n1994 585
R921 VSS.n2040 VSS.n1991 585
R922 VSS.n1991 VSS.n1990 585
R923 VSS.n2055 VSS.n2054 585
R924 VSS.n2054 VSS.t284 585
R925 VSS.n2067 VSS.n2066 585
R926 VSS.n2068 VSS.n2067 585
R927 VSS.n2039 VSS.n2038 585
R928 VSS.n2038 VSS.n2037 585
R929 VSS.n2034 VSS.n2033 585
R930 VSS.n2035 VSS.n2034 585
R931 VSS.n2024 VSS.n1998 585
R932 VSS.n2028 VSS.n1998 585
R933 VSS.n1989 VSS.n1988 585
R934 VSS.n2053 VSS.n1989 585
R935 VSS.n1980 VSS.n1979 585
R936 VSS.n2069 VSS.n1980 585
R937 VSS.n1761 VSS.n1760 585
R938 VSS.n1760 VSS.n1759 585
R939 VSS.n2077 VSS.n2074 585
R940 VSS.n2296 VSS.n2074 585
R941 VSS.n2104 VSS.n2103 585
R942 VSS.n2280 VSS.n2104 585
R943 VSS.n2267 VSS.n2266 585
R944 VSS.n2266 VSS.n2265 585
R945 VSS.n2187 VSS.n2186 585
R946 VSS.n2188 VSS.n2187 585
R947 VSS.n2195 VSS.n2194 585
R948 VSS.t473 VSS.n2195 585
R949 VSS.n2176 VSS.n2174 585
R950 VSS.n2229 VSS.n2176 585
R951 VSS.n2227 VSS.n2226 585
R952 VSS.n2228 VSS.n2227 585
R953 VSS.n2193 VSS.n2175 585
R954 VSS.n2196 VSS.n2175 585
R955 VSS.n2190 VSS.n2157 585
R956 VSS.n2190 VSS.n2189 585
R957 VSS.n2283 VSS.n2282 585
R958 VSS.n2282 VSS.n2281 585
R959 VSS.n2268 VSS.n2106 585
R960 VSS.n2106 VSS.n2105 585
R961 VSS.n2204 VSS.n2203 585
R962 VSS.n2071 VSS.n2070 585
R963 VSS.n2294 VSS.n2293 585
R964 VSS.n2295 VSS.n2294 585
R965 VSS.n1837 VSS.n1836 585
R966 VSS.n1839 VSS.n1837 585
R967 VSS.n1865 VSS.n1864 585
R968 VSS.n1866 VSS.n1865 585
R969 VSS.n1822 VSS.n1820 585
R970 VSS.n1870 VSS.n1822 585
R971 VSS.n1792 VSS.n1790 585
R972 VSS.n1901 VSS.n1792 585
R973 VSS.n1770 VSS.n1769 585
R974 VSS.n1902 VSS.n1769 585
R975 VSS.n1778 VSS.n1768 585
R976 VSS.n1933 VSS.n1768 585
R977 VSS.n1899 VSS.n1898 585
R978 VSS.n1900 VSS.n1899 585
R979 VSS.n1868 VSS.n1802 585
R980 VSS.n1869 VSS.n1868 585
R981 VSS.n1863 VSS.n1821 585
R982 VSS.n1867 VSS.n1821 585
R983 VSS.n1799 VSS.n1798 585
R984 VSS.n1903 VSS.n1799 585
R985 VSS.n1935 VSS.n1767 585
R986 VSS.n1935 VSS.n1934 585
R987 VSS.n1842 VSS.n1841 585
R988 VSS.n1841 VSS.n1840 585
R989 VSS.n2955 VSS.n2944 585
R990 VSS.n2957 VSS.n2944 585
R991 VSS.n2943 VSS.n2942 585
R992 VSS.n3162 VSS.n2943 585
R993 VSS.n3182 VSS.n3181 585
R994 VSS.n3183 VSS.n3182 585
R995 VSS.n2910 VSS.n2909 585
R996 VSS.n2909 VSS.n2908 585
R997 VSS.n3217 VSS.n3216 585
R998 VSS.n3216 VSS.t313 585
R999 VSS.n3235 VSS.n3234 585
R1000 VSS.n3236 VSS.n3235 585
R1001 VSS.n2928 VSS.n2926 585
R1002 VSS.n3185 VSS.n2928 585
R1003 VSS.n2927 VSS.n2925 585
R1004 VSS.n3184 VSS.n2927 585
R1005 VSS.n3165 VSS.n3164 585
R1006 VSS.n3164 VSS.n3163 585
R1007 VSS.n2907 VSS.n2906 585
R1008 VSS.n3215 VSS.n2907 585
R1009 VSS.n2892 VSS.n2891 585
R1010 VSS.n3237 VSS.n2892 585
R1011 VSS.n2960 VSS.n2959 585
R1012 VSS.n2959 VSS.n2958 585
R1013 VSS.n3248 VSS.n3244 585
R1014 VSS.n3252 VSS.n3244 585
R1015 VSS.n3296 VSS.n3295 585
R1016 VSS.n3297 VSS.n3296 585
R1017 VSS.n2869 VSS.n2867 585
R1018 VSS.n3299 VSS.n2869 585
R1019 VSS.n3352 VSS.n3351 585
R1020 VSS.n3351 VSS.n3350 585
R1021 VSS.n2835 VSS.n2834 585
R1022 VSS.t575 VSS.n2835 585
R1023 VSS.n3394 VSS.n3393 585
R1024 VSS.n3395 VSS.n3394 585
R1025 VSS.n3392 VSS.n2822 585
R1026 VSS.n3396 VSS.n2822 585
R1027 VSS.n3372 VSS.n3371 585
R1028 VSS.n3371 VSS.n3370 585
R1029 VSS.n3353 VSS.n2837 585
R1030 VSS.n2837 VSS.n2836 585
R1031 VSS.n2872 VSS.n2871 585
R1032 VSS.n2871 VSS.n2870 585
R1033 VSS.n3302 VSS.n3301 585
R1034 VSS.n3301 VSS.n3300 585
R1035 VSS.n3397 VSS.n2823 585
R1036 VSS.n3239 VSS.n3238 585
R1037 VSS.n3250 VSS.n3249 585
R1038 VSS.n3251 VSS.n3250 585
R1039 VSS.n3036 VSS.n3035 585
R1040 VSS.n3038 VSS.n3036 585
R1041 VSS.n3064 VSS.n3063 585
R1042 VSS.n3065 VSS.n3064 585
R1043 VSS.n3021 VSS.n3019 585
R1044 VSS.n3069 VSS.n3021 585
R1045 VSS.n2991 VSS.n2989 585
R1046 VSS.n3100 VSS.n2991 585
R1047 VSS.n2969 VSS.n2968 585
R1048 VSS.n3101 VSS.n2968 585
R1049 VSS.n2977 VSS.n2967 585
R1050 VSS.n3132 VSS.n2967 585
R1051 VSS.n3098 VSS.n3097 585
R1052 VSS.n3099 VSS.n3098 585
R1053 VSS.n3067 VSS.n3001 585
R1054 VSS.n3068 VSS.n3067 585
R1055 VSS.n3062 VSS.n3020 585
R1056 VSS.n3066 VSS.n3020 585
R1057 VSS.n2998 VSS.n2997 585
R1058 VSS.n3102 VSS.n2998 585
R1059 VSS.n3134 VSS.n2966 585
R1060 VSS.n3134 VSS.n3133 585
R1061 VSS.n3041 VSS.n3040 585
R1062 VSS.n3040 VSS.n3039 585
R1063 VSS.n3547 VSS.n3536 585
R1064 VSS.n3549 VSS.n3536 585
R1065 VSS.n3535 VSS.n3534 585
R1066 VSS.n3754 VSS.n3535 585
R1067 VSS.n3774 VSS.n3773 585
R1068 VSS.n3775 VSS.n3774 585
R1069 VSS.n3502 VSS.n3501 585
R1070 VSS.n3501 VSS.n3500 585
R1071 VSS.n3809 VSS.n3808 585
R1072 VSS.n3808 VSS.t294 585
R1073 VSS.n3827 VSS.n3826 585
R1074 VSS.n3828 VSS.n3827 585
R1075 VSS.n3520 VSS.n3518 585
R1076 VSS.n3777 VSS.n3520 585
R1077 VSS.n3519 VSS.n3517 585
R1078 VSS.n3776 VSS.n3519 585
R1079 VSS.n3757 VSS.n3756 585
R1080 VSS.n3756 VSS.n3755 585
R1081 VSS.n3499 VSS.n3498 585
R1082 VSS.n3807 VSS.n3499 585
R1083 VSS.n3484 VSS.n3483 585
R1084 VSS.n3829 VSS.n3484 585
R1085 VSS.n3552 VSS.n3551 585
R1086 VSS.n3551 VSS.n3550 585
R1087 VSS.n3840 VSS.n3836 585
R1088 VSS.n3844 VSS.n3836 585
R1089 VSS.n3888 VSS.n3887 585
R1090 VSS.n3889 VSS.n3888 585
R1091 VSS.n3461 VSS.n3459 585
R1092 VSS.n3891 VSS.n3461 585
R1093 VSS.n3944 VSS.n3943 585
R1094 VSS.n3943 VSS.n3942 585
R1095 VSS.n3427 VSS.n3426 585
R1096 VSS.t134 VSS.n3427 585
R1097 VSS.n3986 VSS.n3985 585
R1098 VSS.n3987 VSS.n3986 585
R1099 VSS.n3984 VSS.n3414 585
R1100 VSS.n3988 VSS.n3414 585
R1101 VSS.n3964 VSS.n3963 585
R1102 VSS.n3963 VSS.n3962 585
R1103 VSS.n3945 VSS.n3429 585
R1104 VSS.n3429 VSS.n3428 585
R1105 VSS.n3464 VSS.n3463 585
R1106 VSS.n3463 VSS.n3462 585
R1107 VSS.n3894 VSS.n3893 585
R1108 VSS.n3893 VSS.n3892 585
R1109 VSS.n3989 VSS.n3415 585
R1110 VSS.n3831 VSS.n3830 585
R1111 VSS.n3842 VSS.n3841 585
R1112 VSS.n3843 VSS.n3842 585
R1113 VSS.n3628 VSS.n3627 585
R1114 VSS.n3630 VSS.n3628 585
R1115 VSS.n3656 VSS.n3655 585
R1116 VSS.n3657 VSS.n3656 585
R1117 VSS.n3613 VSS.n3611 585
R1118 VSS.n3661 VSS.n3613 585
R1119 VSS.n3583 VSS.n3581 585
R1120 VSS.n3692 VSS.n3583 585
R1121 VSS.n3561 VSS.n3560 585
R1122 VSS.n3693 VSS.n3560 585
R1123 VSS.n3569 VSS.n3559 585
R1124 VSS.n3724 VSS.n3559 585
R1125 VSS.n3690 VSS.n3689 585
R1126 VSS.n3691 VSS.n3690 585
R1127 VSS.n3659 VSS.n3593 585
R1128 VSS.n3660 VSS.n3659 585
R1129 VSS.n3654 VSS.n3612 585
R1130 VSS.n3658 VSS.n3612 585
R1131 VSS.n3590 VSS.n3589 585
R1132 VSS.n3694 VSS.n3590 585
R1133 VSS.n3726 VSS.n3558 585
R1134 VSS.n3726 VSS.n3725 585
R1135 VSS.n3633 VSS.n3632 585
R1136 VSS.n3632 VSS.n3631 585
R1137 VSS.n4139 VSS.n4128 585
R1138 VSS.n4141 VSS.n4128 585
R1139 VSS.n4127 VSS.n4126 585
R1140 VSS.n4346 VSS.n4127 585
R1141 VSS.n4366 VSS.n4365 585
R1142 VSS.n4367 VSS.n4366 585
R1143 VSS.n4094 VSS.n4093 585
R1144 VSS.n4093 VSS.n4092 585
R1145 VSS.n4401 VSS.n4400 585
R1146 VSS.n4400 VSS.t75 585
R1147 VSS.n4419 VSS.n4418 585
R1148 VSS.n4420 VSS.n4419 585
R1149 VSS.n4112 VSS.n4110 585
R1150 VSS.n4369 VSS.n4112 585
R1151 VSS.n4111 VSS.n4109 585
R1152 VSS.n4368 VSS.n4111 585
R1153 VSS.n4349 VSS.n4348 585
R1154 VSS.n4348 VSS.n4347 585
R1155 VSS.n4091 VSS.n4090 585
R1156 VSS.n4399 VSS.n4091 585
R1157 VSS.n4076 VSS.n4075 585
R1158 VSS.n4421 VSS.n4076 585
R1159 VSS.n4144 VSS.n4143 585
R1160 VSS.n4143 VSS.n4142 585
R1161 VSS.n4432 VSS.n4428 585
R1162 VSS.n4436 VSS.n4428 585
R1163 VSS.n4480 VSS.n4479 585
R1164 VSS.n4481 VSS.n4480 585
R1165 VSS.n4053 VSS.n4051 585
R1166 VSS.n4483 VSS.n4053 585
R1167 VSS.n4536 VSS.n4535 585
R1168 VSS.n4535 VSS.n4534 585
R1169 VSS.n4019 VSS.n4018 585
R1170 VSS.t269 VSS.n4019 585
R1171 VSS.n4578 VSS.n4577 585
R1172 VSS.n4579 VSS.n4578 585
R1173 VSS.n4576 VSS.n4006 585
R1174 VSS.n4580 VSS.n4006 585
R1175 VSS.n4556 VSS.n4555 585
R1176 VSS.n4555 VSS.n4554 585
R1177 VSS.n4537 VSS.n4021 585
R1178 VSS.n4021 VSS.n4020 585
R1179 VSS.n4056 VSS.n4055 585
R1180 VSS.n4055 VSS.n4054 585
R1181 VSS.n4486 VSS.n4485 585
R1182 VSS.n4485 VSS.n4484 585
R1183 VSS.n4581 VSS.n4007 585
R1184 VSS.n4423 VSS.n4422 585
R1185 VSS.n4434 VSS.n4433 585
R1186 VSS.n4435 VSS.n4434 585
R1187 VSS.n4220 VSS.n4219 585
R1188 VSS.n4222 VSS.n4220 585
R1189 VSS.n4248 VSS.n4247 585
R1190 VSS.n4249 VSS.n4248 585
R1191 VSS.n4205 VSS.n4203 585
R1192 VSS.n4253 VSS.n4205 585
R1193 VSS.n4175 VSS.n4173 585
R1194 VSS.n4284 VSS.n4175 585
R1195 VSS.n4153 VSS.n4152 585
R1196 VSS.n4285 VSS.n4152 585
R1197 VSS.n4161 VSS.n4151 585
R1198 VSS.n4316 VSS.n4151 585
R1199 VSS.n4282 VSS.n4281 585
R1200 VSS.n4283 VSS.n4282 585
R1201 VSS.n4251 VSS.n4185 585
R1202 VSS.n4252 VSS.n4251 585
R1203 VSS.n4246 VSS.n4204 585
R1204 VSS.n4250 VSS.n4204 585
R1205 VSS.n4182 VSS.n4181 585
R1206 VSS.n4286 VSS.n4182 585
R1207 VSS.n4318 VSS.n4150 585
R1208 VSS.n4318 VSS.n4317 585
R1209 VSS.n4225 VSS.n4224 585
R1210 VSS.n4224 VSS.n4223 585
R1211 VSS.n4731 VSS.n4720 585
R1212 VSS.n4733 VSS.n4720 585
R1213 VSS.n4719 VSS.n4718 585
R1214 VSS.n4938 VSS.n4719 585
R1215 VSS.n4958 VSS.n4957 585
R1216 VSS.n4959 VSS.n4958 585
R1217 VSS.n4686 VSS.n4685 585
R1218 VSS.n4685 VSS.n4684 585
R1219 VSS.n4993 VSS.n4992 585
R1220 VSS.n4992 VSS.t364 585
R1221 VSS.n5011 VSS.n5010 585
R1222 VSS.n5012 VSS.n5011 585
R1223 VSS.n4704 VSS.n4702 585
R1224 VSS.n4961 VSS.n4704 585
R1225 VSS.n4703 VSS.n4701 585
R1226 VSS.n4960 VSS.n4703 585
R1227 VSS.n4941 VSS.n4940 585
R1228 VSS.n4940 VSS.n4939 585
R1229 VSS.n4683 VSS.n4682 585
R1230 VSS.n4991 VSS.n4683 585
R1231 VSS.n4668 VSS.n4667 585
R1232 VSS.n5013 VSS.n4668 585
R1233 VSS.n4736 VSS.n4735 585
R1234 VSS.n4735 VSS.n4734 585
R1235 VSS.n5024 VSS.n5020 585
R1236 VSS.n5028 VSS.n5020 585
R1237 VSS.n5072 VSS.n5071 585
R1238 VSS.n5073 VSS.n5072 585
R1239 VSS.n4645 VSS.n4643 585
R1240 VSS.n5075 VSS.n4645 585
R1241 VSS.n5128 VSS.n5127 585
R1242 VSS.n5127 VSS.n5126 585
R1243 VSS.n4611 VSS.n4610 585
R1244 VSS.t399 VSS.n4611 585
R1245 VSS.n5170 VSS.n5169 585
R1246 VSS.n5171 VSS.n5170 585
R1247 VSS.n5168 VSS.n4598 585
R1248 VSS.n5172 VSS.n4598 585
R1249 VSS.n5148 VSS.n5147 585
R1250 VSS.n5147 VSS.n5146 585
R1251 VSS.n5129 VSS.n4613 585
R1252 VSS.n4613 VSS.n4612 585
R1253 VSS.n4648 VSS.n4647 585
R1254 VSS.n4647 VSS.n4646 585
R1255 VSS.n5078 VSS.n5077 585
R1256 VSS.n5077 VSS.n5076 585
R1257 VSS.n5173 VSS.n4599 585
R1258 VSS.n5015 VSS.n5014 585
R1259 VSS.n5026 VSS.n5025 585
R1260 VSS.n5027 VSS.n5026 585
R1261 VSS.n4812 VSS.n4811 585
R1262 VSS.n4814 VSS.n4812 585
R1263 VSS.n4840 VSS.n4839 585
R1264 VSS.n4841 VSS.n4840 585
R1265 VSS.n4797 VSS.n4795 585
R1266 VSS.n4845 VSS.n4797 585
R1267 VSS.n4767 VSS.n4765 585
R1268 VSS.n4876 VSS.n4767 585
R1269 VSS.n4745 VSS.n4744 585
R1270 VSS.n4877 VSS.n4744 585
R1271 VSS.n4753 VSS.n4743 585
R1272 VSS.n4908 VSS.n4743 585
R1273 VSS.n4874 VSS.n4873 585
R1274 VSS.n4875 VSS.n4874 585
R1275 VSS.n4843 VSS.n4777 585
R1276 VSS.n4844 VSS.n4843 585
R1277 VSS.n4838 VSS.n4796 585
R1278 VSS.n4842 VSS.n4796 585
R1279 VSS.n4774 VSS.n4773 585
R1280 VSS.n4878 VSS.n4774 585
R1281 VSS.n4910 VSS.n4742 585
R1282 VSS.n4910 VSS.n4909 585
R1283 VSS.n4817 VSS.n4816 585
R1284 VSS.n4816 VSS.n4815 585
R1285 VSS.n2599 VSS.n2598 585
R1286 VSS.n2598 VSS.n2597 585
R1287 VSS.n2622 VSS.n2621 585
R1288 VSS.n2623 VSS.n2622 585
R1289 VSS.n2628 VSS.n2591 585
R1290 VSS.n2591 VSS.n2590 585
R1291 VSS.n2636 VSS.n2587 585
R1292 VSS.n2587 VSS.n2586 585
R1293 VSS.n2651 VSS.n2650 585
R1294 VSS.n2650 VSS.t549 585
R1295 VSS.n2663 VSS.n2662 585
R1296 VSS.n2664 VSS.n2663 585
R1297 VSS.n2635 VSS.n2634 585
R1298 VSS.n2634 VSS.n2633 585
R1299 VSS.n2630 VSS.n2629 585
R1300 VSS.n2631 VSS.n2630 585
R1301 VSS.n2620 VSS.n2594 585
R1302 VSS.n2624 VSS.n2594 585
R1303 VSS.n2585 VSS.n2584 585
R1304 VSS.n2649 VSS.n2585 585
R1305 VSS.n2576 VSS.n2575 585
R1306 VSS.n2665 VSS.n2576 585
R1307 VSS.n2357 VSS.n2356 585
R1308 VSS.n2356 VSS.n2355 585
R1309 VSS.n2673 VSS.n2670 585
R1310 VSS.n5261 VSS.n2670 585
R1311 VSS.n2700 VSS.n2699 585
R1312 VSS.n5245 VSS.n2700 585
R1313 VSS.n5232 VSS.n5231 585
R1314 VSS.n5231 VSS.n5230 585
R1315 VSS.n2783 VSS.n2782 585
R1316 VSS.n2784 VSS.n2783 585
R1317 VSS.n2791 VSS.n2790 585
R1318 VSS.t505 VSS.n2791 585
R1319 VSS.n2772 VSS.n2770 585
R1320 VSS.n5194 VSS.n2772 585
R1321 VSS.n5192 VSS.n5191 585
R1322 VSS.n5193 VSS.n5192 585
R1323 VSS.n2789 VSS.n2771 585
R1324 VSS.n2792 VSS.n2771 585
R1325 VSS.n2786 VSS.n2753 585
R1326 VSS.n2786 VSS.n2785 585
R1327 VSS.n5248 VSS.n5247 585
R1328 VSS.n5247 VSS.n5246 585
R1329 VSS.n5233 VSS.n2702 585
R1330 VSS.n2702 VSS.n2701 585
R1331 VSS.n2800 VSS.n2799 585
R1332 VSS.n2667 VSS.n2666 585
R1333 VSS.n5259 VSS.n5258 585
R1334 VSS.n5260 VSS.n5259 585
R1335 VSS.n2433 VSS.n2432 585
R1336 VSS.n2435 VSS.n2433 585
R1337 VSS.n2461 VSS.n2460 585
R1338 VSS.n2462 VSS.n2461 585
R1339 VSS.n2418 VSS.n2416 585
R1340 VSS.n2466 VSS.n2418 585
R1341 VSS.n2388 VSS.n2386 585
R1342 VSS.n2497 VSS.n2388 585
R1343 VSS.n2366 VSS.n2365 585
R1344 VSS.n2498 VSS.n2365 585
R1345 VSS.n2374 VSS.n2364 585
R1346 VSS.n2529 VSS.n2364 585
R1347 VSS.n2495 VSS.n2494 585
R1348 VSS.n2496 VSS.n2495 585
R1349 VSS.n2464 VSS.n2398 585
R1350 VSS.n2465 VSS.n2464 585
R1351 VSS.n2459 VSS.n2417 585
R1352 VSS.n2463 VSS.n2417 585
R1353 VSS.n2395 VSS.n2394 585
R1354 VSS.n2499 VSS.n2395 585
R1355 VSS.n2531 VSS.n2363 585
R1356 VSS.n2531 VSS.n2530 585
R1357 VSS.n2438 VSS.n2437 585
R1358 VSS.n2437 VSS.n2436 585
R1359 VSS.n5560 VSS.n5559 585
R1360 VSS.n5559 VSS.n5558 585
R1361 VSS.n5583 VSS.n5582 585
R1362 VSS.n5584 VSS.n5583 585
R1363 VSS.n5589 VSS.n5552 585
R1364 VSS.n5552 VSS.n5551 585
R1365 VSS.n5597 VSS.n5548 585
R1366 VSS.n5548 VSS.n5547 585
R1367 VSS.n5612 VSS.n5611 585
R1368 VSS.n5611 VSS.t418 585
R1369 VSS.n5624 VSS.n5623 585
R1370 VSS.n5625 VSS.n5624 585
R1371 VSS.n5596 VSS.n5595 585
R1372 VSS.n5595 VSS.n5594 585
R1373 VSS.n5591 VSS.n5590 585
R1374 VSS.n5592 VSS.n5591 585
R1375 VSS.n5581 VSS.n5555 585
R1376 VSS.n5585 VSS.n5555 585
R1377 VSS.n5546 VSS.n5545 585
R1378 VSS.n5610 VSS.n5546 585
R1379 VSS.n5537 VSS.n5536 585
R1380 VSS.n5626 VSS.n5537 585
R1381 VSS.n5318 VSS.n5317 585
R1382 VSS.n5317 VSS.n5316 585
R1383 VSS.n5634 VSS.n5631 585
R1384 VSS.n5834 VSS.n5631 585
R1385 VSS.n5661 VSS.n5660 585
R1386 VSS.n5818 VSS.n5661 585
R1387 VSS.n5805 VSS.n5804 585
R1388 VSS.n5804 VSS.n5803 585
R1389 VSS.n5757 VSS.n5756 585
R1390 VSS.n5758 VSS.n5757 585
R1391 VSS.n5765 VSS.n5764 585
R1392 VSS.t17 VSS.n5765 585
R1393 VSS.n5746 VSS.n5744 585
R1394 VSS.n5767 VSS.n5746 585
R1395 VSS.n5743 VSS.n7 585
R1396 VSS.n9 VSS.n7 585
R1397 VSS.n5763 VSS.n5745 585
R1398 VSS.n5766 VSS.n5745 585
R1399 VSS.n5760 VSS.n5714 585
R1400 VSS.n5760 VSS.n5759 585
R1401 VSS.n5821 VSS.n5820 585
R1402 VSS.n5820 VSS.n5819 585
R1403 VSS.n5806 VSS.n5663 585
R1404 VSS.n5663 VSS.n5662 585
R1405 VSS.n18879 VSS.n8 585
R1406 VSS.n5628 VSS.n5627 585
R1407 VSS.n5832 VSS.n5831 585
R1408 VSS.n5833 VSS.n5832 585
R1409 VSS.n5394 VSS.n5393 585
R1410 VSS.n5396 VSS.n5394 585
R1411 VSS.n5422 VSS.n5421 585
R1412 VSS.n5423 VSS.n5422 585
R1413 VSS.n5379 VSS.n5377 585
R1414 VSS.n5427 VSS.n5379 585
R1415 VSS.n5349 VSS.n5347 585
R1416 VSS.n5458 VSS.n5349 585
R1417 VSS.n5327 VSS.n5326 585
R1418 VSS.n5459 VSS.n5326 585
R1419 VSS.n5335 VSS.n5325 585
R1420 VSS.n5490 VSS.n5325 585
R1421 VSS.n5456 VSS.n5455 585
R1422 VSS.n5457 VSS.n5456 585
R1423 VSS.n5425 VSS.n5359 585
R1424 VSS.n5426 VSS.n5425 585
R1425 VSS.n5420 VSS.n5378 585
R1426 VSS.n5424 VSS.n5378 585
R1427 VSS.n5356 VSS.n5355 585
R1428 VSS.n5460 VSS.n5356 585
R1429 VSS.n5492 VSS.n5324 585
R1430 VSS.n5492 VSS.n5491 585
R1431 VSS.n5399 VSS.n5398 585
R1432 VSS.n5398 VSS.n5397 585
R1433 VSS.n6133 VSS.n6132 585
R1434 VSS.n6132 VSS.n6131 585
R1435 VSS.n6156 VSS.n6155 585
R1436 VSS.n6157 VSS.n6156 585
R1437 VSS.n6162 VSS.n6125 585
R1438 VSS.n6125 VSS.n6124 585
R1439 VSS.n6170 VSS.n6121 585
R1440 VSS.n6121 VSS.n6120 585
R1441 VSS.n6185 VSS.n6184 585
R1442 VSS.n6184 VSS.t81 585
R1443 VSS.n6197 VSS.n6196 585
R1444 VSS.n6198 VSS.n6197 585
R1445 VSS.n6169 VSS.n6168 585
R1446 VSS.n6168 VSS.n6167 585
R1447 VSS.n6164 VSS.n6163 585
R1448 VSS.n6165 VSS.n6164 585
R1449 VSS.n6154 VSS.n6128 585
R1450 VSS.n6158 VSS.n6128 585
R1451 VSS.n6119 VSS.n6118 585
R1452 VSS.n6183 VSS.n6119 585
R1453 VSS.n6110 VSS.n6109 585
R1454 VSS.n6199 VSS.n6110 585
R1455 VSS.n5891 VSS.n5890 585
R1456 VSS.n5890 VSS.n5889 585
R1457 VSS.n6207 VSS.n6204 585
R1458 VSS.n6426 VSS.n6204 585
R1459 VSS.n6234 VSS.n6233 585
R1460 VSS.n6410 VSS.n6234 585
R1461 VSS.n6397 VSS.n6396 585
R1462 VSS.n6396 VSS.n6395 585
R1463 VSS.n6317 VSS.n6316 585
R1464 VSS.n6318 VSS.n6317 585
R1465 VSS.n6325 VSS.n6324 585
R1466 VSS.t31 VSS.n6325 585
R1467 VSS.n6306 VSS.n6304 585
R1468 VSS.n6359 VSS.n6306 585
R1469 VSS.n6357 VSS.n6356 585
R1470 VSS.n6358 VSS.n6357 585
R1471 VSS.n6323 VSS.n6305 585
R1472 VSS.n6326 VSS.n6305 585
R1473 VSS.n6320 VSS.n6287 585
R1474 VSS.n6320 VSS.n6319 585
R1475 VSS.n6413 VSS.n6412 585
R1476 VSS.n6412 VSS.n6411 585
R1477 VSS.n6398 VSS.n6236 585
R1478 VSS.n6236 VSS.n6235 585
R1479 VSS.n6334 VSS.n6333 585
R1480 VSS.n6201 VSS.n6200 585
R1481 VSS.n6424 VSS.n6423 585
R1482 VSS.n6425 VSS.n6424 585
R1483 VSS.n5967 VSS.n5966 585
R1484 VSS.n5969 VSS.n5967 585
R1485 VSS.n5995 VSS.n5994 585
R1486 VSS.n5996 VSS.n5995 585
R1487 VSS.n5952 VSS.n5950 585
R1488 VSS.n6000 VSS.n5952 585
R1489 VSS.n5922 VSS.n5920 585
R1490 VSS.n6031 VSS.n5922 585
R1491 VSS.n5900 VSS.n5899 585
R1492 VSS.n6032 VSS.n5899 585
R1493 VSS.n5908 VSS.n5898 585
R1494 VSS.n6063 VSS.n5898 585
R1495 VSS.n6029 VSS.n6028 585
R1496 VSS.n6030 VSS.n6029 585
R1497 VSS.n5998 VSS.n5932 585
R1498 VSS.n5999 VSS.n5998 585
R1499 VSS.n5993 VSS.n5951 585
R1500 VSS.n5997 VSS.n5951 585
R1501 VSS.n5929 VSS.n5928 585
R1502 VSS.n6033 VSS.n5929 585
R1503 VSS.n6065 VSS.n5897 585
R1504 VSS.n6065 VSS.n6064 585
R1505 VSS.n5972 VSS.n5971 585
R1506 VSS.n5971 VSS.n5970 585
R1507 VSS.n7688 VSS.n7677 585
R1508 VSS.n7690 VSS.n7677 585
R1509 VSS.n7676 VSS.n7675 585
R1510 VSS.n7895 VSS.n7676 585
R1511 VSS.n7915 VSS.n7914 585
R1512 VSS.n7916 VSS.n7915 585
R1513 VSS.n7643 VSS.n7642 585
R1514 VSS.n7642 VSS.n7641 585
R1515 VSS.n7950 VSS.n7949 585
R1516 VSS.n7949 VSS.t72 585
R1517 VSS.n7968 VSS.n7967 585
R1518 VSS.n7969 VSS.n7968 585
R1519 VSS.n7661 VSS.n7659 585
R1520 VSS.n7918 VSS.n7661 585
R1521 VSS.n7660 VSS.n7658 585
R1522 VSS.n7917 VSS.n7660 585
R1523 VSS.n7898 VSS.n7897 585
R1524 VSS.n7897 VSS.n7896 585
R1525 VSS.n7640 VSS.n7639 585
R1526 VSS.n7948 VSS.n7640 585
R1527 VSS.n7625 VSS.n7624 585
R1528 VSS.n7970 VSS.n7625 585
R1529 VSS.n7693 VSS.n7692 585
R1530 VSS.n7692 VSS.n7691 585
R1531 VSS.n7981 VSS.n7977 585
R1532 VSS.n7985 VSS.n7977 585
R1533 VSS.n8029 VSS.n8028 585
R1534 VSS.n8030 VSS.n8029 585
R1535 VSS.n7602 VSS.n7600 585
R1536 VSS.n8032 VSS.n7602 585
R1537 VSS.n8085 VSS.n8084 585
R1538 VSS.n8084 VSS.n8083 585
R1539 VSS.n7568 VSS.n7567 585
R1540 VSS.t361 VSS.n7568 585
R1541 VSS.n8127 VSS.n8126 585
R1542 VSS.n8128 VSS.n8127 585
R1543 VSS.n8125 VSS.n7555 585
R1544 VSS.n8129 VSS.n7555 585
R1545 VSS.n8105 VSS.n8104 585
R1546 VSS.n8104 VSS.n8103 585
R1547 VSS.n8086 VSS.n7570 585
R1548 VSS.n7570 VSS.n7569 585
R1549 VSS.n7605 VSS.n7604 585
R1550 VSS.n7604 VSS.n7603 585
R1551 VSS.n8035 VSS.n8034 585
R1552 VSS.n8034 VSS.n8033 585
R1553 VSS.n8130 VSS.n7556 585
R1554 VSS.n7972 VSS.n7971 585
R1555 VSS.n7983 VSS.n7982 585
R1556 VSS.n7984 VSS.n7983 585
R1557 VSS.n7769 VSS.n7768 585
R1558 VSS.n7771 VSS.n7769 585
R1559 VSS.n7797 VSS.n7796 585
R1560 VSS.n7798 VSS.n7797 585
R1561 VSS.n7754 VSS.n7752 585
R1562 VSS.n7802 VSS.n7754 585
R1563 VSS.n7724 VSS.n7722 585
R1564 VSS.n7833 VSS.n7724 585
R1565 VSS.n7702 VSS.n7701 585
R1566 VSS.n7834 VSS.n7701 585
R1567 VSS.n7710 VSS.n7700 585
R1568 VSS.n7865 VSS.n7700 585
R1569 VSS.n7831 VSS.n7830 585
R1570 VSS.n7832 VSS.n7831 585
R1571 VSS.n7800 VSS.n7734 585
R1572 VSS.n7801 VSS.n7800 585
R1573 VSS.n7795 VSS.n7753 585
R1574 VSS.n7799 VSS.n7753 585
R1575 VSS.n7731 VSS.n7730 585
R1576 VSS.n7835 VSS.n7731 585
R1577 VSS.n7867 VSS.n7699 585
R1578 VSS.n7867 VSS.n7866 585
R1579 VSS.n7774 VSS.n7773 585
R1580 VSS.n7773 VSS.n7772 585
R1581 VSS.n8280 VSS.n8269 585
R1582 VSS.n8282 VSS.n8269 585
R1583 VSS.n8268 VSS.n8267 585
R1584 VSS.n8487 VSS.n8268 585
R1585 VSS.n8507 VSS.n8506 585
R1586 VSS.n8508 VSS.n8507 585
R1587 VSS.n8235 VSS.n8234 585
R1588 VSS.n8234 VSS.n8233 585
R1589 VSS.n8542 VSS.n8541 585
R1590 VSS.n8541 VSS.t93 585
R1591 VSS.n8560 VSS.n8559 585
R1592 VSS.n8561 VSS.n8560 585
R1593 VSS.n8253 VSS.n8251 585
R1594 VSS.n8510 VSS.n8253 585
R1595 VSS.n8252 VSS.n8250 585
R1596 VSS.n8509 VSS.n8252 585
R1597 VSS.n8490 VSS.n8489 585
R1598 VSS.n8489 VSS.n8488 585
R1599 VSS.n8232 VSS.n8231 585
R1600 VSS.n8540 VSS.n8232 585
R1601 VSS.n8217 VSS.n8216 585
R1602 VSS.n8562 VSS.n8217 585
R1603 VSS.n8285 VSS.n8284 585
R1604 VSS.n8284 VSS.n8283 585
R1605 VSS.n8573 VSS.n8569 585
R1606 VSS.n8577 VSS.n8569 585
R1607 VSS.n8621 VSS.n8620 585
R1608 VSS.n8622 VSS.n8621 585
R1609 VSS.n8194 VSS.n8192 585
R1610 VSS.n8624 VSS.n8194 585
R1611 VSS.n8677 VSS.n8676 585
R1612 VSS.n8676 VSS.n8675 585
R1613 VSS.n8160 VSS.n8159 585
R1614 VSS.t494 VSS.n8160 585
R1615 VSS.n8719 VSS.n8718 585
R1616 VSS.n8720 VSS.n8719 585
R1617 VSS.n8717 VSS.n8147 585
R1618 VSS.n8721 VSS.n8147 585
R1619 VSS.n8697 VSS.n8696 585
R1620 VSS.n8696 VSS.n8695 585
R1621 VSS.n8678 VSS.n8162 585
R1622 VSS.n8162 VSS.n8161 585
R1623 VSS.n8197 VSS.n8196 585
R1624 VSS.n8196 VSS.n8195 585
R1625 VSS.n8627 VSS.n8626 585
R1626 VSS.n8626 VSS.n8625 585
R1627 VSS.n8722 VSS.n8148 585
R1628 VSS.n8564 VSS.n8563 585
R1629 VSS.n8575 VSS.n8574 585
R1630 VSS.n8576 VSS.n8575 585
R1631 VSS.n8361 VSS.n8360 585
R1632 VSS.n8363 VSS.n8361 585
R1633 VSS.n8389 VSS.n8388 585
R1634 VSS.n8390 VSS.n8389 585
R1635 VSS.n8346 VSS.n8344 585
R1636 VSS.n8394 VSS.n8346 585
R1637 VSS.n8316 VSS.n8314 585
R1638 VSS.n8425 VSS.n8316 585
R1639 VSS.n8294 VSS.n8293 585
R1640 VSS.n8426 VSS.n8293 585
R1641 VSS.n8302 VSS.n8292 585
R1642 VSS.n8457 VSS.n8292 585
R1643 VSS.n8423 VSS.n8422 585
R1644 VSS.n8424 VSS.n8423 585
R1645 VSS.n8392 VSS.n8326 585
R1646 VSS.n8393 VSS.n8392 585
R1647 VSS.n8387 VSS.n8345 585
R1648 VSS.n8391 VSS.n8345 585
R1649 VSS.n8323 VSS.n8322 585
R1650 VSS.n8427 VSS.n8323 585
R1651 VSS.n8459 VSS.n8291 585
R1652 VSS.n8459 VSS.n8458 585
R1653 VSS.n8366 VSS.n8365 585
R1654 VSS.n8365 VSS.n8364 585
R1655 VSS.n8872 VSS.n8861 585
R1656 VSS.n8874 VSS.n8861 585
R1657 VSS.n8860 VSS.n8859 585
R1658 VSS.n9079 VSS.n8860 585
R1659 VSS.n9099 VSS.n9098 585
R1660 VSS.n9100 VSS.n9099 585
R1661 VSS.n8827 VSS.n8826 585
R1662 VSS.n8826 VSS.n8825 585
R1663 VSS.n9134 VSS.n9133 585
R1664 VSS.n9133 VSS.t85 585
R1665 VSS.n9152 VSS.n9151 585
R1666 VSS.n9153 VSS.n9152 585
R1667 VSS.n8845 VSS.n8843 585
R1668 VSS.n9102 VSS.n8845 585
R1669 VSS.n8844 VSS.n8842 585
R1670 VSS.n9101 VSS.n8844 585
R1671 VSS.n9082 VSS.n9081 585
R1672 VSS.n9081 VSS.n9080 585
R1673 VSS.n8824 VSS.n8823 585
R1674 VSS.n9132 VSS.n8824 585
R1675 VSS.n8809 VSS.n8808 585
R1676 VSS.n9154 VSS.n8809 585
R1677 VSS.n8877 VSS.n8876 585
R1678 VSS.n8876 VSS.n8875 585
R1679 VSS.n9165 VSS.n9161 585
R1680 VSS.n9169 VSS.n9161 585
R1681 VSS.n9213 VSS.n9212 585
R1682 VSS.n9214 VSS.n9213 585
R1683 VSS.n8786 VSS.n8784 585
R1684 VSS.n9216 VSS.n8786 585
R1685 VSS.n9269 VSS.n9268 585
R1686 VSS.n9268 VSS.n9267 585
R1687 VSS.n8752 VSS.n8751 585
R1688 VSS.t406 VSS.n8752 585
R1689 VSS.n9311 VSS.n9310 585
R1690 VSS.n9312 VSS.n9311 585
R1691 VSS.n9309 VSS.n8739 585
R1692 VSS.n9313 VSS.n8739 585
R1693 VSS.n9289 VSS.n9288 585
R1694 VSS.n9288 VSS.n9287 585
R1695 VSS.n9270 VSS.n8754 585
R1696 VSS.n8754 VSS.n8753 585
R1697 VSS.n8789 VSS.n8788 585
R1698 VSS.n8788 VSS.n8787 585
R1699 VSS.n9219 VSS.n9218 585
R1700 VSS.n9218 VSS.n9217 585
R1701 VSS.n9314 VSS.n8740 585
R1702 VSS.n9156 VSS.n9155 585
R1703 VSS.n9167 VSS.n9166 585
R1704 VSS.n9168 VSS.n9167 585
R1705 VSS.n8953 VSS.n8952 585
R1706 VSS.n8955 VSS.n8953 585
R1707 VSS.n8981 VSS.n8980 585
R1708 VSS.n8982 VSS.n8981 585
R1709 VSS.n8938 VSS.n8936 585
R1710 VSS.n8986 VSS.n8938 585
R1711 VSS.n8908 VSS.n8906 585
R1712 VSS.n9017 VSS.n8908 585
R1713 VSS.n8886 VSS.n8885 585
R1714 VSS.n9018 VSS.n8885 585
R1715 VSS.n8894 VSS.n8884 585
R1716 VSS.n9049 VSS.n8884 585
R1717 VSS.n9015 VSS.n9014 585
R1718 VSS.n9016 VSS.n9015 585
R1719 VSS.n8984 VSS.n8918 585
R1720 VSS.n8985 VSS.n8984 585
R1721 VSS.n8979 VSS.n8937 585
R1722 VSS.n8983 VSS.n8937 585
R1723 VSS.n8915 VSS.n8914 585
R1724 VSS.n9019 VSS.n8915 585
R1725 VSS.n9051 VSS.n8883 585
R1726 VSS.n9051 VSS.n9050 585
R1727 VSS.n8958 VSS.n8957 585
R1728 VSS.n8957 VSS.n8956 585
R1729 VSS.n10056 VSS.n10045 585
R1730 VSS.n10058 VSS.n10045 585
R1731 VSS.n10044 VSS.n10043 585
R1732 VSS.n10263 VSS.n10044 585
R1733 VSS.n10283 VSS.n10282 585
R1734 VSS.n10284 VSS.n10283 585
R1735 VSS.n10011 VSS.n10010 585
R1736 VSS.n10010 VSS.n10009 585
R1737 VSS.n10318 VSS.n10317 585
R1738 VSS.n10317 VSS.t100 585
R1739 VSS.n10336 VSS.n10335 585
R1740 VSS.n10337 VSS.n10336 585
R1741 VSS.n10029 VSS.n10027 585
R1742 VSS.n10286 VSS.n10029 585
R1743 VSS.n10028 VSS.n10026 585
R1744 VSS.n10285 VSS.n10028 585
R1745 VSS.n10266 VSS.n10265 585
R1746 VSS.n10265 VSS.n10264 585
R1747 VSS.n10008 VSS.n10007 585
R1748 VSS.n10316 VSS.n10008 585
R1749 VSS.n9993 VSS.n9992 585
R1750 VSS.n10338 VSS.n9993 585
R1751 VSS.n10061 VSS.n10060 585
R1752 VSS.n10060 VSS.n10059 585
R1753 VSS.n10349 VSS.n10345 585
R1754 VSS.n10353 VSS.n10345 585
R1755 VSS.n10397 VSS.n10396 585
R1756 VSS.n10398 VSS.n10397 585
R1757 VSS.n9970 VSS.n9968 585
R1758 VSS.n10400 VSS.n9970 585
R1759 VSS.n10453 VSS.n10452 585
R1760 VSS.n10452 VSS.n10451 585
R1761 VSS.n9936 VSS.n9935 585
R1762 VSS.t378 VSS.n9936 585
R1763 VSS.n10495 VSS.n10494 585
R1764 VSS.n10496 VSS.n10495 585
R1765 VSS.n10493 VSS.n9923 585
R1766 VSS.n10497 VSS.n9923 585
R1767 VSS.n10473 VSS.n10472 585
R1768 VSS.n10472 VSS.n10471 585
R1769 VSS.n10454 VSS.n9938 585
R1770 VSS.n9938 VSS.n9937 585
R1771 VSS.n9973 VSS.n9972 585
R1772 VSS.n9972 VSS.n9971 585
R1773 VSS.n10403 VSS.n10402 585
R1774 VSS.n10402 VSS.n10401 585
R1775 VSS.n10498 VSS.n9924 585
R1776 VSS.n10340 VSS.n10339 585
R1777 VSS.n10351 VSS.n10350 585
R1778 VSS.n10352 VSS.n10351 585
R1779 VSS.n10137 VSS.n10136 585
R1780 VSS.n10139 VSS.n10137 585
R1781 VSS.n10165 VSS.n10164 585
R1782 VSS.n10166 VSS.n10165 585
R1783 VSS.n10122 VSS.n10120 585
R1784 VSS.n10170 VSS.n10122 585
R1785 VSS.n10092 VSS.n10090 585
R1786 VSS.n10201 VSS.n10092 585
R1787 VSS.n10070 VSS.n10069 585
R1788 VSS.n10202 VSS.n10069 585
R1789 VSS.n10078 VSS.n10068 585
R1790 VSS.n10233 VSS.n10068 585
R1791 VSS.n10199 VSS.n10198 585
R1792 VSS.n10200 VSS.n10199 585
R1793 VSS.n10168 VSS.n10102 585
R1794 VSS.n10169 VSS.n10168 585
R1795 VSS.n10163 VSS.n10121 585
R1796 VSS.n10167 VSS.n10121 585
R1797 VSS.n10099 VSS.n10098 585
R1798 VSS.n10203 VSS.n10099 585
R1799 VSS.n10235 VSS.n10067 585
R1800 VSS.n10235 VSS.n10234 585
R1801 VSS.n10142 VSS.n10141 585
R1802 VSS.n10141 VSS.n10140 585
R1803 VSS.n10648 VSS.n10637 585
R1804 VSS.n10650 VSS.n10637 585
R1805 VSS.n10636 VSS.n10635 585
R1806 VSS.n10855 VSS.n10636 585
R1807 VSS.n10875 VSS.n10874 585
R1808 VSS.n10876 VSS.n10875 585
R1809 VSS.n10603 VSS.n10602 585
R1810 VSS.n10602 VSS.n10601 585
R1811 VSS.n10910 VSS.n10909 585
R1812 VSS.n10909 VSS.t519 585
R1813 VSS.n10928 VSS.n10927 585
R1814 VSS.n10929 VSS.n10928 585
R1815 VSS.n10621 VSS.n10619 585
R1816 VSS.n10878 VSS.n10621 585
R1817 VSS.n10620 VSS.n10618 585
R1818 VSS.n10877 VSS.n10620 585
R1819 VSS.n10858 VSS.n10857 585
R1820 VSS.n10857 VSS.n10856 585
R1821 VSS.n10600 VSS.n10599 585
R1822 VSS.n10908 VSS.n10600 585
R1823 VSS.n10585 VSS.n10584 585
R1824 VSS.n10930 VSS.n10585 585
R1825 VSS.n10653 VSS.n10652 585
R1826 VSS.n10652 VSS.n10651 585
R1827 VSS.n10941 VSS.n10937 585
R1828 VSS.n10945 VSS.n10937 585
R1829 VSS.n10989 VSS.n10988 585
R1830 VSS.n10990 VSS.n10989 585
R1831 VSS.n10562 VSS.n10560 585
R1832 VSS.n10992 VSS.n10562 585
R1833 VSS.n11045 VSS.n11044 585
R1834 VSS.n11044 VSS.n11043 585
R1835 VSS.n10528 VSS.n10527 585
R1836 VSS.t164 VSS.n10528 585
R1837 VSS.n11087 VSS.n11086 585
R1838 VSS.n11088 VSS.n11087 585
R1839 VSS.n11085 VSS.n10515 585
R1840 VSS.n11089 VSS.n10515 585
R1841 VSS.n11065 VSS.n11064 585
R1842 VSS.n11064 VSS.n11063 585
R1843 VSS.n11046 VSS.n10530 585
R1844 VSS.n10530 VSS.n10529 585
R1845 VSS.n10565 VSS.n10564 585
R1846 VSS.n10564 VSS.n10563 585
R1847 VSS.n10995 VSS.n10994 585
R1848 VSS.n10994 VSS.n10993 585
R1849 VSS.n11090 VSS.n10516 585
R1850 VSS.n10932 VSS.n10931 585
R1851 VSS.n10943 VSS.n10942 585
R1852 VSS.n10944 VSS.n10943 585
R1853 VSS.n10729 VSS.n10728 585
R1854 VSS.n10731 VSS.n10729 585
R1855 VSS.n10757 VSS.n10756 585
R1856 VSS.n10758 VSS.n10757 585
R1857 VSS.n10714 VSS.n10712 585
R1858 VSS.n10762 VSS.n10714 585
R1859 VSS.n10684 VSS.n10682 585
R1860 VSS.n10793 VSS.n10684 585
R1861 VSS.n10662 VSS.n10661 585
R1862 VSS.n10794 VSS.n10661 585
R1863 VSS.n10670 VSS.n10660 585
R1864 VSS.n10825 VSS.n10660 585
R1865 VSS.n10791 VSS.n10790 585
R1866 VSS.n10792 VSS.n10791 585
R1867 VSS.n10760 VSS.n10694 585
R1868 VSS.n10761 VSS.n10760 585
R1869 VSS.n10755 VSS.n10713 585
R1870 VSS.n10759 VSS.n10713 585
R1871 VSS.n10691 VSS.n10690 585
R1872 VSS.n10795 VSS.n10691 585
R1873 VSS.n10827 VSS.n10659 585
R1874 VSS.n10827 VSS.n10826 585
R1875 VSS.n10734 VSS.n10733 585
R1876 VSS.n10733 VSS.n10732 585
R1877 VSS.n11240 VSS.n11229 585
R1878 VSS.n11242 VSS.n11229 585
R1879 VSS.n11228 VSS.n11227 585
R1880 VSS.n11447 VSS.n11228 585
R1881 VSS.n11467 VSS.n11466 585
R1882 VSS.n11468 VSS.n11467 585
R1883 VSS.n11195 VSS.n11194 585
R1884 VSS.n11194 VSS.n11193 585
R1885 VSS.n11502 VSS.n11501 585
R1886 VSS.n11501 VSS.t395 585
R1887 VSS.n11520 VSS.n11519 585
R1888 VSS.n11521 VSS.n11520 585
R1889 VSS.n11213 VSS.n11211 585
R1890 VSS.n11470 VSS.n11213 585
R1891 VSS.n11212 VSS.n11210 585
R1892 VSS.n11469 VSS.n11212 585
R1893 VSS.n11450 VSS.n11449 585
R1894 VSS.n11449 VSS.n11448 585
R1895 VSS.n11192 VSS.n11191 585
R1896 VSS.n11500 VSS.n11192 585
R1897 VSS.n11177 VSS.n11176 585
R1898 VSS.n11522 VSS.n11177 585
R1899 VSS.n11245 VSS.n11244 585
R1900 VSS.n11244 VSS.n11243 585
R1901 VSS.n11533 VSS.n11529 585
R1902 VSS.n11537 VSS.n11529 585
R1903 VSS.n11581 VSS.n11580 585
R1904 VSS.n11582 VSS.n11581 585
R1905 VSS.n11154 VSS.n11152 585
R1906 VSS.n11584 VSS.n11154 585
R1907 VSS.n11637 VSS.n11636 585
R1908 VSS.n11636 VSS.n11635 585
R1909 VSS.n11120 VSS.n11119 585
R1910 VSS.t58 VSS.n11120 585
R1911 VSS.n11679 VSS.n11678 585
R1912 VSS.n11680 VSS.n11679 585
R1913 VSS.n11677 VSS.n11107 585
R1914 VSS.n11681 VSS.n11107 585
R1915 VSS.n11657 VSS.n11656 585
R1916 VSS.n11656 VSS.n11655 585
R1917 VSS.n11638 VSS.n11122 585
R1918 VSS.n11122 VSS.n11121 585
R1919 VSS.n11157 VSS.n11156 585
R1920 VSS.n11156 VSS.n11155 585
R1921 VSS.n11587 VSS.n11586 585
R1922 VSS.n11586 VSS.n11585 585
R1923 VSS.n11682 VSS.n11108 585
R1924 VSS.n11524 VSS.n11523 585
R1925 VSS.n11535 VSS.n11534 585
R1926 VSS.n11536 VSS.n11535 585
R1927 VSS.n11321 VSS.n11320 585
R1928 VSS.n11323 VSS.n11321 585
R1929 VSS.n11349 VSS.n11348 585
R1930 VSS.n11350 VSS.n11349 585
R1931 VSS.n11306 VSS.n11304 585
R1932 VSS.n11354 VSS.n11306 585
R1933 VSS.n11276 VSS.n11274 585
R1934 VSS.n11385 VSS.n11276 585
R1935 VSS.n11254 VSS.n11253 585
R1936 VSS.n11386 VSS.n11253 585
R1937 VSS.n11262 VSS.n11252 585
R1938 VSS.n11417 VSS.n11252 585
R1939 VSS.n11383 VSS.n11382 585
R1940 VSS.n11384 VSS.n11383 585
R1941 VSS.n11352 VSS.n11286 585
R1942 VSS.n11353 VSS.n11352 585
R1943 VSS.n11347 VSS.n11305 585
R1944 VSS.n11351 VSS.n11305 585
R1945 VSS.n11283 VSS.n11282 585
R1946 VSS.n11387 VSS.n11283 585
R1947 VSS.n11419 VSS.n11251 585
R1948 VSS.n11419 VSS.n11418 585
R1949 VSS.n11326 VSS.n11325 585
R1950 VSS.n11325 VSS.n11324 585
R1951 VSS.n11832 VSS.n11821 585
R1952 VSS.n11834 VSS.n11821 585
R1953 VSS.n11820 VSS.n11819 585
R1954 VSS.n12039 VSS.n11820 585
R1955 VSS.n12059 VSS.n12058 585
R1956 VSS.n12060 VSS.n12059 585
R1957 VSS.n11787 VSS.n11786 585
R1958 VSS.n11786 VSS.n11785 585
R1959 VSS.n12094 VSS.n12093 585
R1960 VSS.n12093 VSS.t244 585
R1961 VSS.n12112 VSS.n12111 585
R1962 VSS.n12113 VSS.n12112 585
R1963 VSS.n11805 VSS.n11803 585
R1964 VSS.n12062 VSS.n11805 585
R1965 VSS.n11804 VSS.n11802 585
R1966 VSS.n12061 VSS.n11804 585
R1967 VSS.n12042 VSS.n12041 585
R1968 VSS.n12041 VSS.n12040 585
R1969 VSS.n11784 VSS.n11783 585
R1970 VSS.n12092 VSS.n11784 585
R1971 VSS.n11769 VSS.n11768 585
R1972 VSS.n12114 VSS.n11769 585
R1973 VSS.n11837 VSS.n11836 585
R1974 VSS.n11836 VSS.n11835 585
R1975 VSS.n12125 VSS.n12121 585
R1976 VSS.n12129 VSS.n12121 585
R1977 VSS.n12173 VSS.n12172 585
R1978 VSS.n12174 VSS.n12173 585
R1979 VSS.n11746 VSS.n11744 585
R1980 VSS.n12176 VSS.n11746 585
R1981 VSS.n12229 VSS.n12228 585
R1982 VSS.n12228 VSS.n12227 585
R1983 VSS.n11712 VSS.n11711 585
R1984 VSS.t259 VSS.n11712 585
R1985 VSS.n12271 VSS.n12270 585
R1986 VSS.n12272 VSS.n12271 585
R1987 VSS.n12269 VSS.n11699 585
R1988 VSS.n12273 VSS.n11699 585
R1989 VSS.n12249 VSS.n12248 585
R1990 VSS.n12248 VSS.n12247 585
R1991 VSS.n12230 VSS.n11714 585
R1992 VSS.n11714 VSS.n11713 585
R1993 VSS.n11749 VSS.n11748 585
R1994 VSS.n11748 VSS.n11747 585
R1995 VSS.n12179 VSS.n12178 585
R1996 VSS.n12178 VSS.n12177 585
R1997 VSS.n12274 VSS.n11700 585
R1998 VSS.n12116 VSS.n12115 585
R1999 VSS.n12127 VSS.n12126 585
R2000 VSS.n12128 VSS.n12127 585
R2001 VSS.n11913 VSS.n11912 585
R2002 VSS.n11915 VSS.n11913 585
R2003 VSS.n11941 VSS.n11940 585
R2004 VSS.n11942 VSS.n11941 585
R2005 VSS.n11898 VSS.n11896 585
R2006 VSS.n11946 VSS.n11898 585
R2007 VSS.n11868 VSS.n11866 585
R2008 VSS.n11977 VSS.n11868 585
R2009 VSS.n11846 VSS.n11845 585
R2010 VSS.n11978 VSS.n11845 585
R2011 VSS.n11854 VSS.n11844 585
R2012 VSS.n12009 VSS.n11844 585
R2013 VSS.n11975 VSS.n11974 585
R2014 VSS.n11976 VSS.n11975 585
R2015 VSS.n11944 VSS.n11878 585
R2016 VSS.n11945 VSS.n11944 585
R2017 VSS.n11939 VSS.n11897 585
R2018 VSS.n11943 VSS.n11897 585
R2019 VSS.n11875 VSS.n11874 585
R2020 VSS.n11979 VSS.n11875 585
R2021 VSS.n12011 VSS.n11843 585
R2022 VSS.n12011 VSS.n12010 585
R2023 VSS.n11918 VSS.n11917 585
R2024 VSS.n11917 VSS.n11916 585
R2025 VSS.n12424 VSS.n12413 585
R2026 VSS.n12426 VSS.n12413 585
R2027 VSS.n12412 VSS.n12411 585
R2028 VSS.n12631 VSS.n12412 585
R2029 VSS.n12651 VSS.n12650 585
R2030 VSS.n12652 VSS.n12651 585
R2031 VSS.n12379 VSS.n12378 585
R2032 VSS.n12378 VSS.n12377 585
R2033 VSS.n12686 VSS.n12685 585
R2034 VSS.n12685 VSS.t221 585
R2035 VSS.n12704 VSS.n12703 585
R2036 VSS.n12705 VSS.n12704 585
R2037 VSS.n12397 VSS.n12395 585
R2038 VSS.n12654 VSS.n12397 585
R2039 VSS.n12396 VSS.n12394 585
R2040 VSS.n12653 VSS.n12396 585
R2041 VSS.n12634 VSS.n12633 585
R2042 VSS.n12633 VSS.n12632 585
R2043 VSS.n12376 VSS.n12375 585
R2044 VSS.n12684 VSS.n12376 585
R2045 VSS.n12361 VSS.n12360 585
R2046 VSS.n12706 VSS.n12361 585
R2047 VSS.n12429 VSS.n12428 585
R2048 VSS.n12428 VSS.n12427 585
R2049 VSS.n12717 VSS.n12713 585
R2050 VSS.n12721 VSS.n12713 585
R2051 VSS.n12765 VSS.n12764 585
R2052 VSS.n12766 VSS.n12765 585
R2053 VSS.n12338 VSS.n12336 585
R2054 VSS.n12768 VSS.n12338 585
R2055 VSS.n12821 VSS.n12820 585
R2056 VSS.n12820 VSS.n12819 585
R2057 VSS.n12304 VSS.n12303 585
R2058 VSS.t441 VSS.n12304 585
R2059 VSS.n12863 VSS.n12862 585
R2060 VSS.n12864 VSS.n12863 585
R2061 VSS.n12861 VSS.n12291 585
R2062 VSS.n12865 VSS.n12291 585
R2063 VSS.n12841 VSS.n12840 585
R2064 VSS.n12840 VSS.n12839 585
R2065 VSS.n12822 VSS.n12306 585
R2066 VSS.n12306 VSS.n12305 585
R2067 VSS.n12341 VSS.n12340 585
R2068 VSS.n12340 VSS.n12339 585
R2069 VSS.n12771 VSS.n12770 585
R2070 VSS.n12770 VSS.n12769 585
R2071 VSS.n12866 VSS.n12292 585
R2072 VSS.n12708 VSS.n12707 585
R2073 VSS.n12719 VSS.n12718 585
R2074 VSS.n12720 VSS.n12719 585
R2075 VSS.n12505 VSS.n12504 585
R2076 VSS.n12507 VSS.n12505 585
R2077 VSS.n12533 VSS.n12532 585
R2078 VSS.n12534 VSS.n12533 585
R2079 VSS.n12490 VSS.n12488 585
R2080 VSS.n12538 VSS.n12490 585
R2081 VSS.n12460 VSS.n12458 585
R2082 VSS.n12569 VSS.n12460 585
R2083 VSS.n12438 VSS.n12437 585
R2084 VSS.n12570 VSS.n12437 585
R2085 VSS.n12446 VSS.n12436 585
R2086 VSS.n12601 VSS.n12436 585
R2087 VSS.n12567 VSS.n12566 585
R2088 VSS.n12568 VSS.n12567 585
R2089 VSS.n12536 VSS.n12470 585
R2090 VSS.n12537 VSS.n12536 585
R2091 VSS.n12531 VSS.n12489 585
R2092 VSS.n12535 VSS.n12489 585
R2093 VSS.n12467 VSS.n12466 585
R2094 VSS.n12571 VSS.n12467 585
R2095 VSS.n12603 VSS.n12435 585
R2096 VSS.n12603 VSS.n12602 585
R2097 VSS.n12510 VSS.n12509 585
R2098 VSS.n12509 VSS.n12508 585
R2099 VSS.n13016 VSS.n13005 585
R2100 VSS.n13018 VSS.n13005 585
R2101 VSS.n13004 VSS.n13003 585
R2102 VSS.n13223 VSS.n13004 585
R2103 VSS.n13243 VSS.n13242 585
R2104 VSS.n13244 VSS.n13243 585
R2105 VSS.n12971 VSS.n12970 585
R2106 VSS.n12970 VSS.n12969 585
R2107 VSS.n13278 VSS.n13277 585
R2108 VSS.n13277 VSS.t168 585
R2109 VSS.n13296 VSS.n13295 585
R2110 VSS.n13297 VSS.n13296 585
R2111 VSS.n12989 VSS.n12987 585
R2112 VSS.n13246 VSS.n12989 585
R2113 VSS.n12988 VSS.n12986 585
R2114 VSS.n13245 VSS.n12988 585
R2115 VSS.n13226 VSS.n13225 585
R2116 VSS.n13225 VSS.n13224 585
R2117 VSS.n12968 VSS.n12967 585
R2118 VSS.n13276 VSS.n12968 585
R2119 VSS.n12953 VSS.n12952 585
R2120 VSS.n13298 VSS.n12953 585
R2121 VSS.n13021 VSS.n13020 585
R2122 VSS.n13020 VSS.n13019 585
R2123 VSS.n13309 VSS.n13305 585
R2124 VSS.n13313 VSS.n13305 585
R2125 VSS.n13357 VSS.n13356 585
R2126 VSS.n13358 VSS.n13357 585
R2127 VSS.n12930 VSS.n12928 585
R2128 VSS.n13360 VSS.n12930 585
R2129 VSS.n13413 VSS.n13412 585
R2130 VSS.n13412 VSS.n13411 585
R2131 VSS.n12896 VSS.n12895 585
R2132 VSS.t3 VSS.n12896 585
R2133 VSS.n13455 VSS.n13454 585
R2134 VSS.n13456 VSS.n13455 585
R2135 VSS.n13453 VSS.n12883 585
R2136 VSS.n13457 VSS.n12883 585
R2137 VSS.n13433 VSS.n13432 585
R2138 VSS.n13432 VSS.n13431 585
R2139 VSS.n13414 VSS.n12898 585
R2140 VSS.n12898 VSS.n12897 585
R2141 VSS.n12933 VSS.n12932 585
R2142 VSS.n12932 VSS.n12931 585
R2143 VSS.n13363 VSS.n13362 585
R2144 VSS.n13362 VSS.n13361 585
R2145 VSS.n13458 VSS.n12884 585
R2146 VSS.n13300 VSS.n13299 585
R2147 VSS.n13311 VSS.n13310 585
R2148 VSS.n13312 VSS.n13311 585
R2149 VSS.n13097 VSS.n13096 585
R2150 VSS.n13099 VSS.n13097 585
R2151 VSS.n13125 VSS.n13124 585
R2152 VSS.n13126 VSS.n13125 585
R2153 VSS.n13082 VSS.n13080 585
R2154 VSS.n13130 VSS.n13082 585
R2155 VSS.n13052 VSS.n13050 585
R2156 VSS.n13161 VSS.n13052 585
R2157 VSS.n13030 VSS.n13029 585
R2158 VSS.n13162 VSS.n13029 585
R2159 VSS.n13038 VSS.n13028 585
R2160 VSS.n13193 VSS.n13028 585
R2161 VSS.n13159 VSS.n13158 585
R2162 VSS.n13160 VSS.n13159 585
R2163 VSS.n13128 VSS.n13062 585
R2164 VSS.n13129 VSS.n13128 585
R2165 VSS.n13123 VSS.n13081 585
R2166 VSS.n13127 VSS.n13081 585
R2167 VSS.n13059 VSS.n13058 585
R2168 VSS.n13163 VSS.n13059 585
R2169 VSS.n13195 VSS.n13027 585
R2170 VSS.n13195 VSS.n13194 585
R2171 VSS.n13102 VSS.n13101 585
R2172 VSS.n13101 VSS.n13100 585
R2173 VSS.n13608 VSS.n13597 585
R2174 VSS.n13610 VSS.n13597 585
R2175 VSS.n13596 VSS.n13595 585
R2176 VSS.n13815 VSS.n13596 585
R2177 VSS.n13835 VSS.n13834 585
R2178 VSS.n13836 VSS.n13835 585
R2179 VSS.n13563 VSS.n13562 585
R2180 VSS.n13562 VSS.n13561 585
R2181 VSS.n13870 VSS.n13869 585
R2182 VSS.n13869 VSS.t43 585
R2183 VSS.n13888 VSS.n13887 585
R2184 VSS.n13889 VSS.n13888 585
R2185 VSS.n13581 VSS.n13579 585
R2186 VSS.n13838 VSS.n13581 585
R2187 VSS.n13580 VSS.n13578 585
R2188 VSS.n13837 VSS.n13580 585
R2189 VSS.n13818 VSS.n13817 585
R2190 VSS.n13817 VSS.n13816 585
R2191 VSS.n13560 VSS.n13559 585
R2192 VSS.n13868 VSS.n13560 585
R2193 VSS.n13545 VSS.n13544 585
R2194 VSS.n13890 VSS.n13545 585
R2195 VSS.n13613 VSS.n13612 585
R2196 VSS.n13612 VSS.n13611 585
R2197 VSS.n13901 VSS.n13897 585
R2198 VSS.n13905 VSS.n13897 585
R2199 VSS.n13949 VSS.n13948 585
R2200 VSS.n13950 VSS.n13949 585
R2201 VSS.n13522 VSS.n13520 585
R2202 VSS.n13952 VSS.n13522 585
R2203 VSS.n14005 VSS.n14004 585
R2204 VSS.n14004 VSS.n14003 585
R2205 VSS.n13488 VSS.n13487 585
R2206 VSS.t460 VSS.n13488 585
R2207 VSS.n14047 VSS.n14046 585
R2208 VSS.n14048 VSS.n14047 585
R2209 VSS.n14045 VSS.n13475 585
R2210 VSS.n14049 VSS.n13475 585
R2211 VSS.n14025 VSS.n14024 585
R2212 VSS.n14024 VSS.n14023 585
R2213 VSS.n14006 VSS.n13490 585
R2214 VSS.n13490 VSS.n13489 585
R2215 VSS.n13525 VSS.n13524 585
R2216 VSS.n13524 VSS.n13523 585
R2217 VSS.n13955 VSS.n13954 585
R2218 VSS.n13954 VSS.n13953 585
R2219 VSS.n14050 VSS.n13476 585
R2220 VSS.n13892 VSS.n13891 585
R2221 VSS.n13903 VSS.n13902 585
R2222 VSS.n13904 VSS.n13903 585
R2223 VSS.n13689 VSS.n13688 585
R2224 VSS.n13691 VSS.n13689 585
R2225 VSS.n13717 VSS.n13716 585
R2226 VSS.n13718 VSS.n13717 585
R2227 VSS.n13674 VSS.n13672 585
R2228 VSS.n13722 VSS.n13674 585
R2229 VSS.n13644 VSS.n13642 585
R2230 VSS.n13753 VSS.n13644 585
R2231 VSS.n13622 VSS.n13621 585
R2232 VSS.n13754 VSS.n13621 585
R2233 VSS.n13630 VSS.n13620 585
R2234 VSS.n13785 VSS.n13620 585
R2235 VSS.n13751 VSS.n13750 585
R2236 VSS.n13752 VSS.n13751 585
R2237 VSS.n13720 VSS.n13654 585
R2238 VSS.n13721 VSS.n13720 585
R2239 VSS.n13715 VSS.n13673 585
R2240 VSS.n13719 VSS.n13673 585
R2241 VSS.n13651 VSS.n13650 585
R2242 VSS.n13755 VSS.n13651 585
R2243 VSS.n13787 VSS.n13619 585
R2244 VSS.n13787 VSS.n13786 585
R2245 VSS.n13694 VSS.n13693 585
R2246 VSS.n13693 VSS.n13692 585
R2247 VSS.n14200 VSS.n14189 585
R2248 VSS.n14202 VSS.n14189 585
R2249 VSS.n14188 VSS.n14187 585
R2250 VSS.n14407 VSS.n14188 585
R2251 VSS.n14427 VSS.n14426 585
R2252 VSS.n14428 VSS.n14427 585
R2253 VSS.n14155 VSS.n14154 585
R2254 VSS.n14154 VSS.n14153 585
R2255 VSS.n14462 VSS.n14461 585
R2256 VSS.n14461 VSS.t161 585
R2257 VSS.n14480 VSS.n14479 585
R2258 VSS.n14481 VSS.n14480 585
R2259 VSS.n14173 VSS.n14171 585
R2260 VSS.n14430 VSS.n14173 585
R2261 VSS.n14172 VSS.n14170 585
R2262 VSS.n14429 VSS.n14172 585
R2263 VSS.n14410 VSS.n14409 585
R2264 VSS.n14409 VSS.n14408 585
R2265 VSS.n14152 VSS.n14151 585
R2266 VSS.n14460 VSS.n14152 585
R2267 VSS.n14137 VSS.n14136 585
R2268 VSS.n14482 VSS.n14137 585
R2269 VSS.n14205 VSS.n14204 585
R2270 VSS.n14204 VSS.n14203 585
R2271 VSS.n14493 VSS.n14489 585
R2272 VSS.n14497 VSS.n14489 585
R2273 VSS.n14541 VSS.n14540 585
R2274 VSS.n14542 VSS.n14541 585
R2275 VSS.n14114 VSS.n14112 585
R2276 VSS.n14544 VSS.n14114 585
R2277 VSS.n14597 VSS.n14596 585
R2278 VSS.n14596 VSS.n14595 585
R2279 VSS.n14080 VSS.n14079 585
R2280 VSS.t39 VSS.n14080 585
R2281 VSS.n14639 VSS.n14638 585
R2282 VSS.n14640 VSS.n14639 585
R2283 VSS.n14637 VSS.n14067 585
R2284 VSS.n14641 VSS.n14067 585
R2285 VSS.n14617 VSS.n14616 585
R2286 VSS.n14616 VSS.n14615 585
R2287 VSS.n14598 VSS.n14082 585
R2288 VSS.n14082 VSS.n14081 585
R2289 VSS.n14117 VSS.n14116 585
R2290 VSS.n14116 VSS.n14115 585
R2291 VSS.n14547 VSS.n14546 585
R2292 VSS.n14546 VSS.n14545 585
R2293 VSS.n14642 VSS.n14068 585
R2294 VSS.n14484 VSS.n14483 585
R2295 VSS.n14495 VSS.n14494 585
R2296 VSS.n14496 VSS.n14495 585
R2297 VSS.n14281 VSS.n14280 585
R2298 VSS.n14283 VSS.n14281 585
R2299 VSS.n14309 VSS.n14308 585
R2300 VSS.n14310 VSS.n14309 585
R2301 VSS.n14266 VSS.n14264 585
R2302 VSS.n14314 VSS.n14266 585
R2303 VSS.n14236 VSS.n14234 585
R2304 VSS.n14345 VSS.n14236 585
R2305 VSS.n14214 VSS.n14213 585
R2306 VSS.n14346 VSS.n14213 585
R2307 VSS.n14222 VSS.n14212 585
R2308 VSS.n14377 VSS.n14212 585
R2309 VSS.n14343 VSS.n14342 585
R2310 VSS.n14344 VSS.n14343 585
R2311 VSS.n14312 VSS.n14246 585
R2312 VSS.n14313 VSS.n14312 585
R2313 VSS.n14307 VSS.n14265 585
R2314 VSS.n14311 VSS.n14265 585
R2315 VSS.n14243 VSS.n14242 585
R2316 VSS.n14347 VSS.n14243 585
R2317 VSS.n14379 VSS.n14211 585
R2318 VSS.n14379 VSS.n14378 585
R2319 VSS.n14286 VSS.n14285 585
R2320 VSS.n14285 VSS.n14284 585
R2321 VSS.n14792 VSS.n14781 585
R2322 VSS.n14794 VSS.n14781 585
R2323 VSS.n14780 VSS.n14779 585
R2324 VSS.n14999 VSS.n14780 585
R2325 VSS.n15019 VSS.n15018 585
R2326 VSS.n15020 VSS.n15019 585
R2327 VSS.n14747 VSS.n14746 585
R2328 VSS.n14746 VSS.n14745 585
R2329 VSS.n15054 VSS.n15053 585
R2330 VSS.n15053 VSS.t525 585
R2331 VSS.n15072 VSS.n15071 585
R2332 VSS.n15073 VSS.n15072 585
R2333 VSS.n14765 VSS.n14763 585
R2334 VSS.n15022 VSS.n14765 585
R2335 VSS.n14764 VSS.n14762 585
R2336 VSS.n15021 VSS.n14764 585
R2337 VSS.n15002 VSS.n15001 585
R2338 VSS.n15001 VSS.n15000 585
R2339 VSS.n14744 VSS.n14743 585
R2340 VSS.n15052 VSS.n14744 585
R2341 VSS.n14729 VSS.n14728 585
R2342 VSS.n15074 VSS.n14729 585
R2343 VSS.n14797 VSS.n14796 585
R2344 VSS.n14796 VSS.n14795 585
R2345 VSS.n15085 VSS.n15081 585
R2346 VSS.n15089 VSS.n15081 585
R2347 VSS.n15133 VSS.n15132 585
R2348 VSS.n15134 VSS.n15133 585
R2349 VSS.n14706 VSS.n14704 585
R2350 VSS.n15136 VSS.n14706 585
R2351 VSS.n15189 VSS.n15188 585
R2352 VSS.n15188 VSS.n15187 585
R2353 VSS.n14672 VSS.n14671 585
R2354 VSS.t152 VSS.n14672 585
R2355 VSS.n15231 VSS.n15230 585
R2356 VSS.n15232 VSS.n15231 585
R2357 VSS.n15229 VSS.n14659 585
R2358 VSS.n15233 VSS.n14659 585
R2359 VSS.n15209 VSS.n15208 585
R2360 VSS.n15208 VSS.n15207 585
R2361 VSS.n15190 VSS.n14674 585
R2362 VSS.n14674 VSS.n14673 585
R2363 VSS.n14709 VSS.n14708 585
R2364 VSS.n14708 VSS.n14707 585
R2365 VSS.n15139 VSS.n15138 585
R2366 VSS.n15138 VSS.n15137 585
R2367 VSS.n15234 VSS.n14660 585
R2368 VSS.n15076 VSS.n15075 585
R2369 VSS.n15087 VSS.n15086 585
R2370 VSS.n15088 VSS.n15087 585
R2371 VSS.n14873 VSS.n14872 585
R2372 VSS.n14875 VSS.n14873 585
R2373 VSS.n14901 VSS.n14900 585
R2374 VSS.n14902 VSS.n14901 585
R2375 VSS.n14858 VSS.n14856 585
R2376 VSS.n14906 VSS.n14858 585
R2377 VSS.n14828 VSS.n14826 585
R2378 VSS.n14937 VSS.n14828 585
R2379 VSS.n14806 VSS.n14805 585
R2380 VSS.n14938 VSS.n14805 585
R2381 VSS.n14814 VSS.n14804 585
R2382 VSS.n14969 VSS.n14804 585
R2383 VSS.n14935 VSS.n14934 585
R2384 VSS.n14936 VSS.n14935 585
R2385 VSS.n14904 VSS.n14838 585
R2386 VSS.n14905 VSS.n14904 585
R2387 VSS.n14899 VSS.n14857 585
R2388 VSS.n14903 VSS.n14857 585
R2389 VSS.n14835 VSS.n14834 585
R2390 VSS.n14939 VSS.n14835 585
R2391 VSS.n14971 VSS.n14803 585
R2392 VSS.n14971 VSS.n14970 585
R2393 VSS.n14878 VSS.n14877 585
R2394 VSS.n14877 VSS.n14876 585
R2395 VSS.n15384 VSS.n15373 585
R2396 VSS.n15386 VSS.n15373 585
R2397 VSS.n15372 VSS.n15371 585
R2398 VSS.n15591 VSS.n15372 585
R2399 VSS.n15611 VSS.n15610 585
R2400 VSS.n15612 VSS.n15611 585
R2401 VSS.n15339 VSS.n15338 585
R2402 VSS.n15338 VSS.n15337 585
R2403 VSS.n15646 VSS.n15645 585
R2404 VSS.n15645 VSS.t179 585
R2405 VSS.n15664 VSS.n15663 585
R2406 VSS.n15665 VSS.n15664 585
R2407 VSS.n15357 VSS.n15355 585
R2408 VSS.n15614 VSS.n15357 585
R2409 VSS.n15356 VSS.n15354 585
R2410 VSS.n15613 VSS.n15356 585
R2411 VSS.n15594 VSS.n15593 585
R2412 VSS.n15593 VSS.n15592 585
R2413 VSS.n15336 VSS.n15335 585
R2414 VSS.n15644 VSS.n15336 585
R2415 VSS.n15321 VSS.n15320 585
R2416 VSS.n15666 VSS.n15321 585
R2417 VSS.n15389 VSS.n15388 585
R2418 VSS.n15388 VSS.n15387 585
R2419 VSS.n15677 VSS.n15673 585
R2420 VSS.n15681 VSS.n15673 585
R2421 VSS.n15725 VSS.n15724 585
R2422 VSS.n15726 VSS.n15725 585
R2423 VSS.n15298 VSS.n15296 585
R2424 VSS.n15728 VSS.n15298 585
R2425 VSS.n15781 VSS.n15780 585
R2426 VSS.n15780 VSS.n15779 585
R2427 VSS.n15264 VSS.n15263 585
R2428 VSS.t374 VSS.n15264 585
R2429 VSS.n15823 VSS.n15822 585
R2430 VSS.n15824 VSS.n15823 585
R2431 VSS.n15821 VSS.n15251 585
R2432 VSS.n15825 VSS.n15251 585
R2433 VSS.n15801 VSS.n15800 585
R2434 VSS.n15800 VSS.n15799 585
R2435 VSS.n15782 VSS.n15266 585
R2436 VSS.n15266 VSS.n15265 585
R2437 VSS.n15301 VSS.n15300 585
R2438 VSS.n15300 VSS.n15299 585
R2439 VSS.n15731 VSS.n15730 585
R2440 VSS.n15730 VSS.n15729 585
R2441 VSS.n15826 VSS.n15252 585
R2442 VSS.n15668 VSS.n15667 585
R2443 VSS.n15679 VSS.n15678 585
R2444 VSS.n15680 VSS.n15679 585
R2445 VSS.n15465 VSS.n15464 585
R2446 VSS.n15467 VSS.n15465 585
R2447 VSS.n15493 VSS.n15492 585
R2448 VSS.n15494 VSS.n15493 585
R2449 VSS.n15450 VSS.n15448 585
R2450 VSS.n15498 VSS.n15450 585
R2451 VSS.n15420 VSS.n15418 585
R2452 VSS.n15529 VSS.n15420 585
R2453 VSS.n15398 VSS.n15397 585
R2454 VSS.n15530 VSS.n15397 585
R2455 VSS.n15406 VSS.n15396 585
R2456 VSS.n15561 VSS.n15396 585
R2457 VSS.n15527 VSS.n15526 585
R2458 VSS.n15528 VSS.n15527 585
R2459 VSS.n15496 VSS.n15430 585
R2460 VSS.n15497 VSS.n15496 585
R2461 VSS.n15491 VSS.n15449 585
R2462 VSS.n15495 VSS.n15449 585
R2463 VSS.n15427 VSS.n15426 585
R2464 VSS.n15531 VSS.n15427 585
R2465 VSS.n15563 VSS.n15395 585
R2466 VSS.n15563 VSS.n15562 585
R2467 VSS.n15470 VSS.n15469 585
R2468 VSS.n15469 VSS.n15468 585
R2469 VSS.n6739 VSS.n6738 585
R2470 VSS.n6738 VSS.n6737 585
R2471 VSS.n6762 VSS.n6761 585
R2472 VSS.n6763 VSS.n6762 585
R2473 VSS.n6768 VSS.n6731 585
R2474 VSS.n6731 VSS.n6730 585
R2475 VSS.n6776 VSS.n6727 585
R2476 VSS.n6727 VSS.n6726 585
R2477 VSS.n6791 VSS.n6790 585
R2478 VSS.n6790 VSS.t413 585
R2479 VSS.n6803 VSS.n6802 585
R2480 VSS.n6804 VSS.n6803 585
R2481 VSS.n6775 VSS.n6774 585
R2482 VSS.n6774 VSS.n6773 585
R2483 VSS.n6770 VSS.n6769 585
R2484 VSS.n6771 VSS.n6770 585
R2485 VSS.n6760 VSS.n6734 585
R2486 VSS.n6764 VSS.n6734 585
R2487 VSS.n6725 VSS.n6724 585
R2488 VSS.n6789 VSS.n6725 585
R2489 VSS.n6716 VSS.n6715 585
R2490 VSS.n6805 VSS.n6716 585
R2491 VSS.n6497 VSS.n6496 585
R2492 VSS.n6496 VSS.n6495 585
R2493 VSS.n6813 VSS.n6810 585
R2494 VSS.n15914 VSS.n6810 585
R2495 VSS.n6840 VSS.n6839 585
R2496 VSS.n15898 VSS.n6840 585
R2497 VSS.n15885 VSS.n15884 585
R2498 VSS.n15884 VSS.n15883 585
R2499 VSS.n6923 VSS.n6922 585
R2500 VSS.n6924 VSS.n6923 585
R2501 VSS.n6931 VSS.n6930 585
R2502 VSS.t113 VSS.n6931 585
R2503 VSS.n6912 VSS.n6910 585
R2504 VSS.n15847 VSS.n6912 585
R2505 VSS.n15845 VSS.n15844 585
R2506 VSS.n15846 VSS.n15845 585
R2507 VSS.n6929 VSS.n6911 585
R2508 VSS.n6932 VSS.n6911 585
R2509 VSS.n6926 VSS.n6893 585
R2510 VSS.n6926 VSS.n6925 585
R2511 VSS.n15901 VSS.n15900 585
R2512 VSS.n15900 VSS.n15899 585
R2513 VSS.n15886 VSS.n6842 585
R2514 VSS.n6842 VSS.n6841 585
R2515 VSS.n6940 VSS.n6939 585
R2516 VSS.n6807 VSS.n6806 585
R2517 VSS.n15912 VSS.n15911 585
R2518 VSS.n15913 VSS.n15912 585
R2519 VSS.n6573 VSS.n6572 585
R2520 VSS.n6575 VSS.n6573 585
R2521 VSS.n6601 VSS.n6600 585
R2522 VSS.n6602 VSS.n6601 585
R2523 VSS.n6558 VSS.n6556 585
R2524 VSS.n6606 VSS.n6558 585
R2525 VSS.n6528 VSS.n6526 585
R2526 VSS.n6637 VSS.n6528 585
R2527 VSS.n6506 VSS.n6505 585
R2528 VSS.n6638 VSS.n6505 585
R2529 VSS.n6514 VSS.n6504 585
R2530 VSS.n6669 VSS.n6504 585
R2531 VSS.n6635 VSS.n6634 585
R2532 VSS.n6636 VSS.n6635 585
R2533 VSS.n6604 VSS.n6538 585
R2534 VSS.n6605 VSS.n6604 585
R2535 VSS.n6599 VSS.n6557 585
R2536 VSS.n6603 VSS.n6557 585
R2537 VSS.n6535 VSS.n6534 585
R2538 VSS.n6639 VSS.n6535 585
R2539 VSS.n6671 VSS.n6503 585
R2540 VSS.n6671 VSS.n6670 585
R2541 VSS.n6578 VSS.n6577 585
R2542 VSS.n6577 VSS.n6576 585
R2543 VSS.n7095 VSS.n7084 585
R2544 VSS.n7097 VSS.n7084 585
R2545 VSS.n7083 VSS.n7082 585
R2546 VSS.n7303 VSS.n7083 585
R2547 VSS.n7323 VSS.n7322 585
R2548 VSS.n7324 VSS.n7323 585
R2549 VSS.n7050 VSS.n7049 585
R2550 VSS.n7049 VSS.n7048 585
R2551 VSS.n7358 VSS.n7357 585
R2552 VSS.n7357 VSS.t385 585
R2553 VSS.n7376 VSS.n7375 585
R2554 VSS.n7377 VSS.n7376 585
R2555 VSS.n7068 VSS.n7066 585
R2556 VSS.n7326 VSS.n7068 585
R2557 VSS.n7067 VSS.n7065 585
R2558 VSS.n7325 VSS.n7067 585
R2559 VSS.n7306 VSS.n7305 585
R2560 VSS.n7305 VSS.n7304 585
R2561 VSS.n7047 VSS.n7046 585
R2562 VSS.n7356 VSS.n7047 585
R2563 VSS.n7032 VSS.n7031 585
R2564 VSS.n7378 VSS.n7032 585
R2565 VSS.n7100 VSS.n7099 585
R2566 VSS.n7099 VSS.n7098 585
R2567 VSS.n7389 VSS.n7385 585
R2568 VSS.n7393 VSS.n7385 585
R2569 VSS.n7437 VSS.n7436 585
R2570 VSS.n7438 VSS.n7437 585
R2571 VSS.n7009 VSS.n7007 585
R2572 VSS.n7440 VSS.n7009 585
R2573 VSS.n7493 VSS.n7492 585
R2574 VSS.n7492 VSS.n7491 585
R2575 VSS.n6975 VSS.n6974 585
R2576 VSS.t437 VSS.n6975 585
R2577 VSS.n7535 VSS.n7534 585
R2578 VSS.n7536 VSS.n7535 585
R2579 VSS.n7533 VSS.n6962 585
R2580 VSS.n7537 VSS.n6962 585
R2581 VSS.n7513 VSS.n7512 585
R2582 VSS.n7512 VSS.n7511 585
R2583 VSS.n7494 VSS.n6977 585
R2584 VSS.n6977 VSS.n6976 585
R2585 VSS.n7012 VSS.n7011 585
R2586 VSS.n7011 VSS.n7010 585
R2587 VSS.n7443 VSS.n7442 585
R2588 VSS.n7442 VSS.n7441 585
R2589 VSS.n7538 VSS.n6963 585
R2590 VSS.n7380 VSS.n7379 585
R2591 VSS.n7391 VSS.n7390 585
R2592 VSS.n7392 VSS.n7391 585
R2593 VSS.n7170 VSS.n7159 585
R2594 VSS.n7172 VSS.n7159 585
R2595 VSS.n7158 VSS.n7157 585
R2596 VSS.n7198 VSS.n7158 585
R2597 VSS.n7218 VSS.n7217 585
R2598 VSS.n7219 VSS.n7218 585
R2599 VSS.n7125 VSS.n7124 585
R2600 VSS.n7124 VSS.n7123 585
R2601 VSS.n7254 VSS.n7253 585
R2602 VSS.n7253 VSS.n7252 585
R2603 VSS.n7272 VSS.n7271 585
R2604 VSS.n7273 VSS.n7272 585
R2605 VSS.n7145 VSS.n7143 585
R2606 VSS.n7221 VSS.n7145 585
R2607 VSS.n7144 VSS.n7142 585
R2608 VSS.n7220 VSS.n7144 585
R2609 VSS.n7201 VSS.n7200 585
R2610 VSS.n7200 VSS.n7199 585
R2611 VSS.n7122 VSS.n7121 585
R2612 VSS.n7251 VSS.n7122 585
R2613 VSS.n7107 VSS.n7106 585
R2614 VSS.n7274 VSS.n7107 585
R2615 VSS.n7175 VSS.n7174 585
R2616 VSS.n7174 VSS.n7173 585
R2617 VSS.n202 VSS.n182 585
R2618 VSS.n200 VSS.n182 585
R2619 VSS.n181 VSS.n180 585
R2620 VSS.n18615 VSS.n181 585
R2621 VSS.n18635 VSS.n18634 585
R2622 VSS.n18636 VSS.n18635 585
R2623 VSS.n148 VSS.n147 585
R2624 VSS.n147 VSS.n146 585
R2625 VSS.n18670 VSS.n18669 585
R2626 VSS.n18669 VSS.t129 585
R2627 VSS.n18688 VSS.n18687 585
R2628 VSS.n18689 VSS.n18688 585
R2629 VSS.n166 VSS.n164 585
R2630 VSS.n18638 VSS.n166 585
R2631 VSS.n165 VSS.n163 585
R2632 VSS.n18637 VSS.n165 585
R2633 VSS.n18618 VSS.n18617 585
R2634 VSS.n18617 VSS.n18616 585
R2635 VSS.n145 VSS.n144 585
R2636 VSS.n18668 VSS.n145 585
R2637 VSS.n130 VSS.n129 585
R2638 VSS.n18690 VSS.n130 585
R2639 VSS.n204 VSS.n203 585
R2640 VSS.n204 VSS.n201 585
R2641 VSS.n18701 VSS.n18697 585
R2642 VSS.n18705 VSS.n18697 585
R2643 VSS.n18749 VSS.n18748 585
R2644 VSS.n18750 VSS.n18749 585
R2645 VSS.n107 VSS.n105 585
R2646 VSS.n18752 VSS.n107 585
R2647 VSS.n18805 VSS.n18804 585
R2648 VSS.n18804 VSS.n18803 585
R2649 VSS.n73 VSS.n72 585
R2650 VSS.t182 VSS.n73 585
R2651 VSS.n18847 VSS.n18846 585
R2652 VSS.n18848 VSS.n18847 585
R2653 VSS.n18845 VSS.n60 585
R2654 VSS.n18849 VSS.n60 585
R2655 VSS.n18825 VSS.n18824 585
R2656 VSS.n18824 VSS.n18823 585
R2657 VSS.n18806 VSS.n75 585
R2658 VSS.n75 VSS.n74 585
R2659 VSS.n110 VSS.n109 585
R2660 VSS.n109 VSS.n108 585
R2661 VSS.n18755 VSS.n18754 585
R2662 VSS.n18754 VSS.n18753 585
R2663 VSS.n18850 VSS.n61 585
R2664 VSS.n18692 VSS.n18691 585
R2665 VSS.n18703 VSS.n18702 585
R2666 VSS.n18704 VSS.n18703 585
R2667 VSS.n358 VSS.n357 585
R2668 VSS.n359 VSS.n358 585
R2669 VSS.n363 VSS.n362 585
R2670 VSS.n362 VSS.n361 585
R2671 VSS.n339 VSS.n338 585
R2672 VSS.n374 VSS.n339 585
R2673 VSS.n335 VSS.n334 585
R2674 VSS.n383 VSS.n335 585
R2675 VSS.n398 VSS.n397 585
R2676 VSS.n399 VSS.n398 585
R2677 VSS.n403 VSS.n402 585
R2678 VSS.n402 VSS.n401 585
R2679 VSS.n381 VSS.n380 585
R2680 VSS.n382 VSS.n381 585
R2681 VSS.n377 VSS.n376 585
R2682 VSS.n376 VSS.n375 585
R2683 VSS.n364 VSS.n341 585
R2684 VSS.n341 VSS.n340 585
R2685 VSS.n394 VSS.n331 585
R2686 VSS.n331 VSS.n330 585
R2687 VSS.n198 VSS.n197 585
R2688 VSS.n199 VSS.n198 585
R2689 VSS.n290 VSS.n289 585
R2690 VSS.n289 VSS.n288 585
R2691 VSS.n18238 VSS.n18237 585
R2692 VSS.n18237 VSS.n18236 585
R2693 VSS.n18261 VSS.n18260 585
R2694 VSS.n18262 VSS.n18261 585
R2695 VSS.n18267 VSS.n18230 585
R2696 VSS.n18230 VSS.n18229 585
R2697 VSS.n18275 VSS.n18226 585
R2698 VSS.n18226 VSS.n18225 585
R2699 VSS.n18290 VSS.n18289 585
R2700 VSS.n18289 VSS.t69 585
R2701 VSS.n18302 VSS.n18301 585
R2702 VSS.n18303 VSS.n18302 585
R2703 VSS.n18274 VSS.n18273 585
R2704 VSS.n18273 VSS.n18272 585
R2705 VSS.n18269 VSS.n18268 585
R2706 VSS.n18270 VSS.n18269 585
R2707 VSS.n18259 VSS.n18233 585
R2708 VSS.n18263 VSS.n18233 585
R2709 VSS.n18224 VSS.n18223 585
R2710 VSS.n18288 VSS.n18224 585
R2711 VSS.n18215 VSS.n18214 585
R2712 VSS.n18304 VSS.n18215 585
R2713 VSS.n211 VSS.n210 585
R2714 VSS.n210 VSS.n209 585
R2715 VSS.n18312 VSS.n18309 585
R2716 VSS.n18531 VSS.n18309 585
R2717 VSS.n18366 VSS.n18362 585
R2718 VSS.n18370 VSS.n18362 585
R2719 VSS.n18381 VSS.n18380 585
R2720 VSS.n18382 VSS.n18381 585
R2721 VSS.n18493 VSS.n18492 585
R2722 VSS.n18494 VSS.n18493 585
R2723 VSS.n18442 VSS.n18440 585
R2724 VSS.t349 VSS.n18440 585
R2725 VSS.n18456 VSS.n18455 585
R2726 VSS.n18457 VSS.n18456 585
R2727 VSS.n18454 VSS.n18437 585
R2728 VSS.n18458 VSS.n18437 585
R2729 VSS.n18452 VSS.n18420 585
R2730 VSS.n18452 VSS.n18451 585
R2731 VSS.n18491 VSS.n18385 585
R2732 VSS.n18385 VSS.n18384 585
R2733 VSS.n18368 VSS.n18367 585
R2734 VSS.n18369 VSS.n18368 585
R2735 VSS.n18373 VSS.n18344 585
R2736 VSS.n18373 VSS.n18361 585
R2737 VSS.n18459 VSS.n18438 585
R2738 VSS.n18306 VSS.n18305 585
R2739 VSS.n18529 VSS.n18528 585
R2740 VSS.n18530 VSS.n18529 585
R2741 VSS.n564 VSS.n563 585
R2742 VSS.n563 VSS.n562 585
R2743 VSS.n585 VSS.n584 585
R2744 VSS.n586 VSS.n585 585
R2745 VSS.n591 VSS.n551 585
R2746 VSS.n551 VSS.n550 585
R2747 VSS.n599 VSS.n547 585
R2748 VSS.n547 VSS.n546 585
R2749 VSS.n614 VSS.n613 585
R2750 VSS.n613 VSS.t126 585
R2751 VSS.n626 VSS.n625 585
R2752 VSS.n627 VSS.n626 585
R2753 VSS.n598 VSS.n597 585
R2754 VSS.n597 VSS.n596 585
R2755 VSS.n593 VSS.n592 585
R2756 VSS.n594 VSS.n593 585
R2757 VSS.n583 VSS.n554 585
R2758 VSS.n587 VSS.n554 585
R2759 VSS.n545 VSS.n544 585
R2760 VSS.n612 VSS.n545 585
R2761 VSS.n536 VSS.n535 585
R2762 VSS.n628 VSS.n536 585
R2763 VSS.n558 VSS.n557 585
R2764 VSS.n561 VSS.n558 585
R2765 VSS.n762 VSS.n761 585
R2766 VSS.n761 VSS.n760 585
R2767 VSS.n800 VSS.n665 585
R2768 VSS.n665 VSS.n664 585
R2769 VSS.n799 VSS.n798 585
R2770 VSS.n798 VSS.n797 585
R2771 VSS.n815 VSS.n814 585
R2772 VSS.n814 VSS.n813 585
R2773 VSS.n630 VSS.n629 585
R2774 VSS.n636 VSS.n633 585
R2775 VSS.n828 VSS.n633 585
R2776 VSS.n826 VSS.n825 585
R2777 VSS.n827 VSS.n826 585
R2778 VSS.n663 VSS.n662 585
R2779 VSS.n812 VSS.n663 585
R2780 VSS.n757 VSS.n716 585
R2781 VSS.n757 VSS.n745 585
R2782 VSS.n756 VSS.n754 585
R2783 VSS.n756 VSS.n755 585
R2784 VSS.n744 VSS.n743 585
R2785 VSS.t335 VSS.n744 585
R2786 VSS.n18867 VSS.n45 585
R2787 VSS.n18871 VSS.n45 585
R2788 VSS.n18869 VSS.n18868 585
R2789 VSS.n18870 VSS.n18869 585
R2790 VSS.n42 VSS.n41 585
R2791 VSS.n907 VSS.n906 585
R2792 VSS.n906 VSS.n905 585
R2793 VSS.n928 VSS.n927 585
R2794 VSS.n929 VSS.n928 585
R2795 VSS.n934 VSS.n899 585
R2796 VSS.n899 VSS.n898 585
R2797 VSS.n942 VSS.n894 585
R2798 VSS.n894 VSS.n893 585
R2799 VSS.n958 VSS.n957 585
R2800 VSS.n957 VSS.n956 585
R2801 VSS.n970 VSS.n969 585
R2802 VSS.n971 VSS.n970 585
R2803 VSS.n941 VSS.n940 585
R2804 VSS.n940 VSS.n939 585
R2805 VSS.n936 VSS.n935 585
R2806 VSS.n937 VSS.n936 585
R2807 VSS.n926 VSS.n902 585
R2808 VSS.n930 VSS.n902 585
R2809 VSS.n892 VSS.n891 585
R2810 VSS.n955 VSS.n892 585
R2811 VSS.n883 VSS.n882 585
R2812 VSS.n972 VSS.n883 585
R2813 VSS.n456 VSS.n455 585
R2814 VSS.n455 VSS.n454 585
R2815 VSS.n1088 VSS.n1087 585
R2816 VSS.n1087 VSS.n1086 585
R2817 VSS.n1109 VSS.n1108 585
R2818 VSS.n1110 VSS.n1109 585
R2819 VSS.n1115 VSS.n1080 585
R2820 VSS.n1080 VSS.n1079 585
R2821 VSS.n1123 VSS.n1075 585
R2822 VSS.n1075 VSS.n1074 585
R2823 VSS.n1139 VSS.n1138 585
R2824 VSS.n1138 VSS.n1137 585
R2825 VSS.n1151 VSS.n1150 585
R2826 VSS.n1152 VSS.n1151 585
R2827 VSS.n1122 VSS.n1121 585
R2828 VSS.n1121 VSS.n1120 585
R2829 VSS.n1117 VSS.n1116 585
R2830 VSS.n1118 VSS.n1117 585
R2831 VSS.n1107 VSS.n1083 585
R2832 VSS.n1111 VSS.n1083 585
R2833 VSS.n1073 VSS.n1072 585
R2834 VSS.n1136 VSS.n1073 585
R2835 VSS.n1064 VSS.n1063 585
R2836 VSS.n1153 VSS.n1064 585
R2837 VSS.n1023 VSS.n1022 585
R2838 VSS.n1022 VSS.n1021 585
R2839 VSS.n17495 VSS.n17494 585
R2840 VSS.n17497 VSS.n17495 585
R2841 VSS.n17523 VSS.n17522 585
R2842 VSS.n17524 VSS.n17523 585
R2843 VSS.n17480 VSS.n17478 585
R2844 VSS.n17528 VSS.n17480 585
R2845 VSS.n17450 VSS.n17448 585
R2846 VSS.n17559 VSS.n17450 585
R2847 VSS.n17428 VSS.n17427 585
R2848 VSS.n17560 VSS.n17427 585
R2849 VSS.n17436 VSS.n17426 585
R2850 VSS.n17591 VSS.n17426 585
R2851 VSS.n17557 VSS.n17556 585
R2852 VSS.n17558 VSS.n17557 585
R2853 VSS.n17526 VSS.n17460 585
R2854 VSS.n17527 VSS.n17526 585
R2855 VSS.n17521 VSS.n17479 585
R2856 VSS.n17525 VSS.n17479 585
R2857 VSS.n17457 VSS.n17456 585
R2858 VSS.n17561 VSS.n17457 585
R2859 VSS.n17593 VSS.n17425 585
R2860 VSS.n17593 VSS.n17592 585
R2861 VSS.n17500 VSS.n17499 585
R2862 VSS.n17499 VSS.n17498 585
R2863 VSS.n1221 VSS.n1220 585
R2864 VSS.n1220 VSS.n1219 585
R2865 VSS.n1244 VSS.n1243 585
R2866 VSS.n1245 VSS.n1244 585
R2867 VSS.n1250 VSS.n1213 585
R2868 VSS.n1213 VSS.n1212 585
R2869 VSS.n1258 VSS.n1209 585
R2870 VSS.n1209 VSS.n1208 585
R2871 VSS.n1273 VSS.n1272 585
R2872 VSS.n1272 VSS.t584 585
R2873 VSS.n1285 VSS.n1284 585
R2874 VSS.n1286 VSS.n1285 585
R2875 VSS.n1257 VSS.n1256 585
R2876 VSS.n1256 VSS.n1255 585
R2877 VSS.n1252 VSS.n1251 585
R2878 VSS.n1253 VSS.n1252 585
R2879 VSS.n1242 VSS.n1216 585
R2880 VSS.n1246 VSS.n1216 585
R2881 VSS.n1207 VSS.n1206 585
R2882 VSS.n1271 VSS.n1207 585
R2883 VSS.n1198 VSS.n1197 585
R2884 VSS.n1287 VSS.n1198 585
R2885 VSS.n1158 VSS.n1157 585
R2886 VSS.n1157 VSS.n1156 585
R2887 VSS.n1295 VSS.n1292 585
R2888 VSS.n17942 VSS.n1292 585
R2889 VSS.n1322 VSS.n1321 585
R2890 VSS.n17926 VSS.n1322 585
R2891 VSS.n17913 VSS.n17912 585
R2892 VSS.n17912 VSS.n17911 585
R2893 VSS.n1405 VSS.n1404 585
R2894 VSS.n1406 VSS.n1405 585
R2895 VSS.n1413 VSS.n1412 585
R2896 VSS.t629 VSS.n1413 585
R2897 VSS.n1394 VSS.n1392 585
R2898 VSS.n17875 VSS.n1394 585
R2899 VSS.n17873 VSS.n17872 585
R2900 VSS.n17874 VSS.n17873 585
R2901 VSS.n1411 VSS.n1393 585
R2902 VSS.n1414 VSS.n1393 585
R2903 VSS.n1408 VSS.n1375 585
R2904 VSS.n1408 VSS.n1407 585
R2905 VSS.n17929 VSS.n17928 585
R2906 VSS.n17928 VSS.n17927 585
R2907 VSS.n17914 VSS.n1324 585
R2908 VSS.n1324 VSS.n1323 585
R2909 VSS.n1422 VSS.n1421 585
R2910 VSS.n1289 VSS.n1288 585
R2911 VSS.n17940 VSS.n17939 585
R2912 VSS.n17941 VSS.n17940 585
R2913 VSS.n17943 VSS.n17942 403.461
R2914 VSS.n17925 VSS.n1323 403.461
R2915 VSS.n1407 VSS.n1395 403.461
R2916 VSS.n17876 VSS.n1414 403.461
R2917 VSS.n17874 VSS.n1415 403.461
R2918 VSS.n1247 VSS.n1246 396.599
R2919 VSS.n1254 VSS.n1253 396.599
R2920 VSS.n1255 VSS.n1254 396.599
R2921 VSS.n1271 VSS.n1270 396.599
R2922 VSS.n1286 VSS.n1199 396.599
R2923 VSS.n17910 VSS.n17909 395.849
R2924 VSS.n17909 VSS.n1341 395.849
R2925 VSS.n17120 VSS.n17119 338.954
R2926 VSS.n17167 VSS.n17165 338.954
R2927 VSS.n17236 VSS.n16881 338.954
R2928 VSS.n17237 VSS.n16868 338.954
R2929 VSS.n17264 VSS.n17262 338.954
R2930 VSS.n17712 VSS.n17711 338.954
R2931 VSS.n17759 VSS.n17757 338.954
R2932 VSS.n17828 VSS.n17295 338.954
R2933 VSS.n17829 VSS.n17282 338.954
R2934 VSS.n17856 VSS.n17854 338.954
R2935 VSS.n9762 VSS.n9761 338.954
R2936 VSS.n9809 VSS.n9807 338.954
R2937 VSS.n9878 VSS.n9345 338.954
R2938 VSS.n9879 VSS.n9333 338.954
R2939 VSS.n9907 VSS.n9905 338.954
R2940 VSS.n16705 VSS.n16704 338.954
R2941 VSS.n16752 VSS.n16750 338.954
R2942 VSS.n16821 VSS.n16287 338.954
R2943 VSS.n16822 VSS.n16275 338.954
R2944 VSS.n16850 VSS.n16848 338.954
R2945 VSS.n16112 VSS.n16111 338.954
R2946 VSS.n16159 VSS.n16157 338.954
R2947 VSS.n16228 VSS.n1459 338.954
R2948 VSS.n16229 VSS.n1447 338.954
R2949 VSS.n16257 VSS.n16255 338.954
R2950 VSS.n2297 VSS.n2296 338.954
R2951 VSS.n2279 VSS.n2105 338.954
R2952 VSS.n2189 VSS.n2177 338.954
R2953 VSS.n2230 VSS.n2196 338.954
R2954 VSS.n2228 VSS.n2197 338.954
R2955 VSS.n3253 VSS.n3252 338.954
R2956 VSS.n3300 VSS.n3298 338.954
R2957 VSS.n3369 VSS.n2836 338.954
R2958 VSS.n3370 VSS.n2824 338.954
R2959 VSS.n3398 VSS.n3396 338.954
R2960 VSS.n3845 VSS.n3844 338.954
R2961 VSS.n3892 VSS.n3890 338.954
R2962 VSS.n3961 VSS.n3428 338.954
R2963 VSS.n3962 VSS.n3416 338.954
R2964 VSS.n3990 VSS.n3988 338.954
R2965 VSS.n4437 VSS.n4436 338.954
R2966 VSS.n4484 VSS.n4482 338.954
R2967 VSS.n4553 VSS.n4020 338.954
R2968 VSS.n4554 VSS.n4008 338.954
R2969 VSS.n4582 VSS.n4580 338.954
R2970 VSS.n5029 VSS.n5028 338.954
R2971 VSS.n5076 VSS.n5074 338.954
R2972 VSS.n5145 VSS.n4612 338.954
R2973 VSS.n5146 VSS.n4600 338.954
R2974 VSS.n5174 VSS.n5172 338.954
R2975 VSS.n5262 VSS.n5261 338.954
R2976 VSS.n5244 VSS.n2701 338.954
R2977 VSS.n2785 VSS.n2773 338.954
R2978 VSS.n5195 VSS.n2792 338.954
R2979 VSS.n5193 VSS.n2793 338.954
R2980 VSS.n5835 VSS.n5834 338.954
R2981 VSS.n5817 VSS.n5662 338.954
R2982 VSS.n5759 VSS.n5747 338.954
R2983 VSS.n5768 VSS.n5766 338.954
R2984 VSS.n18880 VSS.n9 338.954
R2985 VSS.n6427 VSS.n6426 338.954
R2986 VSS.n6409 VSS.n6235 338.954
R2987 VSS.n6319 VSS.n6307 338.954
R2988 VSS.n6360 VSS.n6326 338.954
R2989 VSS.n6358 VSS.n6327 338.954
R2990 VSS.n7986 VSS.n7985 338.954
R2991 VSS.n8033 VSS.n8031 338.954
R2992 VSS.n8102 VSS.n7569 338.954
R2993 VSS.n8103 VSS.n7557 338.954
R2994 VSS.n8131 VSS.n8129 338.954
R2995 VSS.n8578 VSS.n8577 338.954
R2996 VSS.n8625 VSS.n8623 338.954
R2997 VSS.n8694 VSS.n8161 338.954
R2998 VSS.n8695 VSS.n8149 338.954
R2999 VSS.n8723 VSS.n8721 338.954
R3000 VSS.n9170 VSS.n9169 338.954
R3001 VSS.n9217 VSS.n9215 338.954
R3002 VSS.n9286 VSS.n8753 338.954
R3003 VSS.n9287 VSS.n8741 338.954
R3004 VSS.n9315 VSS.n9313 338.954
R3005 VSS.n10354 VSS.n10353 338.954
R3006 VSS.n10401 VSS.n10399 338.954
R3007 VSS.n10470 VSS.n9937 338.954
R3008 VSS.n10471 VSS.n9925 338.954
R3009 VSS.n10499 VSS.n10497 338.954
R3010 VSS.n10946 VSS.n10945 338.954
R3011 VSS.n10993 VSS.n10991 338.954
R3012 VSS.n11062 VSS.n10529 338.954
R3013 VSS.n11063 VSS.n10517 338.954
R3014 VSS.n11091 VSS.n11089 338.954
R3015 VSS.n11538 VSS.n11537 338.954
R3016 VSS.n11585 VSS.n11583 338.954
R3017 VSS.n11654 VSS.n11121 338.954
R3018 VSS.n11655 VSS.n11109 338.954
R3019 VSS.n11683 VSS.n11681 338.954
R3020 VSS.n12130 VSS.n12129 338.954
R3021 VSS.n12177 VSS.n12175 338.954
R3022 VSS.n12246 VSS.n11713 338.954
R3023 VSS.n12247 VSS.n11701 338.954
R3024 VSS.n12275 VSS.n12273 338.954
R3025 VSS.n12722 VSS.n12721 338.954
R3026 VSS.n12769 VSS.n12767 338.954
R3027 VSS.n12838 VSS.n12305 338.954
R3028 VSS.n12839 VSS.n12293 338.954
R3029 VSS.n12867 VSS.n12865 338.954
R3030 VSS.n13314 VSS.n13313 338.954
R3031 VSS.n13361 VSS.n13359 338.954
R3032 VSS.n13430 VSS.n12897 338.954
R3033 VSS.n13431 VSS.n12885 338.954
R3034 VSS.n13459 VSS.n13457 338.954
R3035 VSS.n13906 VSS.n13905 338.954
R3036 VSS.n13953 VSS.n13951 338.954
R3037 VSS.n14022 VSS.n13489 338.954
R3038 VSS.n14023 VSS.n13477 338.954
R3039 VSS.n14051 VSS.n14049 338.954
R3040 VSS.n14498 VSS.n14497 338.954
R3041 VSS.n14545 VSS.n14543 338.954
R3042 VSS.n14614 VSS.n14081 338.954
R3043 VSS.n14615 VSS.n14069 338.954
R3044 VSS.n14643 VSS.n14641 338.954
R3045 VSS.n15090 VSS.n15089 338.954
R3046 VSS.n15137 VSS.n15135 338.954
R3047 VSS.n15206 VSS.n14673 338.954
R3048 VSS.n15207 VSS.n14661 338.954
R3049 VSS.n15235 VSS.n15233 338.954
R3050 VSS.n15682 VSS.n15681 338.954
R3051 VSS.n15729 VSS.n15727 338.954
R3052 VSS.n15798 VSS.n15265 338.954
R3053 VSS.n15799 VSS.n15253 338.954
R3054 VSS.n15827 VSS.n15825 338.954
R3055 VSS.n15915 VSS.n15914 338.954
R3056 VSS.n15897 VSS.n6841 338.954
R3057 VSS.n6925 VSS.n6913 338.954
R3058 VSS.n15848 VSS.n6932 338.954
R3059 VSS.n15846 VSS.n6933 338.954
R3060 VSS.n7394 VSS.n7393 338.954
R3061 VSS.n7441 VSS.n7439 338.954
R3062 VSS.n7510 VSS.n6976 338.954
R3063 VSS.n7511 VSS.n6964 338.954
R3064 VSS.n7539 VSS.n7537 338.954
R3065 VSS.n18706 VSS.n18705 338.954
R3066 VSS.n18753 VSS.n18751 338.954
R3067 VSS.n18822 VSS.n74 338.954
R3068 VSS.n18823 VSS.n62 338.954
R3069 VSS.n18851 VSS.n18849 338.954
R3070 VSS.n18532 VSS.n18531 338.954
R3071 VSS.n18371 VSS.n18361 338.954
R3072 VSS.n18450 VSS.n18384 338.954
R3073 VSS.n18451 VSS.n18439 338.954
R3074 VSS.n18460 VSS.n18458 338.954
R3075 VSS.n829 VSS.n828 338.954
R3076 VSS.n811 VSS.n664 338.954
R3077 VSS.n759 VSS.n745 338.954
R3078 VSS.n760 VSS.n46 338.954
R3079 VSS.n18872 VSS.n18871 338.954
R3080 VSS.n17215 VSS.n16893 332.558
R3081 VSS.n17216 VSS.n17215 332.558
R3082 VSS.n17807 VSS.n17307 332.558
R3083 VSS.n17808 VSS.n17807 332.558
R3084 VSS.n9857 VSS.n9357 332.558
R3085 VSS.n9858 VSS.n9857 332.558
R3086 VSS.n16800 VSS.n16299 332.558
R3087 VSS.n16801 VSS.n16800 332.558
R3088 VSS.n16207 VSS.n1471 332.558
R3089 VSS.n16208 VSS.n16207 332.558
R3090 VSS.n2264 VSS.n2263 332.558
R3091 VSS.n2263 VSS.n2123 332.558
R3092 VSS.n3348 VSS.n2848 332.558
R3093 VSS.n3349 VSS.n3348 332.558
R3094 VSS.n3940 VSS.n3440 332.558
R3095 VSS.n3941 VSS.n3940 332.558
R3096 VSS.n4532 VSS.n4032 332.558
R3097 VSS.n4533 VSS.n4532 332.558
R3098 VSS.n5124 VSS.n4624 332.558
R3099 VSS.n5125 VSS.n5124 332.558
R3100 VSS.n5229 VSS.n5228 332.558
R3101 VSS.n5228 VSS.n2719 332.558
R3102 VSS.n5802 VSS.n5801 332.558
R3103 VSS.n5801 VSS.n5680 332.558
R3104 VSS.n6394 VSS.n6393 332.558
R3105 VSS.n6393 VSS.n6253 332.558
R3106 VSS.n8081 VSS.n7581 332.558
R3107 VSS.n8082 VSS.n8081 332.558
R3108 VSS.n8673 VSS.n8173 332.558
R3109 VSS.n8674 VSS.n8673 332.558
R3110 VSS.n9265 VSS.n8765 332.558
R3111 VSS.n9266 VSS.n9265 332.558
R3112 VSS.n10449 VSS.n9949 332.558
R3113 VSS.n10450 VSS.n10449 332.558
R3114 VSS.n11041 VSS.n10541 332.558
R3115 VSS.n11042 VSS.n11041 332.558
R3116 VSS.n11633 VSS.n11133 332.558
R3117 VSS.n11634 VSS.n11633 332.558
R3118 VSS.n12225 VSS.n11725 332.558
R3119 VSS.n12226 VSS.n12225 332.558
R3120 VSS.n12817 VSS.n12317 332.558
R3121 VSS.n12818 VSS.n12817 332.558
R3122 VSS.n13409 VSS.n12909 332.558
R3123 VSS.n13410 VSS.n13409 332.558
R3124 VSS.n14001 VSS.n13501 332.558
R3125 VSS.n14002 VSS.n14001 332.558
R3126 VSS.n14593 VSS.n14093 332.558
R3127 VSS.n14594 VSS.n14593 332.558
R3128 VSS.n15185 VSS.n14685 332.558
R3129 VSS.n15186 VSS.n15185 332.558
R3130 VSS.n15777 VSS.n15277 332.558
R3131 VSS.n15778 VSS.n15777 332.558
R3132 VSS.n15882 VSS.n15881 332.558
R3133 VSS.n15881 VSS.n6859 332.558
R3134 VSS.n7489 VSS.n6988 332.558
R3135 VSS.n7490 VSS.n7489 332.558
R3136 VSS.n18801 VSS.n86 332.558
R3137 VSS.n18802 VSS.n18801 332.558
R3138 VSS.n18496 VSS.n18383 332.558
R3139 VSS.n18496 VSS.n18495 332.558
R3140 VSS.n796 VSS.n795 332.558
R3141 VSS.n795 VSS.n682 332.558
R3142 VSS.n10171 VSS.n10167 329.844
R3143 VSS.n10169 VSS.n10100 329.844
R3144 VSS.n10200 VSS.n10100 329.844
R3145 VSS.n10204 VSS.n10203 329.844
R3146 VSS.n10233 VSS.n10232 329.844
R3147 VSS.n17030 VSS.n16974 329.38
R3148 VSS.n17053 VSS.n17051 329.38
R3149 VSS.n17053 VSS.n17052 329.38
R3150 VSS.n17082 VSS.n17081 329.38
R3151 VSS.n17103 VSS.n16938 329.38
R3152 VSS.n17622 VSS.n17388 329.38
R3153 VSS.n17645 VSS.n17643 329.38
R3154 VSS.n17645 VSS.n17644 329.38
R3155 VSS.n17674 VSS.n17673 329.38
R3156 VSS.n17695 VSS.n17352 329.38
R3157 VSS.n18106 VSS.n18102 329.38
R3158 VSS.n18104 VSS.n250 329.38
R3159 VSS.n18135 VSS.n250 329.38
R3160 VSS.n18139 VSS.n18138 329.38
R3161 VSS.n18168 VSS.n18167 329.38
R3162 VSS.n9672 VSS.n9438 329.38
R3163 VSS.n9695 VSS.n9693 329.38
R3164 VSS.n9695 VSS.n9694 329.38
R3165 VSS.n9724 VSS.n9723 329.38
R3166 VSS.n9745 VSS.n9402 329.38
R3167 VSS.n16615 VSS.n16380 329.38
R3168 VSS.n16638 VSS.n16636 329.38
R3169 VSS.n16638 VSS.n16637 329.38
R3170 VSS.n16667 VSS.n16666 329.38
R3171 VSS.n16688 VSS.n16344 329.38
R3172 VSS.n16510 VSS.n16457 329.38
R3173 VSS.n16533 VSS.n16531 329.38
R3174 VSS.n16533 VSS.n16532 329.38
R3175 VSS.n16562 VSS.n16561 329.38
R3176 VSS.n16584 VSS.n16419 329.38
R3177 VSS.n16022 VSS.n1552 329.38
R3178 VSS.n16045 VSS.n16043 329.38
R3179 VSS.n16045 VSS.n16044 329.38
R3180 VSS.n16074 VSS.n16073 329.38
R3181 VSS.n16095 VSS.n1516 329.38
R3182 VSS.n1675 VSS.n1622 329.38
R3183 VSS.n1698 VSS.n1696 329.38
R3184 VSS.n1698 VSS.n1697 329.38
R3185 VSS.n1727 VSS.n1726 329.38
R3186 VSS.n1749 VSS.n1584 329.38
R3187 VSS.n2029 VSS.n2028 329.38
R3188 VSS.n2036 VSS.n2035 329.38
R3189 VSS.n2037 VSS.n2036 329.38
R3190 VSS.n2053 VSS.n2052 329.38
R3191 VSS.n2068 VSS.n1981 329.38
R3192 VSS.n1871 VSS.n1867 329.38
R3193 VSS.n1869 VSS.n1800 329.38
R3194 VSS.n1900 VSS.n1800 329.38
R3195 VSS.n1904 VSS.n1903 329.38
R3196 VSS.n1933 VSS.n1932 329.38
R3197 VSS.n3163 VSS.n2929 329.38
R3198 VSS.n3186 VSS.n3184 329.38
R3199 VSS.n3186 VSS.n3185 329.38
R3200 VSS.n3215 VSS.n3214 329.38
R3201 VSS.n3236 VSS.n2893 329.38
R3202 VSS.n3070 VSS.n3066 329.38
R3203 VSS.n3068 VSS.n2999 329.38
R3204 VSS.n3099 VSS.n2999 329.38
R3205 VSS.n3103 VSS.n3102 329.38
R3206 VSS.n3132 VSS.n3131 329.38
R3207 VSS.n3755 VSS.n3521 329.38
R3208 VSS.n3778 VSS.n3776 329.38
R3209 VSS.n3778 VSS.n3777 329.38
R3210 VSS.n3807 VSS.n3806 329.38
R3211 VSS.n3828 VSS.n3485 329.38
R3212 VSS.n3662 VSS.n3658 329.38
R3213 VSS.n3660 VSS.n3591 329.38
R3214 VSS.n3691 VSS.n3591 329.38
R3215 VSS.n3695 VSS.n3694 329.38
R3216 VSS.n3724 VSS.n3723 329.38
R3217 VSS.n4347 VSS.n4113 329.38
R3218 VSS.n4370 VSS.n4368 329.38
R3219 VSS.n4370 VSS.n4369 329.38
R3220 VSS.n4399 VSS.n4398 329.38
R3221 VSS.n4420 VSS.n4077 329.38
R3222 VSS.n4254 VSS.n4250 329.38
R3223 VSS.n4252 VSS.n4183 329.38
R3224 VSS.n4283 VSS.n4183 329.38
R3225 VSS.n4287 VSS.n4286 329.38
R3226 VSS.n4316 VSS.n4315 329.38
R3227 VSS.n4939 VSS.n4705 329.38
R3228 VSS.n4962 VSS.n4960 329.38
R3229 VSS.n4962 VSS.n4961 329.38
R3230 VSS.n4991 VSS.n4990 329.38
R3231 VSS.n5012 VSS.n4669 329.38
R3232 VSS.n4846 VSS.n4842 329.38
R3233 VSS.n4844 VSS.n4775 329.38
R3234 VSS.n4875 VSS.n4775 329.38
R3235 VSS.n4879 VSS.n4878 329.38
R3236 VSS.n4908 VSS.n4907 329.38
R3237 VSS.n2625 VSS.n2624 329.38
R3238 VSS.n2632 VSS.n2631 329.38
R3239 VSS.n2633 VSS.n2632 329.38
R3240 VSS.n2649 VSS.n2648 329.38
R3241 VSS.n2664 VSS.n2577 329.38
R3242 VSS.n2467 VSS.n2463 329.38
R3243 VSS.n2465 VSS.n2396 329.38
R3244 VSS.n2496 VSS.n2396 329.38
R3245 VSS.n2500 VSS.n2499 329.38
R3246 VSS.n2529 VSS.n2528 329.38
R3247 VSS.n5586 VSS.n5585 329.38
R3248 VSS.n5593 VSS.n5592 329.38
R3249 VSS.n5594 VSS.n5593 329.38
R3250 VSS.n5610 VSS.n5609 329.38
R3251 VSS.n5625 VSS.n5538 329.38
R3252 VSS.n5428 VSS.n5424 329.38
R3253 VSS.n5426 VSS.n5357 329.38
R3254 VSS.n5457 VSS.n5357 329.38
R3255 VSS.n5461 VSS.n5460 329.38
R3256 VSS.n5490 VSS.n5489 329.38
R3257 VSS.n6159 VSS.n6158 329.38
R3258 VSS.n6166 VSS.n6165 329.38
R3259 VSS.n6167 VSS.n6166 329.38
R3260 VSS.n6183 VSS.n6182 329.38
R3261 VSS.n6198 VSS.n6111 329.38
R3262 VSS.n6001 VSS.n5997 329.38
R3263 VSS.n5999 VSS.n5930 329.38
R3264 VSS.n6030 VSS.n5930 329.38
R3265 VSS.n6034 VSS.n6033 329.38
R3266 VSS.n6063 VSS.n6062 329.38
R3267 VSS.n7896 VSS.n7662 329.38
R3268 VSS.n7919 VSS.n7917 329.38
R3269 VSS.n7919 VSS.n7918 329.38
R3270 VSS.n7948 VSS.n7947 329.38
R3271 VSS.n7969 VSS.n7626 329.38
R3272 VSS.n7803 VSS.n7799 329.38
R3273 VSS.n7801 VSS.n7732 329.38
R3274 VSS.n7832 VSS.n7732 329.38
R3275 VSS.n7836 VSS.n7835 329.38
R3276 VSS.n7865 VSS.n7864 329.38
R3277 VSS.n8488 VSS.n8254 329.38
R3278 VSS.n8511 VSS.n8509 329.38
R3279 VSS.n8511 VSS.n8510 329.38
R3280 VSS.n8540 VSS.n8539 329.38
R3281 VSS.n8561 VSS.n8218 329.38
R3282 VSS.n8395 VSS.n8391 329.38
R3283 VSS.n8393 VSS.n8324 329.38
R3284 VSS.n8424 VSS.n8324 329.38
R3285 VSS.n8428 VSS.n8427 329.38
R3286 VSS.n8457 VSS.n8456 329.38
R3287 VSS.n9080 VSS.n8846 329.38
R3288 VSS.n9103 VSS.n9101 329.38
R3289 VSS.n9103 VSS.n9102 329.38
R3290 VSS.n9132 VSS.n9131 329.38
R3291 VSS.n9153 VSS.n8810 329.38
R3292 VSS.n8987 VSS.n8983 329.38
R3293 VSS.n8985 VSS.n8916 329.38
R3294 VSS.n9016 VSS.n8916 329.38
R3295 VSS.n9020 VSS.n9019 329.38
R3296 VSS.n9049 VSS.n9048 329.38
R3297 VSS.n10264 VSS.n10030 329.38
R3298 VSS.n10287 VSS.n10285 329.38
R3299 VSS.n10287 VSS.n10286 329.38
R3300 VSS.n10316 VSS.n10315 329.38
R3301 VSS.n10337 VSS.n9994 329.38
R3302 VSS.n10856 VSS.n10622 329.38
R3303 VSS.n10879 VSS.n10877 329.38
R3304 VSS.n10879 VSS.n10878 329.38
R3305 VSS.n10908 VSS.n10907 329.38
R3306 VSS.n10929 VSS.n10586 329.38
R3307 VSS.n10763 VSS.n10759 329.38
R3308 VSS.n10761 VSS.n10692 329.38
R3309 VSS.n10792 VSS.n10692 329.38
R3310 VSS.n10796 VSS.n10795 329.38
R3311 VSS.n10825 VSS.n10824 329.38
R3312 VSS.n11448 VSS.n11214 329.38
R3313 VSS.n11471 VSS.n11469 329.38
R3314 VSS.n11471 VSS.n11470 329.38
R3315 VSS.n11500 VSS.n11499 329.38
R3316 VSS.n11521 VSS.n11178 329.38
R3317 VSS.n11355 VSS.n11351 329.38
R3318 VSS.n11353 VSS.n11284 329.38
R3319 VSS.n11384 VSS.n11284 329.38
R3320 VSS.n11388 VSS.n11387 329.38
R3321 VSS.n11417 VSS.n11416 329.38
R3322 VSS.n12040 VSS.n11806 329.38
R3323 VSS.n12063 VSS.n12061 329.38
R3324 VSS.n12063 VSS.n12062 329.38
R3325 VSS.n12092 VSS.n12091 329.38
R3326 VSS.n12113 VSS.n11770 329.38
R3327 VSS.n11947 VSS.n11943 329.38
R3328 VSS.n11945 VSS.n11876 329.38
R3329 VSS.n11976 VSS.n11876 329.38
R3330 VSS.n11980 VSS.n11979 329.38
R3331 VSS.n12009 VSS.n12008 329.38
R3332 VSS.n12632 VSS.n12398 329.38
R3333 VSS.n12655 VSS.n12653 329.38
R3334 VSS.n12655 VSS.n12654 329.38
R3335 VSS.n12684 VSS.n12683 329.38
R3336 VSS.n12705 VSS.n12362 329.38
R3337 VSS.n12539 VSS.n12535 329.38
R3338 VSS.n12537 VSS.n12468 329.38
R3339 VSS.n12568 VSS.n12468 329.38
R3340 VSS.n12572 VSS.n12571 329.38
R3341 VSS.n12601 VSS.n12600 329.38
R3342 VSS.n13224 VSS.n12990 329.38
R3343 VSS.n13247 VSS.n13245 329.38
R3344 VSS.n13247 VSS.n13246 329.38
R3345 VSS.n13276 VSS.n13275 329.38
R3346 VSS.n13297 VSS.n12954 329.38
R3347 VSS.n13131 VSS.n13127 329.38
R3348 VSS.n13129 VSS.n13060 329.38
R3349 VSS.n13160 VSS.n13060 329.38
R3350 VSS.n13164 VSS.n13163 329.38
R3351 VSS.n13193 VSS.n13192 329.38
R3352 VSS.n13816 VSS.n13582 329.38
R3353 VSS.n13839 VSS.n13837 329.38
R3354 VSS.n13839 VSS.n13838 329.38
R3355 VSS.n13868 VSS.n13867 329.38
R3356 VSS.n13889 VSS.n13546 329.38
R3357 VSS.n13723 VSS.n13719 329.38
R3358 VSS.n13721 VSS.n13652 329.38
R3359 VSS.n13752 VSS.n13652 329.38
R3360 VSS.n13756 VSS.n13755 329.38
R3361 VSS.n13785 VSS.n13784 329.38
R3362 VSS.n14408 VSS.n14174 329.38
R3363 VSS.n14431 VSS.n14429 329.38
R3364 VSS.n14431 VSS.n14430 329.38
R3365 VSS.n14460 VSS.n14459 329.38
R3366 VSS.n14481 VSS.n14138 329.38
R3367 VSS.n14315 VSS.n14311 329.38
R3368 VSS.n14313 VSS.n14244 329.38
R3369 VSS.n14344 VSS.n14244 329.38
R3370 VSS.n14348 VSS.n14347 329.38
R3371 VSS.n14377 VSS.n14376 329.38
R3372 VSS.n15000 VSS.n14766 329.38
R3373 VSS.n15023 VSS.n15021 329.38
R3374 VSS.n15023 VSS.n15022 329.38
R3375 VSS.n15052 VSS.n15051 329.38
R3376 VSS.n15073 VSS.n14730 329.38
R3377 VSS.n14907 VSS.n14903 329.38
R3378 VSS.n14905 VSS.n14836 329.38
R3379 VSS.n14936 VSS.n14836 329.38
R3380 VSS.n14940 VSS.n14939 329.38
R3381 VSS.n14969 VSS.n14968 329.38
R3382 VSS.n15592 VSS.n15358 329.38
R3383 VSS.n15615 VSS.n15613 329.38
R3384 VSS.n15615 VSS.n15614 329.38
R3385 VSS.n15644 VSS.n15643 329.38
R3386 VSS.n15665 VSS.n15322 329.38
R3387 VSS.n15499 VSS.n15495 329.38
R3388 VSS.n15497 VSS.n15428 329.38
R3389 VSS.n15528 VSS.n15428 329.38
R3390 VSS.n15532 VSS.n15531 329.38
R3391 VSS.n15561 VSS.n15560 329.38
R3392 VSS.n6765 VSS.n6764 329.38
R3393 VSS.n6772 VSS.n6771 329.38
R3394 VSS.n6773 VSS.n6772 329.38
R3395 VSS.n6789 VSS.n6788 329.38
R3396 VSS.n6804 VSS.n6717 329.38
R3397 VSS.n6607 VSS.n6603 329.38
R3398 VSS.n6605 VSS.n6536 329.38
R3399 VSS.n6636 VSS.n6536 329.38
R3400 VSS.n6640 VSS.n6639 329.38
R3401 VSS.n6669 VSS.n6668 329.38
R3402 VSS.n7304 VSS.n7069 329.38
R3403 VSS.n7327 VSS.n7325 329.38
R3404 VSS.n7327 VSS.n7326 329.38
R3405 VSS.n7356 VSS.n7355 329.38
R3406 VSS.n7377 VSS.n7033 329.38
R3407 VSS.n7199 VSS.n7146 329.38
R3408 VSS.n7222 VSS.n7220 329.38
R3409 VSS.n7222 VSS.n7221 329.38
R3410 VSS.n7251 VSS.n7250 329.38
R3411 VSS.n7273 VSS.n7108 329.38
R3412 VSS.n18616 VSS.n167 329.38
R3413 VSS.n18639 VSS.n18637 329.38
R3414 VSS.n18639 VSS.n18638 329.38
R3415 VSS.n18668 VSS.n18667 329.38
R3416 VSS.n18689 VSS.n131 329.38
R3417 VSS.n373 VSS.n340 329.38
R3418 VSS.n375 VSS.n336 329.38
R3419 VSS.n382 VSS.n336 329.38
R3420 VSS.n384 VSS.n330 329.38
R3421 VSS.n401 VSS.n400 329.38
R3422 VSS.n18264 VSS.n18263 329.38
R3423 VSS.n18271 VSS.n18270 329.38
R3424 VSS.n18272 VSS.n18271 329.38
R3425 VSS.n18288 VSS.n18287 329.38
R3426 VSS.n18303 VSS.n18216 329.38
R3427 VSS.n588 VSS.n587 329.38
R3428 VSS.n595 VSS.n594 329.38
R3429 VSS.n596 VSS.n595 329.38
R3430 VSS.n612 VSS.n611 329.38
R3431 VSS.n627 VSS.n537 329.38
R3432 VSS.n931 VSS.n930 329.38
R3433 VSS.n938 VSS.n937 329.38
R3434 VSS.n939 VSS.n938 329.38
R3435 VSS.n955 VSS.n954 329.38
R3436 VSS.n971 VSS.n884 329.38
R3437 VSS.n1112 VSS.n1111 329.38
R3438 VSS.n1119 VSS.n1118 329.38
R3439 VSS.n1120 VSS.n1119 329.38
R3440 VSS.n1136 VSS.n1135 329.38
R3441 VSS.n1152 VSS.n1065 329.38
R3442 VSS.n9579 VSS.n9575 328.914
R3443 VSS.n9577 VSS.n9508 328.914
R3444 VSS.n9608 VSS.n9508 328.914
R3445 VSS.n9612 VSS.n9611 328.914
R3446 VSS.n9641 VSS.n9640 328.914
R3447 VSS.t198 VSS.n1293 304.498
R3448 VSS.n17214 VSS.n17213 292.5
R3449 VSS.n17215 VSS.n17214 292.5
R3450 VSS.n17806 VSS.n17805 292.5
R3451 VSS.n17807 VSS.n17806 292.5
R3452 VSS.n9856 VSS.n9855 292.5
R3453 VSS.n9857 VSS.n9856 292.5
R3454 VSS.n16799 VSS.n16798 292.5
R3455 VSS.n16800 VSS.n16799 292.5
R3456 VSS.n16206 VSS.n16205 292.5
R3457 VSS.n16207 VSS.n16206 292.5
R3458 VSS.n2262 VSS.n2261 292.5
R3459 VSS.n2263 VSS.n2262 292.5
R3460 VSS.n3347 VSS.n3346 292.5
R3461 VSS.n3348 VSS.n3347 292.5
R3462 VSS.n3939 VSS.n3938 292.5
R3463 VSS.n3940 VSS.n3939 292.5
R3464 VSS.n4531 VSS.n4530 292.5
R3465 VSS.n4532 VSS.n4531 292.5
R3466 VSS.n5123 VSS.n5122 292.5
R3467 VSS.n5124 VSS.n5123 292.5
R3468 VSS.n5227 VSS.n5226 292.5
R3469 VSS.n5228 VSS.n5227 292.5
R3470 VSS.n5800 VSS.n5799 292.5
R3471 VSS.n5801 VSS.n5800 292.5
R3472 VSS.n6392 VSS.n6391 292.5
R3473 VSS.n6393 VSS.n6392 292.5
R3474 VSS.n8080 VSS.n8079 292.5
R3475 VSS.n8081 VSS.n8080 292.5
R3476 VSS.n8672 VSS.n8671 292.5
R3477 VSS.n8673 VSS.n8672 292.5
R3478 VSS.n9264 VSS.n9263 292.5
R3479 VSS.n9265 VSS.n9264 292.5
R3480 VSS.n10448 VSS.n10447 292.5
R3481 VSS.n10449 VSS.n10448 292.5
R3482 VSS.n11040 VSS.n11039 292.5
R3483 VSS.n11041 VSS.n11040 292.5
R3484 VSS.n11632 VSS.n11631 292.5
R3485 VSS.n11633 VSS.n11632 292.5
R3486 VSS.n12224 VSS.n12223 292.5
R3487 VSS.n12225 VSS.n12224 292.5
R3488 VSS.n12816 VSS.n12815 292.5
R3489 VSS.n12817 VSS.n12816 292.5
R3490 VSS.n13408 VSS.n13407 292.5
R3491 VSS.n13409 VSS.n13408 292.5
R3492 VSS.n14000 VSS.n13999 292.5
R3493 VSS.n14001 VSS.n14000 292.5
R3494 VSS.n14592 VSS.n14591 292.5
R3495 VSS.n14593 VSS.n14592 292.5
R3496 VSS.n15184 VSS.n15183 292.5
R3497 VSS.n15185 VSS.n15184 292.5
R3498 VSS.n15776 VSS.n15775 292.5
R3499 VSS.n15777 VSS.n15776 292.5
R3500 VSS.n15880 VSS.n15879 292.5
R3501 VSS.n15881 VSS.n15880 292.5
R3502 VSS.n7488 VSS.n7487 292.5
R3503 VSS.n7489 VSS.n7488 292.5
R3504 VSS.n18800 VSS.n18799 292.5
R3505 VSS.n18801 VSS.n18800 292.5
R3506 VSS.n18498 VSS.n18497 292.5
R3507 VSS.n18497 VSS.n18496 292.5
R3508 VSS.n794 VSS.n793 292.5
R3509 VSS.n795 VSS.n794 292.5
R3510 VSS.n17908 VSS.n17907 292.5
R3511 VSS.n17909 VSS.n17908 292.5
R3512 VSS.n17123 VSS.n17122 290.906
R3513 VSS.n17266 VSS.n16865 290.906
R3514 VSS.n17715 VSS.n17714 290.906
R3515 VSS.n17858 VSS.n17279 290.906
R3516 VSS.n18535 VSS.n18534 290.906
R3517 VSS.n18462 VSS.n18436 290.906
R3518 VSS.n9765 VSS.n9764 290.906
R3519 VSS.n9909 VSS.n9330 290.906
R3520 VSS.n16708 VSS.n16707 290.906
R3521 VSS.n16852 VSS.n16272 290.906
R3522 VSS.n16115 VSS.n16114 290.906
R3523 VSS.n16259 VSS.n1444 290.906
R3524 VSS.n2300 VSS.n2299 290.906
R3525 VSS.n2206 VSS.n2205 290.906
R3526 VSS.n3256 VSS.n3255 290.906
R3527 VSS.n3400 VSS.n2821 290.906
R3528 VSS.n3848 VSS.n3847 290.906
R3529 VSS.n3992 VSS.n3413 290.906
R3530 VSS.n4440 VSS.n4439 290.906
R3531 VSS.n4584 VSS.n4005 290.906
R3532 VSS.n5032 VSS.n5031 290.906
R3533 VSS.n5176 VSS.n4597 290.906
R3534 VSS.n5265 VSS.n5264 290.906
R3535 VSS.n2802 VSS.n2801 290.906
R3536 VSS.n5838 VSS.n5837 290.906
R3537 VSS.n18882 VSS.n6 290.906
R3538 VSS.n6430 VSS.n6429 290.906
R3539 VSS.n6336 VSS.n6335 290.906
R3540 VSS.n7989 VSS.n7988 290.906
R3541 VSS.n8133 VSS.n7554 290.906
R3542 VSS.n8581 VSS.n8580 290.906
R3543 VSS.n8725 VSS.n8146 290.906
R3544 VSS.n9173 VSS.n9172 290.906
R3545 VSS.n9317 VSS.n8738 290.906
R3546 VSS.n10357 VSS.n10356 290.906
R3547 VSS.n10501 VSS.n9922 290.906
R3548 VSS.n10949 VSS.n10948 290.906
R3549 VSS.n11093 VSS.n10514 290.906
R3550 VSS.n11541 VSS.n11540 290.906
R3551 VSS.n11685 VSS.n11106 290.906
R3552 VSS.n12133 VSS.n12132 290.906
R3553 VSS.n12277 VSS.n11698 290.906
R3554 VSS.n12725 VSS.n12724 290.906
R3555 VSS.n12869 VSS.n12290 290.906
R3556 VSS.n13317 VSS.n13316 290.906
R3557 VSS.n13461 VSS.n12882 290.906
R3558 VSS.n13909 VSS.n13908 290.906
R3559 VSS.n14053 VSS.n13474 290.906
R3560 VSS.n14501 VSS.n14500 290.906
R3561 VSS.n14645 VSS.n14066 290.906
R3562 VSS.n15093 VSS.n15092 290.906
R3563 VSS.n15237 VSS.n14658 290.906
R3564 VSS.n15685 VSS.n15684 290.906
R3565 VSS.n15829 VSS.n15250 290.906
R3566 VSS.n15918 VSS.n15917 290.906
R3567 VSS.n6942 VSS.n6941 290.906
R3568 VSS.n7397 VSS.n7396 290.906
R3569 VSS.n7541 VSS.n6961 290.906
R3570 VSS.n18709 VSS.n18708 290.906
R3571 VSS.n18853 VSS.n59 290.906
R3572 VSS.n832 VSS.n831 290.906
R3573 VSS.n18875 VSS.n18874 290.906
R3574 VSS.n17946 VSS.n17945 290.906
R3575 VSS.n1424 VSS.n1423 290.906
R3576 VSS.n17948 VSS.t196 269.807
R3577 VSS.n17112 VSS.t598 255.815
R3578 VSS.n17704 VSS.t120 255.815
R3579 VSS.n9754 VSS.t35 255.815
R3580 VSS.n16697 VSS.t490 255.815
R3581 VSS.n16104 VSS.t561 255.815
R3582 VSS.t78 VSS.n2075 255.815
R3583 VSS.n3245 VSS.t464 255.815
R3584 VSS.n3837 VSS.t611 255.815
R3585 VSS.n4429 VSS.t516 255.815
R3586 VSS.n5021 VSS.t176 255.815
R3587 VSS.t214 VSS.n2671 255.815
R3588 VSS.t116 VSS.n5632 255.815
R3589 VSS.t618 VSS.n6205 255.815
R3590 VSS.n7978 VSS.t239 255.815
R3591 VSS.n8570 VSS.t499 255.815
R3592 VSS.n9162 VSS.t541 255.815
R3593 VSS.n10346 VSS.t276 255.815
R3594 VSS.n10938 VSS.t587 255.815
R3595 VSS.n11530 VSS.t224 255.815
R3596 VSS.n12122 VSS.t306 255.815
R3597 VSS.n12714 VSS.t27 255.815
R3598 VSS.n13306 VSS.t328 255.815
R3599 VSS.n13898 VSS.t537 255.815
R3600 VSS.n14490 VSS.t316 255.815
R3601 VSS.n15082 VSS.t580 255.815
R3602 VSS.n15674 VSS.t594 255.815
R3603 VSS.t290 VSS.n6811 255.815
R3604 VSS.n7386 VSS.t431 255.815
R3605 VSS.n18698 VSS.t341 255.815
R3606 VSS.t286 VSS.n18310 255.815
R3607 VSS.t187 VSS.n634 255.815
R3608 VSS.t370 VSS.n1217 239.457
R3609 VSS.n17028 VSS.t523 198.87
R3610 VSS.n17620 VSS.t351 198.87
R3611 VSS.n9670 VSS.t477 198.87
R3612 VSS.n16613 VSS.t10 198.87
R3613 VSS.n16020 VSS.t344 198.87
R3614 VSS.t132 VSS.n1999 198.87
R3615 VSS.n3161 VSS.t591 198.87
R3616 VSS.n3753 VSS.t310 198.87
R3617 VSS.n4345 VSS.t212 198.87
R3618 VSS.n4937 VSS.t552 198.87
R3619 VSS.t91 VSS.n2595 198.87
R3620 VSS.t453 VSS.n5556 198.87
R3621 VSS.t219 VSS.n6129 198.87
R3622 VSS.n7894 VSS.t546 198.87
R3623 VSS.n8486 VSS.t483 198.87
R3624 VSS.n9078 VSS.t274 198.87
R3625 VSS.n10262 VSS.t124 198.87
R3626 VSS.n10854 VSS.t97 198.87
R3627 VSS.n11446 VSS.t203 198.87
R3628 VSS.n12038 VSS.t146 198.87
R3629 VSS.n12630 VSS.t252 198.87
R3630 VSS.n13222 VSS.t103 198.87
R3631 VSS.n13814 VSS.t446 198.87
R3632 VSS.n14406 VSS.t156 198.87
R3633 VSS.n14998 VSS.t159 198.87
R3634 VSS.n15590 VSS.t333 198.87
R3635 VSS.t480 VSS.n6735 198.87
R3636 VSS.n7302 VSS.t558 198.87
R3637 VSS.n18614 VSS.t391 198.87
R3638 VSS.t298 VSS.n18234 198.87
R3639 VSS.t573 VSS.n555 198.87
R3640 VSS.t106 VSS.n10123 192.929
R3641 VSS.t486 VSS.n273 192.655
R3642 VSS.n16508 VSS.t532 192.655
R3643 VSS.n1673 VSS.t53 192.655
R3644 VSS.t357 VSS.n1823 192.655
R3645 VSS.t209 VSS.n3022 192.655
R3646 VSS.t633 VSS.n3614 192.655
R3647 VSS.t565 VSS.n4206 192.655
R3648 VSS.t262 VSS.n4798 192.655
R3649 VSS.t509 VSS.n2419 192.655
R3650 VSS.t229 VSS.n5380 192.655
R3651 VSS.t24 VSS.n5953 192.655
R3652 VSS.t49 VSS.n7755 192.655
R3653 VSS.t326 VSS.n8347 192.655
R3654 VSS.t425 VSS.n8939 192.655
R3655 VSS.t608 VSS.n10715 192.655
R3656 VSS.t236 VSS.n11307 192.655
R3657 VSS.t338 VSS.n11899 192.655
R3658 VSS.t626 VSS.n12491 192.655
R3659 VSS.t355 VSS.n13083 192.655
R3660 VSS.t416 VSS.n13675 192.655
R3661 VSS.t555 VSS.n14267 192.655
R3662 VSS.t7 VSS.n14859 192.655
R3663 VSS.t605 VSS.n15451 192.655
R3664 VSS.t139 VSS.n6559 192.655
R3665 VSS.n7197 VSS.t21 192.655
R3666 VSS.n360 VSS.t389 192.655
R3667 VSS.t232 VSS.n903 192.655
R3668 VSS.t422 VSS.n1084 192.655
R3669 VSS.t88 VSS.n9531 192.385
R3670 VSS.n17125 VSS.t600 188.758
R3671 VSS.n17717 VSS.t122 188.758
R3672 VSS.n9767 VSS.t37 188.758
R3673 VSS.n16710 VSS.t492 188.758
R3674 VSS.n16117 VSS.t563 188.758
R3675 VSS.n2302 VSS.t80 188.758
R3676 VSS.n3258 VSS.t462 188.758
R3677 VSS.n3850 VSS.t613 188.758
R3678 VSS.n4442 VSS.t518 188.758
R3679 VSS.n5034 VSS.t178 188.758
R3680 VSS.n5267 VSS.t216 188.758
R3681 VSS.n5840 VSS.t118 188.758
R3682 VSS.n6432 VSS.t620 188.758
R3683 VSS.n7991 VSS.t241 188.758
R3684 VSS.n8583 VSS.t501 188.758
R3685 VSS.n9175 VSS.t543 188.758
R3686 VSS.n10359 VSS.t278 188.758
R3687 VSS.n10951 VSS.t589 188.758
R3688 VSS.n11543 VSS.t226 188.758
R3689 VSS.n12135 VSS.t308 188.758
R3690 VSS.n12727 VSS.t29 188.758
R3691 VSS.n13319 VSS.t330 188.758
R3692 VSS.n13911 VSS.t539 188.758
R3693 VSS.n14503 VSS.t318 188.758
R3694 VSS.n15095 VSS.t582 188.758
R3695 VSS.n15687 VSS.t596 188.758
R3696 VSS.n15920 VSS.t292 188.758
R3697 VSS.n7399 VSS.t433 188.758
R3698 VSS.n18711 VSS.t343 188.758
R3699 VSS.n18537 VSS.t288 188.758
R3700 VSS.n834 VSS.t189 188.758
R3701 VSS.n1219 VSS.t370 157.143
R3702 VSS.n10139 VSS.t106 136.917
R3703 VSS.n18074 VSS.t486 136.724
R3704 VSS.n16483 VSS.t532 136.724
R3705 VSS.n1648 VSS.t53 136.724
R3706 VSS.n1839 VSS.t357 136.724
R3707 VSS.n3038 VSS.t209 136.724
R3708 VSS.n3630 VSS.t633 136.724
R3709 VSS.n4222 VSS.t565 136.724
R3710 VSS.n4814 VSS.t262 136.724
R3711 VSS.n2435 VSS.t509 136.724
R3712 VSS.n5396 VSS.t229 136.724
R3713 VSS.n5969 VSS.t24 136.724
R3714 VSS.n7771 VSS.t49 136.724
R3715 VSS.n8363 VSS.t326 136.724
R3716 VSS.n8955 VSS.t425 136.724
R3717 VSS.n10731 VSS.t608 136.724
R3718 VSS.n11323 VSS.t236 136.724
R3719 VSS.n11915 VSS.t338 136.724
R3720 VSS.n12507 VSS.t626 136.724
R3721 VSS.n13099 VSS.t355 136.724
R3722 VSS.n13691 VSS.t416 136.724
R3723 VSS.n14283 VSS.t555 136.724
R3724 VSS.n14875 VSS.t7 136.724
R3725 VSS.n15467 VSS.t605 136.724
R3726 VSS.n6575 VSS.t139 136.724
R3727 VSS.n7172 VSS.t21 136.724
R3728 VSS.t389 VSS.n359 136.724
R3729 VSS.n905 VSS.t232 136.724
R3730 VSS.n1086 VSS.t422 136.724
R3731 VSS.n9547 VSS.t88 136.53
R3732 VSS.n17002 VSS.t523 130.508
R3733 VSS.n17416 VSS.t351 130.508
R3734 VSS.n9466 VSS.t477 130.508
R3735 VSS.n16408 VSS.t10 130.508
R3736 VSS.n1751 VSS.t344 130.508
R3737 VSS.n2001 VSS.t132 130.508
R3738 VSS.n2957 VSS.t591 130.508
R3739 VSS.n3549 VSS.t310 130.508
R3740 VSS.n4141 VSS.t212 130.508
R3741 VSS.n4733 VSS.t552 130.508
R3742 VSS.n2597 VSS.t91 130.508
R3743 VSS.n5558 VSS.t453 130.508
R3744 VSS.n6131 VSS.t219 130.508
R3745 VSS.n7690 VSS.t546 130.508
R3746 VSS.n8282 VSS.t483 130.508
R3747 VSS.n8874 VSS.t274 130.508
R3748 VSS.n10058 VSS.t124 130.508
R3749 VSS.n10650 VSS.t97 130.508
R3750 VSS.n11242 VSS.t203 130.508
R3751 VSS.n11834 VSS.t146 130.508
R3752 VSS.n12426 VSS.t252 130.508
R3753 VSS.n13018 VSS.t103 130.508
R3754 VSS.n13610 VSS.t446 130.508
R3755 VSS.n14202 VSS.t156 130.508
R3756 VSS.n14794 VSS.t159 130.508
R3757 VSS.n15386 VSS.t333 130.508
R3758 VSS.n6737 VSS.t480 130.508
R3759 VSS.n7097 VSS.t558 130.508
R3760 VSS.n200 VSS.t391 130.508
R3761 VSS.n18236 VSS.t298 130.508
R3762 VSS.n562 VSS.t573 130.508
R3763 VSS.n17529 VSS.n17525 128.415
R3764 VSS.n17527 VSS.n17458 128.415
R3765 VSS.n17558 VSS.n17458 128.415
R3766 VSS.n17562 VSS.n17561 128.415
R3767 VSS.n17591 VSS.n17590 128.415
R3768 VSS.n17911 VSS.n17910 121.799
R3769 VSS.n1406 VSS.n1341 121.799
R3770 VSS.n1253 VSS.n1212 112.246
R3771 VSS.n1255 VSS.n1208 112.246
R3772 VSS.n17926 VSS.n17925 106.575
R3773 VSS.t629 VSS.n1395 106.575
R3774 VSS.n17166 VSS.n16893 102.326
R3775 VSS.n17217 VSS.n17216 102.326
R3776 VSS.n17758 VSS.n17307 102.326
R3777 VSS.n17809 VSS.n17808 102.326
R3778 VSS.n9808 VSS.n9357 102.326
R3779 VSS.n9859 VSS.n9858 102.326
R3780 VSS.n16751 VSS.n16299 102.326
R3781 VSS.n16802 VSS.n16801 102.326
R3782 VSS.n16158 VSS.n1471 102.326
R3783 VSS.n16209 VSS.n16208 102.326
R3784 VSS.n2265 VSS.n2264 102.326
R3785 VSS.n2188 VSS.n2123 102.326
R3786 VSS.n3299 VSS.n2848 102.326
R3787 VSS.n3350 VSS.n3349 102.326
R3788 VSS.n3891 VSS.n3440 102.326
R3789 VSS.n3942 VSS.n3941 102.326
R3790 VSS.n4483 VSS.n4032 102.326
R3791 VSS.n4534 VSS.n4533 102.326
R3792 VSS.n5075 VSS.n4624 102.326
R3793 VSS.n5126 VSS.n5125 102.326
R3794 VSS.n5230 VSS.n5229 102.326
R3795 VSS.n2784 VSS.n2719 102.326
R3796 VSS.n5803 VSS.n5802 102.326
R3797 VSS.n5758 VSS.n5680 102.326
R3798 VSS.n6395 VSS.n6394 102.326
R3799 VSS.n6318 VSS.n6253 102.326
R3800 VSS.n8032 VSS.n7581 102.326
R3801 VSS.n8083 VSS.n8082 102.326
R3802 VSS.n8624 VSS.n8173 102.326
R3803 VSS.n8675 VSS.n8674 102.326
R3804 VSS.n9216 VSS.n8765 102.326
R3805 VSS.n9267 VSS.n9266 102.326
R3806 VSS.n10400 VSS.n9949 102.326
R3807 VSS.n10451 VSS.n10450 102.326
R3808 VSS.n10992 VSS.n10541 102.326
R3809 VSS.n11043 VSS.n11042 102.326
R3810 VSS.n11584 VSS.n11133 102.326
R3811 VSS.n11635 VSS.n11634 102.326
R3812 VSS.n12176 VSS.n11725 102.326
R3813 VSS.n12227 VSS.n12226 102.326
R3814 VSS.n12768 VSS.n12317 102.326
R3815 VSS.n12819 VSS.n12818 102.326
R3816 VSS.n13360 VSS.n12909 102.326
R3817 VSS.n13411 VSS.n13410 102.326
R3818 VSS.n13952 VSS.n13501 102.326
R3819 VSS.n14003 VSS.n14002 102.326
R3820 VSS.n14544 VSS.n14093 102.326
R3821 VSS.n14595 VSS.n14594 102.326
R3822 VSS.n15136 VSS.n14685 102.326
R3823 VSS.n15187 VSS.n15186 102.326
R3824 VSS.n15728 VSS.n15277 102.326
R3825 VSS.n15779 VSS.n15778 102.326
R3826 VSS.n15883 VSS.n15882 102.326
R3827 VSS.n6924 VSS.n6859 102.326
R3828 VSS.n7440 VSS.n6988 102.326
R3829 VSS.n7491 VSS.n7490 102.326
R3830 VSS.n18752 VSS.n86 102.326
R3831 VSS.n18803 VSS.n18802 102.326
R3832 VSS.n18383 VSS.n18382 102.326
R3833 VSS.n18495 VSS.n18494 102.326
R3834 VSS.n797 VSS.n796 102.326
R3835 VSS.n755 VSS.n682 102.326
R3836 VSS.n17927 VSS.t198 98.9624
R3837 VSS.n1246 VSS.n1245 97.2794
R3838 VSS.t584 VSS.n1271 97.2794
R3839 VSS.n10170 VSS.n10169 93.3527
R3840 VSS.n10201 VSS.n10200 93.3527
R3841 VSS.n17051 VSS.n17050 93.2208
R3842 VSS.n17052 VSS.n16953 93.2208
R3843 VSS.n17643 VSS.n17642 93.2208
R3844 VSS.n17644 VSS.n17367 93.2208
R3845 VSS.n18105 VSS.n18104 93.2208
R3846 VSS.n18136 VSS.n18135 93.2208
R3847 VSS.n9693 VSS.n9692 93.2208
R3848 VSS.n9694 VSS.n9417 93.2208
R3849 VSS.n16636 VSS.n16635 93.2208
R3850 VSS.n16637 VSS.n16359 93.2208
R3851 VSS.n16531 VSS.n16530 93.2208
R3852 VSS.n16532 VSS.n16434 93.2208
R3853 VSS.n16043 VSS.n16042 93.2208
R3854 VSS.n16044 VSS.n1531 93.2208
R3855 VSS.n1696 VSS.n1695 93.2208
R3856 VSS.n1697 VSS.n1599 93.2208
R3857 VSS.n2035 VSS.n1994 93.2208
R3858 VSS.n2037 VSS.n1990 93.2208
R3859 VSS.n1870 VSS.n1869 93.2208
R3860 VSS.n1901 VSS.n1900 93.2208
R3861 VSS.n3184 VSS.n3183 93.2208
R3862 VSS.n3185 VSS.n2908 93.2208
R3863 VSS.n3069 VSS.n3068 93.2208
R3864 VSS.n3100 VSS.n3099 93.2208
R3865 VSS.n3776 VSS.n3775 93.2208
R3866 VSS.n3777 VSS.n3500 93.2208
R3867 VSS.n3661 VSS.n3660 93.2208
R3868 VSS.n3692 VSS.n3691 93.2208
R3869 VSS.n4368 VSS.n4367 93.2208
R3870 VSS.n4369 VSS.n4092 93.2208
R3871 VSS.n4253 VSS.n4252 93.2208
R3872 VSS.n4284 VSS.n4283 93.2208
R3873 VSS.n4960 VSS.n4959 93.2208
R3874 VSS.n4961 VSS.n4684 93.2208
R3875 VSS.n4845 VSS.n4844 93.2208
R3876 VSS.n4876 VSS.n4875 93.2208
R3877 VSS.n2631 VSS.n2590 93.2208
R3878 VSS.n2633 VSS.n2586 93.2208
R3879 VSS.n2466 VSS.n2465 93.2208
R3880 VSS.n2497 VSS.n2496 93.2208
R3881 VSS.n5592 VSS.n5551 93.2208
R3882 VSS.n5594 VSS.n5547 93.2208
R3883 VSS.n5427 VSS.n5426 93.2208
R3884 VSS.n5458 VSS.n5457 93.2208
R3885 VSS.n6165 VSS.n6124 93.2208
R3886 VSS.n6167 VSS.n6120 93.2208
R3887 VSS.n6000 VSS.n5999 93.2208
R3888 VSS.n6031 VSS.n6030 93.2208
R3889 VSS.n7917 VSS.n7916 93.2208
R3890 VSS.n7918 VSS.n7641 93.2208
R3891 VSS.n7802 VSS.n7801 93.2208
R3892 VSS.n7833 VSS.n7832 93.2208
R3893 VSS.n8509 VSS.n8508 93.2208
R3894 VSS.n8510 VSS.n8233 93.2208
R3895 VSS.n8394 VSS.n8393 93.2208
R3896 VSS.n8425 VSS.n8424 93.2208
R3897 VSS.n9101 VSS.n9100 93.2208
R3898 VSS.n9102 VSS.n8825 93.2208
R3899 VSS.n8986 VSS.n8985 93.2208
R3900 VSS.n9017 VSS.n9016 93.2208
R3901 VSS.n10285 VSS.n10284 93.2208
R3902 VSS.n10286 VSS.n10009 93.2208
R3903 VSS.n10877 VSS.n10876 93.2208
R3904 VSS.n10878 VSS.n10601 93.2208
R3905 VSS.n10762 VSS.n10761 93.2208
R3906 VSS.n10793 VSS.n10792 93.2208
R3907 VSS.n11469 VSS.n11468 93.2208
R3908 VSS.n11470 VSS.n11193 93.2208
R3909 VSS.n11354 VSS.n11353 93.2208
R3910 VSS.n11385 VSS.n11384 93.2208
R3911 VSS.n12061 VSS.n12060 93.2208
R3912 VSS.n12062 VSS.n11785 93.2208
R3913 VSS.n11946 VSS.n11945 93.2208
R3914 VSS.n11977 VSS.n11976 93.2208
R3915 VSS.n12653 VSS.n12652 93.2208
R3916 VSS.n12654 VSS.n12377 93.2208
R3917 VSS.n12538 VSS.n12537 93.2208
R3918 VSS.n12569 VSS.n12568 93.2208
R3919 VSS.n13245 VSS.n13244 93.2208
R3920 VSS.n13246 VSS.n12969 93.2208
R3921 VSS.n13130 VSS.n13129 93.2208
R3922 VSS.n13161 VSS.n13160 93.2208
R3923 VSS.n13837 VSS.n13836 93.2208
R3924 VSS.n13838 VSS.n13561 93.2208
R3925 VSS.n13722 VSS.n13721 93.2208
R3926 VSS.n13753 VSS.n13752 93.2208
R3927 VSS.n14429 VSS.n14428 93.2208
R3928 VSS.n14430 VSS.n14153 93.2208
R3929 VSS.n14314 VSS.n14313 93.2208
R3930 VSS.n14345 VSS.n14344 93.2208
R3931 VSS.n15021 VSS.n15020 93.2208
R3932 VSS.n15022 VSS.n14745 93.2208
R3933 VSS.n14906 VSS.n14905 93.2208
R3934 VSS.n14937 VSS.n14936 93.2208
R3935 VSS.n15613 VSS.n15612 93.2208
R3936 VSS.n15614 VSS.n15337 93.2208
R3937 VSS.n15498 VSS.n15497 93.2208
R3938 VSS.n15529 VSS.n15528 93.2208
R3939 VSS.n6771 VSS.n6730 93.2208
R3940 VSS.n6773 VSS.n6726 93.2208
R3941 VSS.n6606 VSS.n6605 93.2208
R3942 VSS.n6637 VSS.n6636 93.2208
R3943 VSS.n7325 VSS.n7324 93.2208
R3944 VSS.n7326 VSS.n7048 93.2208
R3945 VSS.n7220 VSS.n7219 93.2208
R3946 VSS.n7221 VSS.n7123 93.2208
R3947 VSS.n18637 VSS.n18636 93.2208
R3948 VSS.n18638 VSS.n146 93.2208
R3949 VSS.n375 VSS.n374 93.2208
R3950 VSS.n383 VSS.n382 93.2208
R3951 VSS.n18270 VSS.n18229 93.2208
R3952 VSS.n18272 VSS.n18225 93.2208
R3953 VSS.n594 VSS.n550 93.2208
R3954 VSS.n596 VSS.n546 93.2208
R3955 VSS.n937 VSS.n898 93.2208
R3956 VSS.n939 VSS.n893 93.2208
R3957 VSS.n1118 VSS.n1079 93.2208
R3958 VSS.n1120 VSS.n1074 93.2208
R3959 VSS.n9578 VSS.n9577 93.0894
R3960 VSS.n9609 VSS.n9608 93.0894
R3961 VSS.n17941 VSS.n1293 91.35
R3962 VSS.n17876 VSS.n17875 91.35
R3963 VSS.n17165 VSS.n17164 89.5354
R3964 VSS.t173 VSS.n17236 89.5354
R3965 VSS.n17757 VSS.n17756 89.5354
R3966 VSS.t568 VSS.n17828 89.5354
R3967 VSS.n9807 VSS.n9806 89.5354
R3968 VSS.t449 VSS.n9878 89.5354
R3969 VSS.n16750 VSS.n16749 89.5354
R3970 VSS.t62 VSS.n16821 89.5354
R3971 VSS.n16157 VSS.n16156 89.5354
R3972 VSS.t512 VSS.n16228 89.5354
R3973 VSS.n2280 VSS.n2279 89.5354
R3974 VSS.t473 VSS.n2177 89.5354
R3975 VSS.n3298 VSS.n3297 89.5354
R3976 VSS.t575 VSS.n3369 89.5354
R3977 VSS.n3890 VSS.n3889 89.5354
R3978 VSS.t134 VSS.n3961 89.5354
R3979 VSS.n4482 VSS.n4481 89.5354
R3980 VSS.t269 VSS.n4553 89.5354
R3981 VSS.n5074 VSS.n5073 89.5354
R3982 VSS.t399 VSS.n5145 89.5354
R3983 VSS.n5245 VSS.n5244 89.5354
R3984 VSS.t505 VSS.n2773 89.5354
R3985 VSS.n5818 VSS.n5817 89.5354
R3986 VSS.t17 VSS.n5747 89.5354
R3987 VSS.n6410 VSS.n6409 89.5354
R3988 VSS.t31 VSS.n6307 89.5354
R3989 VSS.n8031 VSS.n8030 89.5354
R3990 VSS.t361 VSS.n8102 89.5354
R3991 VSS.n8623 VSS.n8622 89.5354
R3992 VSS.t494 VSS.n8694 89.5354
R3993 VSS.n9215 VSS.n9214 89.5354
R3994 VSS.t406 VSS.n9286 89.5354
R3995 VSS.n10399 VSS.n10398 89.5354
R3996 VSS.t378 VSS.n10470 89.5354
R3997 VSS.n10991 VSS.n10990 89.5354
R3998 VSS.t164 VSS.n11062 89.5354
R3999 VSS.n11583 VSS.n11582 89.5354
R4000 VSS.t58 VSS.n11654 89.5354
R4001 VSS.n12175 VSS.n12174 89.5354
R4002 VSS.t259 VSS.n12246 89.5354
R4003 VSS.n12767 VSS.n12766 89.5354
R4004 VSS.t441 VSS.n12838 89.5354
R4005 VSS.n13359 VSS.n13358 89.5354
R4006 VSS.t3 VSS.n13430 89.5354
R4007 VSS.n13951 VSS.n13950 89.5354
R4008 VSS.t460 VSS.n14022 89.5354
R4009 VSS.n14543 VSS.n14542 89.5354
R4010 VSS.t39 VSS.n14614 89.5354
R4011 VSS.n15135 VSS.n15134 89.5354
R4012 VSS.t152 VSS.n15206 89.5354
R4013 VSS.n15727 VSS.n15726 89.5354
R4014 VSS.t374 VSS.n15798 89.5354
R4015 VSS.n15898 VSS.n15897 89.5354
R4016 VSS.t113 VSS.n6913 89.5354
R4017 VSS.n7439 VSS.n7438 89.5354
R4018 VSS.t437 VSS.n7510 89.5354
R4019 VSS.n18751 VSS.n18750 89.5354
R4020 VSS.t182 VSS.n18822 89.5354
R4021 VSS.n18371 VSS.n18370 89.5354
R4022 VSS.t349 VSS.n18450 89.5354
R4023 VSS.n812 VSS.n811 89.5354
R4024 VSS.t335 VSS.n759 89.5354
R4025 VSS.t598 VSS.n16915 83.14
R4026 VSS.t120 VSS.n17329 83.14
R4027 VSS.t35 VSS.n9379 83.14
R4028 VSS.t490 VSS.n16321 83.14
R4029 VSS.t561 VSS.n1493 83.14
R4030 VSS.n2281 VSS.t78 83.14
R4031 VSS.t464 VSS.n2870 83.14
R4032 VSS.t611 VSS.n3462 83.14
R4033 VSS.t516 VSS.n4054 83.14
R4034 VSS.t176 VSS.n4646 83.14
R4035 VSS.n5246 VSS.t214 83.14
R4036 VSS.n5819 VSS.t116 83.14
R4037 VSS.n6411 VSS.t618 83.14
R4038 VSS.t239 VSS.n7603 83.14
R4039 VSS.t499 VSS.n8195 83.14
R4040 VSS.t541 VSS.n8787 83.14
R4041 VSS.t276 VSS.n9971 83.14
R4042 VSS.t587 VSS.n10563 83.14
R4043 VSS.t224 VSS.n11155 83.14
R4044 VSS.t306 VSS.n11747 83.14
R4045 VSS.t27 VSS.n12339 83.14
R4046 VSS.t328 VSS.n12931 83.14
R4047 VSS.t537 VSS.n13523 83.14
R4048 VSS.t316 VSS.n14115 83.14
R4049 VSS.t580 VSS.n14707 83.14
R4050 VSS.t594 VSS.n15299 83.14
R4051 VSS.n15899 VSS.t290 83.14
R4052 VSS.t431 VSS.n7010 83.14
R4053 VSS.t341 VSS.n108 83.14
R4054 VSS.n18369 VSS.t286 83.14
R4055 VSS.n813 VSS.t187 83.14
R4056 VSS.n1219 VSS.n1156 82.3134
R4057 VSS.n1287 VSS.n1286 82.3134
R4058 VSS.n17121 VSS.n17111 81.5708
R4059 VSS.n17113 VSS.n16916 81.5708
R4060 VSS.n17168 VSS.n16913 81.5708
R4061 VSS.n17235 VSS.n16882 81.5708
R4062 VSS.n17238 VSS.n16869 81.5708
R4063 VSS.n17265 VSS.n16866 81.5708
R4064 VSS.n17713 VSS.n17703 81.5708
R4065 VSS.n17705 VSS.n17330 81.5708
R4066 VSS.n17760 VSS.n17327 81.5708
R4067 VSS.n17827 VSS.n17296 81.5708
R4068 VSS.n17830 VSS.n17283 81.5708
R4069 VSS.n17857 VSS.n17280 81.5708
R4070 VSS.n18533 VSS.n18309 81.5708
R4071 VSS.n18368 VSS.n18311 81.5708
R4072 VSS.n18373 VSS.n18372 81.5708
R4073 VSS.n18449 VSS.n18385 81.5708
R4074 VSS.n18453 VSS.n18452 81.5708
R4075 VSS.n18461 VSS.n18437 81.5708
R4076 VSS.n9763 VSS.n9753 81.5708
R4077 VSS.n9755 VSS.n9380 81.5708
R4078 VSS.n9810 VSS.n9377 81.5708
R4079 VSS.n9877 VSS.n9346 81.5708
R4080 VSS.n9880 VSS.n9334 81.5708
R4081 VSS.n9908 VSS.n9331 81.5708
R4082 VSS.n16706 VSS.n16696 81.5708
R4083 VSS.n16698 VSS.n16322 81.5708
R4084 VSS.n16753 VSS.n16319 81.5708
R4085 VSS.n16820 VSS.n16288 81.5708
R4086 VSS.n16823 VSS.n16276 81.5708
R4087 VSS.n16851 VSS.n16273 81.5708
R4088 VSS.n16113 VSS.n16103 81.5708
R4089 VSS.n16105 VSS.n1494 81.5708
R4090 VSS.n16160 VSS.n1491 81.5708
R4091 VSS.n16227 VSS.n1460 81.5708
R4092 VSS.n16230 VSS.n1448 81.5708
R4093 VSS.n16258 VSS.n1445 81.5708
R4094 VSS.n2298 VSS.n2074 81.5708
R4095 VSS.n2282 VSS.n2076 81.5708
R4096 VSS.n2278 VSS.n2106 81.5708
R4097 VSS.n2191 VSS.n2190 81.5708
R4098 VSS.n2231 VSS.n2175 81.5708
R4099 VSS.n2227 VSS.n2198 81.5708
R4100 VSS.n3254 VSS.n3244 81.5708
R4101 VSS.n3246 VSS.n2871 81.5708
R4102 VSS.n3301 VSS.n2868 81.5708
R4103 VSS.n3368 VSS.n2837 81.5708
R4104 VSS.n3371 VSS.n2825 81.5708
R4105 VSS.n3399 VSS.n2822 81.5708
R4106 VSS.n3846 VSS.n3836 81.5708
R4107 VSS.n3838 VSS.n3463 81.5708
R4108 VSS.n3893 VSS.n3460 81.5708
R4109 VSS.n3960 VSS.n3429 81.5708
R4110 VSS.n3963 VSS.n3417 81.5708
R4111 VSS.n3991 VSS.n3414 81.5708
R4112 VSS.n4438 VSS.n4428 81.5708
R4113 VSS.n4430 VSS.n4055 81.5708
R4114 VSS.n4485 VSS.n4052 81.5708
R4115 VSS.n4552 VSS.n4021 81.5708
R4116 VSS.n4555 VSS.n4009 81.5708
R4117 VSS.n4583 VSS.n4006 81.5708
R4118 VSS.n5030 VSS.n5020 81.5708
R4119 VSS.n5022 VSS.n4647 81.5708
R4120 VSS.n5077 VSS.n4644 81.5708
R4121 VSS.n5144 VSS.n4613 81.5708
R4122 VSS.n5147 VSS.n4601 81.5708
R4123 VSS.n5175 VSS.n4598 81.5708
R4124 VSS.n5263 VSS.n2670 81.5708
R4125 VSS.n5247 VSS.n2672 81.5708
R4126 VSS.n5243 VSS.n2702 81.5708
R4127 VSS.n2787 VSS.n2786 81.5708
R4128 VSS.n5196 VSS.n2771 81.5708
R4129 VSS.n5192 VSS.n2794 81.5708
R4130 VSS.n5836 VSS.n5631 81.5708
R4131 VSS.n5820 VSS.n5633 81.5708
R4132 VSS.n5816 VSS.n5663 81.5708
R4133 VSS.n5761 VSS.n5760 81.5708
R4134 VSS.n5769 VSS.n5745 81.5708
R4135 VSS.n18881 VSS.n7 81.5708
R4136 VSS.n6428 VSS.n6204 81.5708
R4137 VSS.n6412 VSS.n6206 81.5708
R4138 VSS.n6408 VSS.n6236 81.5708
R4139 VSS.n6321 VSS.n6320 81.5708
R4140 VSS.n6361 VSS.n6305 81.5708
R4141 VSS.n6357 VSS.n6328 81.5708
R4142 VSS.n7987 VSS.n7977 81.5708
R4143 VSS.n7979 VSS.n7604 81.5708
R4144 VSS.n8034 VSS.n7601 81.5708
R4145 VSS.n8101 VSS.n7570 81.5708
R4146 VSS.n8104 VSS.n7558 81.5708
R4147 VSS.n8132 VSS.n7555 81.5708
R4148 VSS.n8579 VSS.n8569 81.5708
R4149 VSS.n8571 VSS.n8196 81.5708
R4150 VSS.n8626 VSS.n8193 81.5708
R4151 VSS.n8693 VSS.n8162 81.5708
R4152 VSS.n8696 VSS.n8150 81.5708
R4153 VSS.n8724 VSS.n8147 81.5708
R4154 VSS.n9171 VSS.n9161 81.5708
R4155 VSS.n9163 VSS.n8788 81.5708
R4156 VSS.n9218 VSS.n8785 81.5708
R4157 VSS.n9285 VSS.n8754 81.5708
R4158 VSS.n9288 VSS.n8742 81.5708
R4159 VSS.n9316 VSS.n8739 81.5708
R4160 VSS.n10355 VSS.n10345 81.5708
R4161 VSS.n10347 VSS.n9972 81.5708
R4162 VSS.n10402 VSS.n9969 81.5708
R4163 VSS.n10469 VSS.n9938 81.5708
R4164 VSS.n10472 VSS.n9926 81.5708
R4165 VSS.n10500 VSS.n9923 81.5708
R4166 VSS.n10947 VSS.n10937 81.5708
R4167 VSS.n10939 VSS.n10564 81.5708
R4168 VSS.n10994 VSS.n10561 81.5708
R4169 VSS.n11061 VSS.n10530 81.5708
R4170 VSS.n11064 VSS.n10518 81.5708
R4171 VSS.n11092 VSS.n10515 81.5708
R4172 VSS.n11539 VSS.n11529 81.5708
R4173 VSS.n11531 VSS.n11156 81.5708
R4174 VSS.n11586 VSS.n11153 81.5708
R4175 VSS.n11653 VSS.n11122 81.5708
R4176 VSS.n11656 VSS.n11110 81.5708
R4177 VSS.n11684 VSS.n11107 81.5708
R4178 VSS.n12131 VSS.n12121 81.5708
R4179 VSS.n12123 VSS.n11748 81.5708
R4180 VSS.n12178 VSS.n11745 81.5708
R4181 VSS.n12245 VSS.n11714 81.5708
R4182 VSS.n12248 VSS.n11702 81.5708
R4183 VSS.n12276 VSS.n11699 81.5708
R4184 VSS.n12723 VSS.n12713 81.5708
R4185 VSS.n12715 VSS.n12340 81.5708
R4186 VSS.n12770 VSS.n12337 81.5708
R4187 VSS.n12837 VSS.n12306 81.5708
R4188 VSS.n12840 VSS.n12294 81.5708
R4189 VSS.n12868 VSS.n12291 81.5708
R4190 VSS.n13315 VSS.n13305 81.5708
R4191 VSS.n13307 VSS.n12932 81.5708
R4192 VSS.n13362 VSS.n12929 81.5708
R4193 VSS.n13429 VSS.n12898 81.5708
R4194 VSS.n13432 VSS.n12886 81.5708
R4195 VSS.n13460 VSS.n12883 81.5708
R4196 VSS.n13907 VSS.n13897 81.5708
R4197 VSS.n13899 VSS.n13524 81.5708
R4198 VSS.n13954 VSS.n13521 81.5708
R4199 VSS.n14021 VSS.n13490 81.5708
R4200 VSS.n14024 VSS.n13478 81.5708
R4201 VSS.n14052 VSS.n13475 81.5708
R4202 VSS.n14499 VSS.n14489 81.5708
R4203 VSS.n14491 VSS.n14116 81.5708
R4204 VSS.n14546 VSS.n14113 81.5708
R4205 VSS.n14613 VSS.n14082 81.5708
R4206 VSS.n14616 VSS.n14070 81.5708
R4207 VSS.n14644 VSS.n14067 81.5708
R4208 VSS.n15091 VSS.n15081 81.5708
R4209 VSS.n15083 VSS.n14708 81.5708
R4210 VSS.n15138 VSS.n14705 81.5708
R4211 VSS.n15205 VSS.n14674 81.5708
R4212 VSS.n15208 VSS.n14662 81.5708
R4213 VSS.n15236 VSS.n14659 81.5708
R4214 VSS.n15683 VSS.n15673 81.5708
R4215 VSS.n15675 VSS.n15300 81.5708
R4216 VSS.n15730 VSS.n15297 81.5708
R4217 VSS.n15797 VSS.n15266 81.5708
R4218 VSS.n15800 VSS.n15254 81.5708
R4219 VSS.n15828 VSS.n15251 81.5708
R4220 VSS.n15916 VSS.n6810 81.5708
R4221 VSS.n15900 VSS.n6812 81.5708
R4222 VSS.n15896 VSS.n6842 81.5708
R4223 VSS.n6927 VSS.n6926 81.5708
R4224 VSS.n15849 VSS.n6911 81.5708
R4225 VSS.n15845 VSS.n6934 81.5708
R4226 VSS.n7395 VSS.n7385 81.5708
R4227 VSS.n7387 VSS.n7011 81.5708
R4228 VSS.n7442 VSS.n7008 81.5708
R4229 VSS.n7509 VSS.n6977 81.5708
R4230 VSS.n7512 VSS.n6965 81.5708
R4231 VSS.n7540 VSS.n6962 81.5708
R4232 VSS.n18707 VSS.n18697 81.5708
R4233 VSS.n18699 VSS.n109 81.5708
R4234 VSS.n18754 VSS.n106 81.5708
R4235 VSS.n18821 VSS.n75 81.5708
R4236 VSS.n18824 VSS.n63 81.5708
R4237 VSS.n18852 VSS.n60 81.5708
R4238 VSS.n830 VSS.n633 81.5708
R4239 VSS.n814 VSS.n635 81.5708
R4240 VSS.n810 VSS.n665 81.5708
R4241 VSS.n758 VSS.n757 81.5708
R4242 VSS.n761 VSS.n47 81.5708
R4243 VSS.n18873 VSS.n45 81.5708
R4244 VSS.n17944 VSS.n1292 81.5708
R4245 VSS.n17928 VSS.n1294 81.5708
R4246 VSS.n17924 VSS.n1324 81.5708
R4247 VSS.n1409 VSS.n1408 81.5708
R4248 VSS.n17877 VSS.n1393 81.5708
R4249 VSS.n17873 VSS.n1416 81.5708
R4250 VSS.n10167 VSS.n10166 80.9057
R4251 VSS.n10203 VSS.n10202 80.9057
R4252 VSS.n17030 VSS.n17029 80.7915
R4253 VSS.t247 VSS.n17082 80.7915
R4254 VSS.n17622 VSS.n17621 80.7915
R4255 VSS.t46 VSS.n17674 80.7915
R4256 VSS.n18102 VSS.n18101 80.7915
R4257 VSS.n18138 VSS.n18137 80.7915
R4258 VSS.n9672 VSS.n9671 80.7915
R4259 VSS.t65 VSS.n9724 80.7915
R4260 VSS.n16615 VSS.n16614 80.7915
R4261 VSS.t143 VSS.n16667 80.7915
R4262 VSS.n16510 VSS.n16509 80.7915
R4263 VSS.n16563 VSS.n16562 80.7915
R4264 VSS.n16022 VSS.n16021 80.7915
R4265 VSS.t455 VSS.n16074 80.7915
R4266 VSS.n1675 VSS.n1674 80.7915
R4267 VSS.n1728 VSS.n1727 80.7915
R4268 VSS.n2028 VSS.n2027 80.7915
R4269 VSS.t284 VSS.n2053 80.7915
R4270 VSS.n1867 VSS.n1866 80.7915
R4271 VSS.n1903 VSS.n1902 80.7915
R4272 VSS.n3163 VSS.n3162 80.7915
R4273 VSS.t313 VSS.n3215 80.7915
R4274 VSS.n3066 VSS.n3065 80.7915
R4275 VSS.n3102 VSS.n3101 80.7915
R4276 VSS.n3755 VSS.n3754 80.7915
R4277 VSS.t294 VSS.n3807 80.7915
R4278 VSS.n3658 VSS.n3657 80.7915
R4279 VSS.n3694 VSS.n3693 80.7915
R4280 VSS.n4347 VSS.n4346 80.7915
R4281 VSS.t75 VSS.n4399 80.7915
R4282 VSS.n4250 VSS.n4249 80.7915
R4283 VSS.n4286 VSS.n4285 80.7915
R4284 VSS.n4939 VSS.n4938 80.7915
R4285 VSS.t364 VSS.n4991 80.7915
R4286 VSS.n4842 VSS.n4841 80.7915
R4287 VSS.n4878 VSS.n4877 80.7915
R4288 VSS.n2624 VSS.n2623 80.7915
R4289 VSS.t549 VSS.n2649 80.7915
R4290 VSS.n2463 VSS.n2462 80.7915
R4291 VSS.n2499 VSS.n2498 80.7915
R4292 VSS.n5585 VSS.n5584 80.7915
R4293 VSS.t418 VSS.n5610 80.7915
R4294 VSS.n5424 VSS.n5423 80.7915
R4295 VSS.n5460 VSS.n5459 80.7915
R4296 VSS.n6158 VSS.n6157 80.7915
R4297 VSS.t81 VSS.n6183 80.7915
R4298 VSS.n5997 VSS.n5996 80.7915
R4299 VSS.n6033 VSS.n6032 80.7915
R4300 VSS.n7896 VSS.n7895 80.7915
R4301 VSS.t72 VSS.n7948 80.7915
R4302 VSS.n7799 VSS.n7798 80.7915
R4303 VSS.n7835 VSS.n7834 80.7915
R4304 VSS.n8488 VSS.n8487 80.7915
R4305 VSS.t93 VSS.n8540 80.7915
R4306 VSS.n8391 VSS.n8390 80.7915
R4307 VSS.n8427 VSS.n8426 80.7915
R4308 VSS.n9080 VSS.n9079 80.7915
R4309 VSS.t85 VSS.n9132 80.7915
R4310 VSS.n8983 VSS.n8982 80.7915
R4311 VSS.n9019 VSS.n9018 80.7915
R4312 VSS.n10264 VSS.n10263 80.7915
R4313 VSS.t100 VSS.n10316 80.7915
R4314 VSS.n10856 VSS.n10855 80.7915
R4315 VSS.t519 VSS.n10908 80.7915
R4316 VSS.n10759 VSS.n10758 80.7915
R4317 VSS.n10795 VSS.n10794 80.7915
R4318 VSS.n11448 VSS.n11447 80.7915
R4319 VSS.t395 VSS.n11500 80.7915
R4320 VSS.n11351 VSS.n11350 80.7915
R4321 VSS.n11387 VSS.n11386 80.7915
R4322 VSS.n12040 VSS.n12039 80.7915
R4323 VSS.t244 VSS.n12092 80.7915
R4324 VSS.n11943 VSS.n11942 80.7915
R4325 VSS.n11979 VSS.n11978 80.7915
R4326 VSS.n12632 VSS.n12631 80.7915
R4327 VSS.t221 VSS.n12684 80.7915
R4328 VSS.n12535 VSS.n12534 80.7915
R4329 VSS.n12571 VSS.n12570 80.7915
R4330 VSS.n13224 VSS.n13223 80.7915
R4331 VSS.t168 VSS.n13276 80.7915
R4332 VSS.n13127 VSS.n13126 80.7915
R4333 VSS.n13163 VSS.n13162 80.7915
R4334 VSS.n13816 VSS.n13815 80.7915
R4335 VSS.t43 VSS.n13868 80.7915
R4336 VSS.n13719 VSS.n13718 80.7915
R4337 VSS.n13755 VSS.n13754 80.7915
R4338 VSS.n14408 VSS.n14407 80.7915
R4339 VSS.t161 VSS.n14460 80.7915
R4340 VSS.n14311 VSS.n14310 80.7915
R4341 VSS.n14347 VSS.n14346 80.7915
R4342 VSS.n15000 VSS.n14999 80.7915
R4343 VSS.t525 VSS.n15052 80.7915
R4344 VSS.n14903 VSS.n14902 80.7915
R4345 VSS.n14939 VSS.n14938 80.7915
R4346 VSS.n15592 VSS.n15591 80.7915
R4347 VSS.t179 VSS.n15644 80.7915
R4348 VSS.n15495 VSS.n15494 80.7915
R4349 VSS.n15531 VSS.n15530 80.7915
R4350 VSS.n6764 VSS.n6763 80.7915
R4351 VSS.t413 VSS.n6789 80.7915
R4352 VSS.n6603 VSS.n6602 80.7915
R4353 VSS.n6639 VSS.n6638 80.7915
R4354 VSS.n7304 VSS.n7303 80.7915
R4355 VSS.t385 VSS.n7356 80.7915
R4356 VSS.n7199 VSS.n7198 80.7915
R4357 VSS.n7252 VSS.n7251 80.7915
R4358 VSS.n18616 VSS.n18615 80.7915
R4359 VSS.t129 VSS.n18668 80.7915
R4360 VSS.n361 VSS.n340 80.7915
R4361 VSS.n399 VSS.n330 80.7915
R4362 VSS.n18263 VSS.n18262 80.7915
R4363 VSS.t69 VSS.n18288 80.7915
R4364 VSS.n587 VSS.n586 80.7915
R4365 VSS.t126 VSS.n612 80.7915
R4366 VSS.n930 VSS.n929 80.7915
R4367 VSS.n956 VSS.n955 80.7915
R4368 VSS.n1111 VSS.n1110 80.7915
R4369 VSS.n1137 VSS.n1136 80.7915
R4370 VSS.n9575 VSS.n9574 80.6775
R4371 VSS.n9611 VSS.n9610 80.6775
R4372 VSS.n17214 VSS.n16894 80.0317
R4373 VSS.n17214 VSS.n16892 80.0317
R4374 VSS.n17806 VSS.n17308 80.0317
R4375 VSS.n17806 VSS.n17306 80.0317
R4376 VSS.n18497 VSS.n18359 80.0317
R4377 VSS.n18497 VSS.n18360 80.0317
R4378 VSS.n9856 VSS.n9358 80.0317
R4379 VSS.n9856 VSS.n9356 80.0317
R4380 VSS.n16799 VSS.n16300 80.0317
R4381 VSS.n16799 VSS.n16298 80.0317
R4382 VSS.n16206 VSS.n1472 80.0317
R4383 VSS.n16206 VSS.n1470 80.0317
R4384 VSS.n2262 VSS.n2122 80.0317
R4385 VSS.n2262 VSS.n2124 80.0317
R4386 VSS.n3347 VSS.n2849 80.0317
R4387 VSS.n3347 VSS.n2847 80.0317
R4388 VSS.n3939 VSS.n3441 80.0317
R4389 VSS.n3939 VSS.n3439 80.0317
R4390 VSS.n4531 VSS.n4033 80.0317
R4391 VSS.n4531 VSS.n4031 80.0317
R4392 VSS.n5123 VSS.n4625 80.0317
R4393 VSS.n5123 VSS.n4623 80.0317
R4394 VSS.n5227 VSS.n2718 80.0317
R4395 VSS.n5227 VSS.n2720 80.0317
R4396 VSS.n5800 VSS.n5679 80.0317
R4397 VSS.n5800 VSS.n5681 80.0317
R4398 VSS.n6392 VSS.n6252 80.0317
R4399 VSS.n6392 VSS.n6254 80.0317
R4400 VSS.n8080 VSS.n7582 80.0317
R4401 VSS.n8080 VSS.n7580 80.0317
R4402 VSS.n8672 VSS.n8174 80.0317
R4403 VSS.n8672 VSS.n8172 80.0317
R4404 VSS.n9264 VSS.n8766 80.0317
R4405 VSS.n9264 VSS.n8764 80.0317
R4406 VSS.n10448 VSS.n9950 80.0317
R4407 VSS.n10448 VSS.n9948 80.0317
R4408 VSS.n11040 VSS.n10542 80.0317
R4409 VSS.n11040 VSS.n10540 80.0317
R4410 VSS.n11632 VSS.n11134 80.0317
R4411 VSS.n11632 VSS.n11132 80.0317
R4412 VSS.n12224 VSS.n11726 80.0317
R4413 VSS.n12224 VSS.n11724 80.0317
R4414 VSS.n12816 VSS.n12318 80.0317
R4415 VSS.n12816 VSS.n12316 80.0317
R4416 VSS.n13408 VSS.n12910 80.0317
R4417 VSS.n13408 VSS.n12908 80.0317
R4418 VSS.n14000 VSS.n13502 80.0317
R4419 VSS.n14000 VSS.n13500 80.0317
R4420 VSS.n14592 VSS.n14094 80.0317
R4421 VSS.n14592 VSS.n14092 80.0317
R4422 VSS.n15184 VSS.n14686 80.0317
R4423 VSS.n15184 VSS.n14684 80.0317
R4424 VSS.n15776 VSS.n15278 80.0317
R4425 VSS.n15776 VSS.n15276 80.0317
R4426 VSS.n15880 VSS.n6858 80.0317
R4427 VSS.n15880 VSS.n6860 80.0317
R4428 VSS.n7488 VSS.n6989 80.0317
R4429 VSS.n7488 VSS.n6987 80.0317
R4430 VSS.n18800 VSS.n87 80.0317
R4431 VSS.n18800 VSS.n85 80.0317
R4432 VSS.n794 VSS.n681 80.0317
R4433 VSS.n794 VSS.n683 80.0317
R4434 VSS.n17908 VSS.n1340 80.0317
R4435 VSS.n17908 VSS.n1342 80.0317
R4436 VSS.n17118 VSS.n17112 76.7447
R4437 VSS.n17261 VSS.n16868 76.7447
R4438 VSS.n17710 VSS.n17704 76.7447
R4439 VSS.n17853 VSS.n17282 76.7447
R4440 VSS.n9760 VSS.n9754 76.7447
R4441 VSS.n9904 VSS.n9333 76.7447
R4442 VSS.n16703 VSS.n16697 76.7447
R4443 VSS.n16847 VSS.n16275 76.7447
R4444 VSS.n16110 VSS.n16104 76.7447
R4445 VSS.n16254 VSS.n1447 76.7447
R4446 VSS.n2295 VSS.n2075 76.7447
R4447 VSS.n2230 VSS.n2229 76.7447
R4448 VSS.n3251 VSS.n3245 76.7447
R4449 VSS.n3395 VSS.n2824 76.7447
R4450 VSS.n3843 VSS.n3837 76.7447
R4451 VSS.n3987 VSS.n3416 76.7447
R4452 VSS.n4435 VSS.n4429 76.7447
R4453 VSS.n4579 VSS.n4008 76.7447
R4454 VSS.n5027 VSS.n5021 76.7447
R4455 VSS.n5171 VSS.n4600 76.7447
R4456 VSS.n5260 VSS.n2671 76.7447
R4457 VSS.n5195 VSS.n5194 76.7447
R4458 VSS.n5833 VSS.n5632 76.7447
R4459 VSS.n5768 VSS.n5767 76.7447
R4460 VSS.n6425 VSS.n6205 76.7447
R4461 VSS.n6360 VSS.n6359 76.7447
R4462 VSS.n7984 VSS.n7978 76.7447
R4463 VSS.n8128 VSS.n7557 76.7447
R4464 VSS.n8576 VSS.n8570 76.7447
R4465 VSS.n8720 VSS.n8149 76.7447
R4466 VSS.n9168 VSS.n9162 76.7447
R4467 VSS.n9312 VSS.n8741 76.7447
R4468 VSS.n10352 VSS.n10346 76.7447
R4469 VSS.n10496 VSS.n9925 76.7447
R4470 VSS.n10944 VSS.n10938 76.7447
R4471 VSS.n11088 VSS.n10517 76.7447
R4472 VSS.n11536 VSS.n11530 76.7447
R4473 VSS.n11680 VSS.n11109 76.7447
R4474 VSS.n12128 VSS.n12122 76.7447
R4475 VSS.n12272 VSS.n11701 76.7447
R4476 VSS.n12720 VSS.n12714 76.7447
R4477 VSS.n12864 VSS.n12293 76.7447
R4478 VSS.n13312 VSS.n13306 76.7447
R4479 VSS.n13456 VSS.n12885 76.7447
R4480 VSS.n13904 VSS.n13898 76.7447
R4481 VSS.n14048 VSS.n13477 76.7447
R4482 VSS.n14496 VSS.n14490 76.7447
R4483 VSS.n14640 VSS.n14069 76.7447
R4484 VSS.n15088 VSS.n15082 76.7447
R4485 VSS.n15232 VSS.n14661 76.7447
R4486 VSS.n15680 VSS.n15674 76.7447
R4487 VSS.n15824 VSS.n15253 76.7447
R4488 VSS.n15913 VSS.n6811 76.7447
R4489 VSS.n15848 VSS.n15847 76.7447
R4490 VSS.n7392 VSS.n7386 76.7447
R4491 VSS.n7536 VSS.n6964 76.7447
R4492 VSS.n18704 VSS.n18698 76.7447
R4493 VSS.n18848 VSS.n62 76.7447
R4494 VSS.n18530 VSS.n18310 76.7447
R4495 VSS.n18457 VSS.n18439 76.7447
R4496 VSS.n827 VSS.n634 76.7447
R4497 VSS.n18870 VSS.n46 76.7447
R4498 VSS.n17943 VSS.n1288 76.1251
R4499 VSS.n1421 VSS.n1415 76.1251
R4500 VSS.t615 VSS.n17481 75.1106
R4501 VSS.n1220 VSS.n1218 74.5791
R4502 VSS.n1248 VSS.n1216 74.5791
R4503 VSS.n1252 VSS.n1211 74.5791
R4504 VSS.n1256 VSS.n1211 74.5791
R4505 VSS.n1269 VSS.n1207 74.5791
R4506 VSS.n1285 VSS.n1200 74.5791
R4507 VSS.n17495 VSS.n17482 74.5791
R4508 VSS.n17530 VSS.n17479 74.5791
R4509 VSS.n17526 VSS.n17459 74.5791
R4510 VSS.n17557 VSS.n17459 74.5791
R4511 VSS.n17563 VSS.n17457 74.5791
R4512 VSS.n17589 VSS.n17426 74.5791
R4513 VSS.n1087 VSS.n1085 74.5791
R4514 VSS.n1113 VSS.n1083 74.5791
R4515 VSS.n1117 VSS.n1078 74.5791
R4516 VSS.n1121 VSS.n1078 74.5791
R4517 VSS.n1134 VSS.n1073 74.5791
R4518 VSS.n1151 VSS.n1066 74.5791
R4519 VSS.n906 VSS.n904 74.5791
R4520 VSS.n932 VSS.n902 74.5791
R4521 VSS.n936 VSS.n897 74.5791
R4522 VSS.n940 VSS.n897 74.5791
R4523 VSS.n953 VSS.n892 74.5791
R4524 VSS.n970 VSS.n885 74.5791
R4525 VSS.n17027 VSS.n16989 74.5791
R4526 VSS.n17031 VSS.n16975 74.5791
R4527 VSS.n17054 VSS.n16972 74.5791
R4528 VSS.n17054 VSS.n16973 74.5791
R4529 VSS.n17080 VSS.n16952 74.5791
R4530 VSS.n17102 VSS.n16939 74.5791
R4531 VSS.n17619 VSS.n17403 74.5791
R4532 VSS.n17623 VSS.n17389 74.5791
R4533 VSS.n17646 VSS.n17386 74.5791
R4534 VSS.n17646 VSS.n17387 74.5791
R4535 VSS.n17672 VSS.n17366 74.5791
R4536 VSS.n17694 VSS.n17353 74.5791
R4537 VSS.n18237 VSS.n18235 74.5791
R4538 VSS.n18265 VSS.n18233 74.5791
R4539 VSS.n18269 VSS.n18228 74.5791
R4540 VSS.n18273 VSS.n18228 74.5791
R4541 VSS.n18286 VSS.n18224 74.5791
R4542 VSS.n18302 VSS.n18217 74.5791
R4543 VSS.n287 VSS.n274 74.5791
R4544 VSS.n18107 VSS.n271 74.5791
R4545 VSS.n18103 VSS.n251 74.5791
R4546 VSS.n18134 VSS.n251 74.5791
R4547 VSS.n18140 VSS.n249 74.5791
R4548 VSS.n18166 VSS.n218 74.5791
R4549 VSS.n9545 VSS.n9532 74.5791
R4550 VSS.n9580 VSS.n9529 74.5791
R4551 VSS.n9576 VSS.n9509 74.5791
R4552 VSS.n9607 VSS.n9509 74.5791
R4553 VSS.n9613 VSS.n9507 74.5791
R4554 VSS.n9639 VSS.n9476 74.5791
R4555 VSS.n9669 VSS.n9453 74.5791
R4556 VSS.n9673 VSS.n9439 74.5791
R4557 VSS.n9696 VSS.n9436 74.5791
R4558 VSS.n9696 VSS.n9437 74.5791
R4559 VSS.n9722 VSS.n9416 74.5791
R4560 VSS.n9744 VSS.n9403 74.5791
R4561 VSS.n16507 VSS.n16470 74.5791
R4562 VSS.n16511 VSS.n16458 74.5791
R4563 VSS.n16534 VSS.n16455 74.5791
R4564 VSS.n16534 VSS.n16456 74.5791
R4565 VSS.n16560 VSS.n16433 74.5791
R4566 VSS.n16583 VSS.n16420 74.5791
R4567 VSS.n16612 VSS.n16395 74.5791
R4568 VSS.n16616 VSS.n16381 74.5791
R4569 VSS.n16639 VSS.n16378 74.5791
R4570 VSS.n16639 VSS.n16379 74.5791
R4571 VSS.n16665 VSS.n16358 74.5791
R4572 VSS.n16687 VSS.n16345 74.5791
R4573 VSS.n1672 VSS.n1635 74.5791
R4574 VSS.n1676 VSS.n1623 74.5791
R4575 VSS.n1699 VSS.n1620 74.5791
R4576 VSS.n1699 VSS.n1621 74.5791
R4577 VSS.n1725 VSS.n1598 74.5791
R4578 VSS.n1748 VSS.n1585 74.5791
R4579 VSS.n16019 VSS.n1567 74.5791
R4580 VSS.n16023 VSS.n1553 74.5791
R4581 VSS.n16046 VSS.n1550 74.5791
R4582 VSS.n16046 VSS.n1551 74.5791
R4583 VSS.n16072 VSS.n1530 74.5791
R4584 VSS.n16094 VSS.n1517 74.5791
R4585 VSS.n1837 VSS.n1824 74.5791
R4586 VSS.n1872 VSS.n1821 74.5791
R4587 VSS.n1868 VSS.n1801 74.5791
R4588 VSS.n1899 VSS.n1801 74.5791
R4589 VSS.n1905 VSS.n1799 74.5791
R4590 VSS.n1931 VSS.n1768 74.5791
R4591 VSS.n2002 VSS.n2000 74.5791
R4592 VSS.n2030 VSS.n1998 74.5791
R4593 VSS.n2034 VSS.n1993 74.5791
R4594 VSS.n2038 VSS.n1993 74.5791
R4595 VSS.n2051 VSS.n1989 74.5791
R4596 VSS.n2067 VSS.n1982 74.5791
R4597 VSS.n3036 VSS.n3023 74.5791
R4598 VSS.n3071 VSS.n3020 74.5791
R4599 VSS.n3067 VSS.n3000 74.5791
R4600 VSS.n3098 VSS.n3000 74.5791
R4601 VSS.n3104 VSS.n2998 74.5791
R4602 VSS.n3130 VSS.n2967 74.5791
R4603 VSS.n3160 VSS.n2944 74.5791
R4604 VSS.n3164 VSS.n2930 74.5791
R4605 VSS.n3187 VSS.n2927 74.5791
R4606 VSS.n3187 VSS.n2928 74.5791
R4607 VSS.n3213 VSS.n2907 74.5791
R4608 VSS.n3235 VSS.n2894 74.5791
R4609 VSS.n3628 VSS.n3615 74.5791
R4610 VSS.n3663 VSS.n3612 74.5791
R4611 VSS.n3659 VSS.n3592 74.5791
R4612 VSS.n3690 VSS.n3592 74.5791
R4613 VSS.n3696 VSS.n3590 74.5791
R4614 VSS.n3722 VSS.n3559 74.5791
R4615 VSS.n3752 VSS.n3536 74.5791
R4616 VSS.n3756 VSS.n3522 74.5791
R4617 VSS.n3779 VSS.n3519 74.5791
R4618 VSS.n3779 VSS.n3520 74.5791
R4619 VSS.n3805 VSS.n3499 74.5791
R4620 VSS.n3827 VSS.n3486 74.5791
R4621 VSS.n4220 VSS.n4207 74.5791
R4622 VSS.n4255 VSS.n4204 74.5791
R4623 VSS.n4251 VSS.n4184 74.5791
R4624 VSS.n4282 VSS.n4184 74.5791
R4625 VSS.n4288 VSS.n4182 74.5791
R4626 VSS.n4314 VSS.n4151 74.5791
R4627 VSS.n4344 VSS.n4128 74.5791
R4628 VSS.n4348 VSS.n4114 74.5791
R4629 VSS.n4371 VSS.n4111 74.5791
R4630 VSS.n4371 VSS.n4112 74.5791
R4631 VSS.n4397 VSS.n4091 74.5791
R4632 VSS.n4419 VSS.n4078 74.5791
R4633 VSS.n4812 VSS.n4799 74.5791
R4634 VSS.n4847 VSS.n4796 74.5791
R4635 VSS.n4843 VSS.n4776 74.5791
R4636 VSS.n4874 VSS.n4776 74.5791
R4637 VSS.n4880 VSS.n4774 74.5791
R4638 VSS.n4906 VSS.n4743 74.5791
R4639 VSS.n4936 VSS.n4720 74.5791
R4640 VSS.n4940 VSS.n4706 74.5791
R4641 VSS.n4963 VSS.n4703 74.5791
R4642 VSS.n4963 VSS.n4704 74.5791
R4643 VSS.n4989 VSS.n4683 74.5791
R4644 VSS.n5011 VSS.n4670 74.5791
R4645 VSS.n2433 VSS.n2420 74.5791
R4646 VSS.n2468 VSS.n2417 74.5791
R4647 VSS.n2464 VSS.n2397 74.5791
R4648 VSS.n2495 VSS.n2397 74.5791
R4649 VSS.n2501 VSS.n2395 74.5791
R4650 VSS.n2527 VSS.n2364 74.5791
R4651 VSS.n2598 VSS.n2596 74.5791
R4652 VSS.n2626 VSS.n2594 74.5791
R4653 VSS.n2630 VSS.n2589 74.5791
R4654 VSS.n2634 VSS.n2589 74.5791
R4655 VSS.n2647 VSS.n2585 74.5791
R4656 VSS.n2663 VSS.n2578 74.5791
R4657 VSS.n5394 VSS.n5381 74.5791
R4658 VSS.n5429 VSS.n5378 74.5791
R4659 VSS.n5425 VSS.n5358 74.5791
R4660 VSS.n5456 VSS.n5358 74.5791
R4661 VSS.n5462 VSS.n5356 74.5791
R4662 VSS.n5488 VSS.n5325 74.5791
R4663 VSS.n5559 VSS.n5557 74.5791
R4664 VSS.n5587 VSS.n5555 74.5791
R4665 VSS.n5591 VSS.n5550 74.5791
R4666 VSS.n5595 VSS.n5550 74.5791
R4667 VSS.n5608 VSS.n5546 74.5791
R4668 VSS.n5624 VSS.n5539 74.5791
R4669 VSS.n5967 VSS.n5954 74.5791
R4670 VSS.n6002 VSS.n5951 74.5791
R4671 VSS.n5998 VSS.n5931 74.5791
R4672 VSS.n6029 VSS.n5931 74.5791
R4673 VSS.n6035 VSS.n5929 74.5791
R4674 VSS.n6061 VSS.n5898 74.5791
R4675 VSS.n6132 VSS.n6130 74.5791
R4676 VSS.n6160 VSS.n6128 74.5791
R4677 VSS.n6164 VSS.n6123 74.5791
R4678 VSS.n6168 VSS.n6123 74.5791
R4679 VSS.n6181 VSS.n6119 74.5791
R4680 VSS.n6197 VSS.n6112 74.5791
R4681 VSS.n7769 VSS.n7756 74.5791
R4682 VSS.n7804 VSS.n7753 74.5791
R4683 VSS.n7800 VSS.n7733 74.5791
R4684 VSS.n7831 VSS.n7733 74.5791
R4685 VSS.n7837 VSS.n7731 74.5791
R4686 VSS.n7863 VSS.n7700 74.5791
R4687 VSS.n7893 VSS.n7677 74.5791
R4688 VSS.n7897 VSS.n7663 74.5791
R4689 VSS.n7920 VSS.n7660 74.5791
R4690 VSS.n7920 VSS.n7661 74.5791
R4691 VSS.n7946 VSS.n7640 74.5791
R4692 VSS.n7968 VSS.n7627 74.5791
R4693 VSS.n8361 VSS.n8348 74.5791
R4694 VSS.n8396 VSS.n8345 74.5791
R4695 VSS.n8392 VSS.n8325 74.5791
R4696 VSS.n8423 VSS.n8325 74.5791
R4697 VSS.n8429 VSS.n8323 74.5791
R4698 VSS.n8455 VSS.n8292 74.5791
R4699 VSS.n8485 VSS.n8269 74.5791
R4700 VSS.n8489 VSS.n8255 74.5791
R4701 VSS.n8512 VSS.n8252 74.5791
R4702 VSS.n8512 VSS.n8253 74.5791
R4703 VSS.n8538 VSS.n8232 74.5791
R4704 VSS.n8560 VSS.n8219 74.5791
R4705 VSS.n8953 VSS.n8940 74.5791
R4706 VSS.n8988 VSS.n8937 74.5791
R4707 VSS.n8984 VSS.n8917 74.5791
R4708 VSS.n9015 VSS.n8917 74.5791
R4709 VSS.n9021 VSS.n8915 74.5791
R4710 VSS.n9047 VSS.n8884 74.5791
R4711 VSS.n9077 VSS.n8861 74.5791
R4712 VSS.n9081 VSS.n8847 74.5791
R4713 VSS.n9104 VSS.n8844 74.5791
R4714 VSS.n9104 VSS.n8845 74.5791
R4715 VSS.n9130 VSS.n8824 74.5791
R4716 VSS.n9152 VSS.n8811 74.5791
R4717 VSS.n10137 VSS.n10124 74.5791
R4718 VSS.n10172 VSS.n10121 74.5791
R4719 VSS.n10168 VSS.n10101 74.5791
R4720 VSS.n10199 VSS.n10101 74.5791
R4721 VSS.n10205 VSS.n10099 74.5791
R4722 VSS.n10231 VSS.n10068 74.5791
R4723 VSS.n10261 VSS.n10045 74.5791
R4724 VSS.n10265 VSS.n10031 74.5791
R4725 VSS.n10288 VSS.n10028 74.5791
R4726 VSS.n10288 VSS.n10029 74.5791
R4727 VSS.n10314 VSS.n10008 74.5791
R4728 VSS.n10336 VSS.n9995 74.5791
R4729 VSS.n10729 VSS.n10716 74.5791
R4730 VSS.n10764 VSS.n10713 74.5791
R4731 VSS.n10760 VSS.n10693 74.5791
R4732 VSS.n10791 VSS.n10693 74.5791
R4733 VSS.n10797 VSS.n10691 74.5791
R4734 VSS.n10823 VSS.n10660 74.5791
R4735 VSS.n10853 VSS.n10637 74.5791
R4736 VSS.n10857 VSS.n10623 74.5791
R4737 VSS.n10880 VSS.n10620 74.5791
R4738 VSS.n10880 VSS.n10621 74.5791
R4739 VSS.n10906 VSS.n10600 74.5791
R4740 VSS.n10928 VSS.n10587 74.5791
R4741 VSS.n11321 VSS.n11308 74.5791
R4742 VSS.n11356 VSS.n11305 74.5791
R4743 VSS.n11352 VSS.n11285 74.5791
R4744 VSS.n11383 VSS.n11285 74.5791
R4745 VSS.n11389 VSS.n11283 74.5791
R4746 VSS.n11415 VSS.n11252 74.5791
R4747 VSS.n11445 VSS.n11229 74.5791
R4748 VSS.n11449 VSS.n11215 74.5791
R4749 VSS.n11472 VSS.n11212 74.5791
R4750 VSS.n11472 VSS.n11213 74.5791
R4751 VSS.n11498 VSS.n11192 74.5791
R4752 VSS.n11520 VSS.n11179 74.5791
R4753 VSS.n11913 VSS.n11900 74.5791
R4754 VSS.n11948 VSS.n11897 74.5791
R4755 VSS.n11944 VSS.n11877 74.5791
R4756 VSS.n11975 VSS.n11877 74.5791
R4757 VSS.n11981 VSS.n11875 74.5791
R4758 VSS.n12007 VSS.n11844 74.5791
R4759 VSS.n12037 VSS.n11821 74.5791
R4760 VSS.n12041 VSS.n11807 74.5791
R4761 VSS.n12064 VSS.n11804 74.5791
R4762 VSS.n12064 VSS.n11805 74.5791
R4763 VSS.n12090 VSS.n11784 74.5791
R4764 VSS.n12112 VSS.n11771 74.5791
R4765 VSS.n12505 VSS.n12492 74.5791
R4766 VSS.n12540 VSS.n12489 74.5791
R4767 VSS.n12536 VSS.n12469 74.5791
R4768 VSS.n12567 VSS.n12469 74.5791
R4769 VSS.n12573 VSS.n12467 74.5791
R4770 VSS.n12599 VSS.n12436 74.5791
R4771 VSS.n12629 VSS.n12413 74.5791
R4772 VSS.n12633 VSS.n12399 74.5791
R4773 VSS.n12656 VSS.n12396 74.5791
R4774 VSS.n12656 VSS.n12397 74.5791
R4775 VSS.n12682 VSS.n12376 74.5791
R4776 VSS.n12704 VSS.n12363 74.5791
R4777 VSS.n13097 VSS.n13084 74.5791
R4778 VSS.n13132 VSS.n13081 74.5791
R4779 VSS.n13128 VSS.n13061 74.5791
R4780 VSS.n13159 VSS.n13061 74.5791
R4781 VSS.n13165 VSS.n13059 74.5791
R4782 VSS.n13191 VSS.n13028 74.5791
R4783 VSS.n13221 VSS.n13005 74.5791
R4784 VSS.n13225 VSS.n12991 74.5791
R4785 VSS.n13248 VSS.n12988 74.5791
R4786 VSS.n13248 VSS.n12989 74.5791
R4787 VSS.n13274 VSS.n12968 74.5791
R4788 VSS.n13296 VSS.n12955 74.5791
R4789 VSS.n13689 VSS.n13676 74.5791
R4790 VSS.n13724 VSS.n13673 74.5791
R4791 VSS.n13720 VSS.n13653 74.5791
R4792 VSS.n13751 VSS.n13653 74.5791
R4793 VSS.n13757 VSS.n13651 74.5791
R4794 VSS.n13783 VSS.n13620 74.5791
R4795 VSS.n13813 VSS.n13597 74.5791
R4796 VSS.n13817 VSS.n13583 74.5791
R4797 VSS.n13840 VSS.n13580 74.5791
R4798 VSS.n13840 VSS.n13581 74.5791
R4799 VSS.n13866 VSS.n13560 74.5791
R4800 VSS.n13888 VSS.n13547 74.5791
R4801 VSS.n14281 VSS.n14268 74.5791
R4802 VSS.n14316 VSS.n14265 74.5791
R4803 VSS.n14312 VSS.n14245 74.5791
R4804 VSS.n14343 VSS.n14245 74.5791
R4805 VSS.n14349 VSS.n14243 74.5791
R4806 VSS.n14375 VSS.n14212 74.5791
R4807 VSS.n14405 VSS.n14189 74.5791
R4808 VSS.n14409 VSS.n14175 74.5791
R4809 VSS.n14432 VSS.n14172 74.5791
R4810 VSS.n14432 VSS.n14173 74.5791
R4811 VSS.n14458 VSS.n14152 74.5791
R4812 VSS.n14480 VSS.n14139 74.5791
R4813 VSS.n14873 VSS.n14860 74.5791
R4814 VSS.n14908 VSS.n14857 74.5791
R4815 VSS.n14904 VSS.n14837 74.5791
R4816 VSS.n14935 VSS.n14837 74.5791
R4817 VSS.n14941 VSS.n14835 74.5791
R4818 VSS.n14967 VSS.n14804 74.5791
R4819 VSS.n14997 VSS.n14781 74.5791
R4820 VSS.n15001 VSS.n14767 74.5791
R4821 VSS.n15024 VSS.n14764 74.5791
R4822 VSS.n15024 VSS.n14765 74.5791
R4823 VSS.n15050 VSS.n14744 74.5791
R4824 VSS.n15072 VSS.n14731 74.5791
R4825 VSS.n15465 VSS.n15452 74.5791
R4826 VSS.n15500 VSS.n15449 74.5791
R4827 VSS.n15496 VSS.n15429 74.5791
R4828 VSS.n15527 VSS.n15429 74.5791
R4829 VSS.n15533 VSS.n15427 74.5791
R4830 VSS.n15559 VSS.n15396 74.5791
R4831 VSS.n15589 VSS.n15373 74.5791
R4832 VSS.n15593 VSS.n15359 74.5791
R4833 VSS.n15616 VSS.n15356 74.5791
R4834 VSS.n15616 VSS.n15357 74.5791
R4835 VSS.n15642 VSS.n15336 74.5791
R4836 VSS.n15664 VSS.n15323 74.5791
R4837 VSS.n6573 VSS.n6560 74.5791
R4838 VSS.n6608 VSS.n6557 74.5791
R4839 VSS.n6604 VSS.n6537 74.5791
R4840 VSS.n6635 VSS.n6537 74.5791
R4841 VSS.n6641 VSS.n6535 74.5791
R4842 VSS.n6667 VSS.n6504 74.5791
R4843 VSS.n6738 VSS.n6736 74.5791
R4844 VSS.n6766 VSS.n6734 74.5791
R4845 VSS.n6770 VSS.n6729 74.5791
R4846 VSS.n6774 VSS.n6729 74.5791
R4847 VSS.n6787 VSS.n6725 74.5791
R4848 VSS.n6803 VSS.n6718 74.5791
R4849 VSS.n7196 VSS.n7159 74.5791
R4850 VSS.n7200 VSS.n7147 74.5791
R4851 VSS.n7223 VSS.n7144 74.5791
R4852 VSS.n7223 VSS.n7145 74.5791
R4853 VSS.n7249 VSS.n7122 74.5791
R4854 VSS.n7272 VSS.n7109 74.5791
R4855 VSS.n7301 VSS.n7084 74.5791
R4856 VSS.n7305 VSS.n7070 74.5791
R4857 VSS.n7328 VSS.n7067 74.5791
R4858 VSS.n7328 VSS.n7068 74.5791
R4859 VSS.n7354 VSS.n7047 74.5791
R4860 VSS.n7376 VSS.n7034 74.5791
R4861 VSS.n358 VSS.n344 74.5791
R4862 VSS.n372 VSS.n341 74.5791
R4863 VSS.n376 VSS.n337 74.5791
R4864 VSS.n381 VSS.n337 74.5791
R4865 VSS.n385 VSS.n331 74.5791
R4866 VSS.n402 VSS.n329 74.5791
R4867 VSS.n18613 VSS.n182 74.5791
R4868 VSS.n18617 VSS.n168 74.5791
R4869 VSS.n18640 VSS.n165 74.5791
R4870 VSS.n18640 VSS.n166 74.5791
R4871 VSS.n18666 VSS.n145 74.5791
R4872 VSS.n18688 VSS.n132 74.5791
R4873 VSS.n563 VSS.n556 74.5791
R4874 VSS.n589 VSS.n554 74.5791
R4875 VSS.n593 VSS.n549 74.5791
R4876 VSS.n597 VSS.n549 74.5791
R4877 VSS.n610 VSS.n545 74.5791
R4878 VSS.n626 VSS.n538 74.5791
R4879 VSS.n10140 VSS.n10139 68.4588
R4880 VSS.n10234 VSS.n10233 68.4588
R4881 VSS.n17003 VSS.n17002 68.3621
R4882 VSS.n17104 VSS.n17103 68.3621
R4883 VSS.n17417 VSS.n17416 68.3621
R4884 VSS.n17696 VSS.n17695 68.3621
R4885 VSS.n18075 VSS.n18074 68.3621
R4886 VSS.n18169 VSS.n18168 68.3621
R4887 VSS.n9467 VSS.n9466 68.3621
R4888 VSS.n9746 VSS.n9745 68.3621
R4889 VSS.n16409 VSS.n16408 68.3621
R4890 VSS.n16689 VSS.n16688 68.3621
R4891 VSS.n16484 VSS.n16483 68.3621
R4892 VSS.n16585 VSS.n16584 68.3621
R4893 VSS.n1752 VSS.n1751 68.3621
R4894 VSS.n16096 VSS.n16095 68.3621
R4895 VSS.n1649 VSS.n1648 68.3621
R4896 VSS.n1750 VSS.n1749 68.3621
R4897 VSS.n2001 VSS.n1759 68.3621
R4898 VSS.n2069 VSS.n2068 68.3621
R4899 VSS.n1840 VSS.n1839 68.3621
R4900 VSS.n1934 VSS.n1933 68.3621
R4901 VSS.n2958 VSS.n2957 68.3621
R4902 VSS.n3237 VSS.n3236 68.3621
R4903 VSS.n3039 VSS.n3038 68.3621
R4904 VSS.n3133 VSS.n3132 68.3621
R4905 VSS.n3550 VSS.n3549 68.3621
R4906 VSS.n3829 VSS.n3828 68.3621
R4907 VSS.n3631 VSS.n3630 68.3621
R4908 VSS.n3725 VSS.n3724 68.3621
R4909 VSS.n4142 VSS.n4141 68.3621
R4910 VSS.n4421 VSS.n4420 68.3621
R4911 VSS.n4223 VSS.n4222 68.3621
R4912 VSS.n4317 VSS.n4316 68.3621
R4913 VSS.n4734 VSS.n4733 68.3621
R4914 VSS.n5013 VSS.n5012 68.3621
R4915 VSS.n4815 VSS.n4814 68.3621
R4916 VSS.n4909 VSS.n4908 68.3621
R4917 VSS.n2597 VSS.n2355 68.3621
R4918 VSS.n2665 VSS.n2664 68.3621
R4919 VSS.n2436 VSS.n2435 68.3621
R4920 VSS.n2530 VSS.n2529 68.3621
R4921 VSS.n5558 VSS.n5316 68.3621
R4922 VSS.n5626 VSS.n5625 68.3621
R4923 VSS.n5397 VSS.n5396 68.3621
R4924 VSS.n5491 VSS.n5490 68.3621
R4925 VSS.n6131 VSS.n5889 68.3621
R4926 VSS.n6199 VSS.n6198 68.3621
R4927 VSS.n5970 VSS.n5969 68.3621
R4928 VSS.n6064 VSS.n6063 68.3621
R4929 VSS.n7691 VSS.n7690 68.3621
R4930 VSS.n7970 VSS.n7969 68.3621
R4931 VSS.n7772 VSS.n7771 68.3621
R4932 VSS.n7866 VSS.n7865 68.3621
R4933 VSS.n8283 VSS.n8282 68.3621
R4934 VSS.n8562 VSS.n8561 68.3621
R4935 VSS.n8364 VSS.n8363 68.3621
R4936 VSS.n8458 VSS.n8457 68.3621
R4937 VSS.n8875 VSS.n8874 68.3621
R4938 VSS.n9154 VSS.n9153 68.3621
R4939 VSS.n8956 VSS.n8955 68.3621
R4940 VSS.n9050 VSS.n9049 68.3621
R4941 VSS.n10059 VSS.n10058 68.3621
R4942 VSS.n10338 VSS.n10337 68.3621
R4943 VSS.n10651 VSS.n10650 68.3621
R4944 VSS.n10930 VSS.n10929 68.3621
R4945 VSS.n10732 VSS.n10731 68.3621
R4946 VSS.n10826 VSS.n10825 68.3621
R4947 VSS.n11243 VSS.n11242 68.3621
R4948 VSS.n11522 VSS.n11521 68.3621
R4949 VSS.n11324 VSS.n11323 68.3621
R4950 VSS.n11418 VSS.n11417 68.3621
R4951 VSS.n11835 VSS.n11834 68.3621
R4952 VSS.n12114 VSS.n12113 68.3621
R4953 VSS.n11916 VSS.n11915 68.3621
R4954 VSS.n12010 VSS.n12009 68.3621
R4955 VSS.n12427 VSS.n12426 68.3621
R4956 VSS.n12706 VSS.n12705 68.3621
R4957 VSS.n12508 VSS.n12507 68.3621
R4958 VSS.n12602 VSS.n12601 68.3621
R4959 VSS.n13019 VSS.n13018 68.3621
R4960 VSS.n13298 VSS.n13297 68.3621
R4961 VSS.n13100 VSS.n13099 68.3621
R4962 VSS.n13194 VSS.n13193 68.3621
R4963 VSS.n13611 VSS.n13610 68.3621
R4964 VSS.n13890 VSS.n13889 68.3621
R4965 VSS.n13692 VSS.n13691 68.3621
R4966 VSS.n13786 VSS.n13785 68.3621
R4967 VSS.n14203 VSS.n14202 68.3621
R4968 VSS.n14482 VSS.n14481 68.3621
R4969 VSS.n14284 VSS.n14283 68.3621
R4970 VSS.n14378 VSS.n14377 68.3621
R4971 VSS.n14795 VSS.n14794 68.3621
R4972 VSS.n15074 VSS.n15073 68.3621
R4973 VSS.n14876 VSS.n14875 68.3621
R4974 VSS.n14970 VSS.n14969 68.3621
R4975 VSS.n15387 VSS.n15386 68.3621
R4976 VSS.n15666 VSS.n15665 68.3621
R4977 VSS.n15468 VSS.n15467 68.3621
R4978 VSS.n15562 VSS.n15561 68.3621
R4979 VSS.n6737 VSS.n6495 68.3621
R4980 VSS.n6805 VSS.n6804 68.3621
R4981 VSS.n6576 VSS.n6575 68.3621
R4982 VSS.n6670 VSS.n6669 68.3621
R4983 VSS.n7098 VSS.n7097 68.3621
R4984 VSS.n7378 VSS.n7377 68.3621
R4985 VSS.n7173 VSS.n7172 68.3621
R4986 VSS.n7274 VSS.n7273 68.3621
R4987 VSS.n201 VSS.n200 68.3621
R4988 VSS.n18690 VSS.n18689 68.3621
R4989 VSS.n359 VSS.n288 68.3621
R4990 VSS.n401 VSS.n199 68.3621
R4991 VSS.n18236 VSS.n209 68.3621
R4992 VSS.n18304 VSS.n18303 68.3621
R4993 VSS.n562 VSS.n561 68.3621
R4994 VSS.n628 VSS.n627 68.3621
R4995 VSS.n905 VSS.n454 68.3621
R4996 VSS.n972 VSS.n971 68.3621
R4997 VSS.n1086 VSS.n1021 68.3621
R4998 VSS.n1153 VSS.n1152 68.3621
R4999 VSS.n9548 VSS.n9547 68.2657
R5000 VSS.n9642 VSS.n9641 68.2657
R5001 VSS.n17120 VSS.n17105 63.954
R5002 VSS.n17264 VSS.n17263 63.954
R5003 VSS.n17712 VSS.n17697 63.954
R5004 VSS.n17856 VSS.n17855 63.954
R5005 VSS.n9762 VSS.n9747 63.954
R5006 VSS.n9907 VSS.n9906 63.954
R5007 VSS.n16705 VSS.n16690 63.954
R5008 VSS.n16850 VSS.n16849 63.954
R5009 VSS.n16112 VSS.n16097 63.954
R5010 VSS.n16257 VSS.n16256 63.954
R5011 VSS.n2297 VSS.n2070 63.954
R5012 VSS.n2203 VSS.n2197 63.954
R5013 VSS.n3253 VSS.n3238 63.954
R5014 VSS.n3398 VSS.n3397 63.954
R5015 VSS.n3845 VSS.n3830 63.954
R5016 VSS.n3990 VSS.n3989 63.954
R5017 VSS.n4437 VSS.n4422 63.954
R5018 VSS.n4582 VSS.n4581 63.954
R5019 VSS.n5029 VSS.n5014 63.954
R5020 VSS.n5174 VSS.n5173 63.954
R5021 VSS.n5262 VSS.n2666 63.954
R5022 VSS.n2799 VSS.n2793 63.954
R5023 VSS.n5835 VSS.n5627 63.954
R5024 VSS.n18880 VSS.n18879 63.954
R5025 VSS.n6427 VSS.n6200 63.954
R5026 VSS.n6333 VSS.n6327 63.954
R5027 VSS.n7986 VSS.n7971 63.954
R5028 VSS.n8131 VSS.n8130 63.954
R5029 VSS.n8578 VSS.n8563 63.954
R5030 VSS.n8723 VSS.n8722 63.954
R5031 VSS.n9170 VSS.n9155 63.954
R5032 VSS.n9315 VSS.n9314 63.954
R5033 VSS.n10354 VSS.n10339 63.954
R5034 VSS.n10499 VSS.n10498 63.954
R5035 VSS.n10946 VSS.n10931 63.954
R5036 VSS.n11091 VSS.n11090 63.954
R5037 VSS.n11538 VSS.n11523 63.954
R5038 VSS.n11683 VSS.n11682 63.954
R5039 VSS.n12130 VSS.n12115 63.954
R5040 VSS.n12275 VSS.n12274 63.954
R5041 VSS.n12722 VSS.n12707 63.954
R5042 VSS.n12867 VSS.n12866 63.954
R5043 VSS.n13314 VSS.n13299 63.954
R5044 VSS.n13459 VSS.n13458 63.954
R5045 VSS.n13906 VSS.n13891 63.954
R5046 VSS.n14051 VSS.n14050 63.954
R5047 VSS.n14498 VSS.n14483 63.954
R5048 VSS.n14643 VSS.n14642 63.954
R5049 VSS.n15090 VSS.n15075 63.954
R5050 VSS.n15235 VSS.n15234 63.954
R5051 VSS.n15682 VSS.n15667 63.954
R5052 VSS.n15827 VSS.n15826 63.954
R5053 VSS.n15915 VSS.n6806 63.954
R5054 VSS.n6939 VSS.n6933 63.954
R5055 VSS.n7394 VSS.n7379 63.954
R5056 VSS.n7539 VSS.n7538 63.954
R5057 VSS.n18706 VSS.n18691 63.954
R5058 VSS.n18851 VSS.n18850 63.954
R5059 VSS.n18532 VSS.n18305 63.954
R5060 VSS.n18460 VSS.n18459 63.954
R5061 VSS.n829 VSS.n629 63.954
R5062 VSS.n18872 VSS.n41 63.954
R5063 VSS.n17497 VSS.t615 53.3045
R5064 VSS.n17947 VSS.n1288 53.2877
R5065 VSS.n1421 VSS.n24 53.2877
R5066 VSS.n494 VSS.t235 46.866
R5067 VSS.n1061 VSS.t256 46.866
R5068 VSS.n17424 VSS.t410 46.866
R5069 VSS.n216 VSS.t467 46.866
R5070 VSS.n9474 VSS.t250 46.866
R5071 VSS.n16416 VSS.t529 46.866
R5072 VSS.n1581 VSS.t324 46.866
R5073 VSS.n1766 VSS.t207 46.866
R5074 VSS.n2965 VSS.t282 46.866
R5075 VSS.n3557 VSS.t265 46.866
R5076 VSS.n4149 VSS.t321 46.866
R5077 VSS.n4741 VSS.t192 46.866
R5078 VSS.n2362 VSS.t149 46.866
R5079 VSS.n5323 VSS.t384 46.866
R5080 VSS.n5896 VSS.t56 46.866
R5081 VSS.n7698 VSS.t428 46.866
R5082 VSS.n8290 VSS.t201 46.866
R5083 VSS.n8882 VSS.t109 46.866
R5084 VSS.n10066 VSS.t636 46.866
R5085 VSS.n10658 VSS.t304 46.866
R5086 VSS.n11250 VSS.t535 46.866
R5087 VSS.n11842 VSS.t603 46.866
R5088 VSS.n12434 VSS.t624 46.866
R5089 VSS.n13026 VSS.t194 46.866
R5090 VSS.n13618 VSS.t368 46.866
R5091 VSS.n14210 VSS.t301 46.866
R5092 VSS.n14802 VSS.t404 46.866
R5093 VSS.n15394 VSS.t471 46.866
R5094 VSS.n6502 VSS.t436 46.866
R5095 VSS.n7105 VSS.t503 46.866
R5096 VSS.n196 VSS.t14 46.866
R5097 VSS.n1195 VSS.t585 46.863
R5098 VSS.n16935 VSS.t248 46.863
R5099 VSS.n17349 VSS.t47 46.863
R5100 VSS.n18212 VSS.t70 46.863
R5101 VSS.n9399 VSS.t66 46.863
R5102 VSS.n16341 VSS.t144 46.863
R5103 VSS.n1513 VSS.t456 46.863
R5104 VSS.n1977 VSS.t285 46.863
R5105 VSS.n2890 VSS.t314 46.863
R5106 VSS.n3482 VSS.t295 46.863
R5107 VSS.n4074 VSS.t76 46.863
R5108 VSS.n4666 VSS.t365 46.863
R5109 VSS.n2573 VSS.t550 46.863
R5110 VSS.n5534 VSS.t419 46.863
R5111 VSS.n6107 VSS.t82 46.863
R5112 VSS.n7623 VSS.t73 46.863
R5113 VSS.n8215 VSS.t94 46.863
R5114 VSS.n8807 VSS.t86 46.863
R5115 VSS.n9991 VSS.t101 46.863
R5116 VSS.n10583 VSS.t520 46.863
R5117 VSS.n11175 VSS.t396 46.863
R5118 VSS.n11767 VSS.t245 46.863
R5119 VSS.n12359 VSS.t222 46.863
R5120 VSS.n12951 VSS.t169 46.863
R5121 VSS.n13543 VSS.t44 46.863
R5122 VSS.n14135 VSS.t162 46.863
R5123 VSS.n14727 VSS.t526 46.863
R5124 VSS.n15319 VSS.t180 46.863
R5125 VSS.n6713 VSS.t414 46.863
R5126 VSS.n7030 VSS.t386 46.863
R5127 VSS.n128 VSS.t130 46.863
R5128 VSS.n533 VSS.t127 46.863
R5129 VSS.n1166 VSS.t371 46.8459
R5130 VSS.n16985 VSS.t524 46.8459
R5131 VSS.n17399 VSS.t352 46.8459
R5132 VSS.n18183 VSS.t299 46.8459
R5133 VSS.n9449 VSS.t478 46.8459
R5134 VSS.n16391 VSS.t11 46.8459
R5135 VSS.n1563 VSS.t345 46.8459
R5136 VSS.n1948 VSS.t133 46.8459
R5137 VSS.n2940 VSS.t592 46.8459
R5138 VSS.n3532 VSS.t311 46.8459
R5139 VSS.n4124 VSS.t213 46.8459
R5140 VSS.n4716 VSS.t553 46.8459
R5141 VSS.n2544 VSS.t92 46.8459
R5142 VSS.n5505 VSS.t454 46.8459
R5143 VSS.n6078 VSS.t220 46.8459
R5144 VSS.n7673 VSS.t547 46.8459
R5145 VSS.n8265 VSS.t484 46.8459
R5146 VSS.n8857 VSS.t275 46.8459
R5147 VSS.n10041 VSS.t125 46.8459
R5148 VSS.n10633 VSS.t98 46.8459
R5149 VSS.n11225 VSS.t204 46.8459
R5150 VSS.n11817 VSS.t147 46.8459
R5151 VSS.n12409 VSS.t253 46.8459
R5152 VSS.n13001 VSS.t104 46.8459
R5153 VSS.n13593 VSS.t447 46.8459
R5154 VSS.n14185 VSS.t157 46.8459
R5155 VSS.n14777 VSS.t160 46.8459
R5156 VSS.n15369 VSS.t334 46.8459
R5157 VSS.n6684 VSS.t481 46.8459
R5158 VSS.n7080 VSS.t559 46.8459
R5159 VSS.n178 VSS.t392 46.8459
R5160 VSS.n504 VSS.t574 46.8459
R5161 VSS.n464 VSS.t233 46.8455
R5162 VSS.n1031 VSS.t423 46.8455
R5163 VSS.n17486 VSS.t616 46.8455
R5164 VSS.n278 VSS.t487 46.8455
R5165 VSS.n9536 VSS.t89 46.8455
R5166 VSS.n16467 VSS.t533 46.8455
R5167 VSS.n1632 VSS.t54 46.8455
R5168 VSS.n1828 VSS.t358 46.8455
R5169 VSS.n3027 VSS.t210 46.8455
R5170 VSS.n3619 VSS.t634 46.8455
R5171 VSS.n4211 VSS.t566 46.8455
R5172 VSS.n4803 VSS.t263 46.8455
R5173 VSS.n2424 VSS.t510 46.8455
R5174 VSS.n5385 VSS.t230 46.8455
R5175 VSS.n5958 VSS.t25 46.8455
R5176 VSS.n7760 VSS.t50 46.8455
R5177 VSS.n8352 VSS.t327 46.8455
R5178 VSS.n8944 VSS.t426 46.8455
R5179 VSS.n10128 VSS.t107 46.8455
R5180 VSS.n10720 VSS.t609 46.8455
R5181 VSS.n11312 VSS.t237 46.8455
R5182 VSS.n11904 VSS.t339 46.8455
R5183 VSS.n12496 VSS.t627 46.8455
R5184 VSS.n13088 VSS.t356 46.8455
R5185 VSS.n13680 VSS.t417 46.8455
R5186 VSS.n14272 VSS.t556 46.8455
R5187 VSS.n14864 VSS.t8 46.8455
R5188 VSS.n15456 VSS.t606 46.8455
R5189 VSS.n6564 VSS.t140 46.8455
R5190 VSS.n7156 VSS.t22 46.8455
R5191 VSS.n298 VSS.t390 46.8455
R5192 VSS.n17250 VSS.t174 46.8085
R5193 VSS.n17842 VSS.t569 46.8085
R5194 VSS.n18426 VSS.t350 46.8085
R5195 VSS.n9893 VSS.t450 46.8085
R5196 VSS.n16836 VSS.t63 46.8085
R5197 VSS.n16243 VSS.t513 46.8085
R5198 VSS.n2213 VSS.t474 46.8085
R5199 VSS.n3384 VSS.t576 46.8085
R5200 VSS.n3976 VSS.t135 46.8085
R5201 VSS.n4568 VSS.t270 46.8085
R5202 VSS.n5160 VSS.t400 46.8085
R5203 VSS.n2809 VSS.t506 46.8085
R5204 VSS.n5735 VSS.t18 46.8085
R5205 VSS.n6343 VSS.t32 46.8085
R5206 VSS.n8117 VSS.t362 46.8085
R5207 VSS.n8709 VSS.t495 46.8085
R5208 VSS.n9301 VSS.t407 46.8085
R5209 VSS.n10485 VSS.t379 46.8085
R5210 VSS.n11077 VSS.t165 46.8085
R5211 VSS.n11669 VSS.t59 46.8085
R5212 VSS.n12261 VSS.t260 46.8085
R5213 VSS.n12853 VSS.t442 46.8085
R5214 VSS.n13445 VSS.t4 46.8085
R5215 VSS.n14037 VSS.t461 46.8085
R5216 VSS.n14629 VSS.t40 46.8085
R5217 VSS.n15221 VSS.t153 46.8085
R5218 VSS.n15813 VSS.t375 46.8085
R5219 VSS.n6949 VSS.t114 46.8085
R5220 VSS.n7525 VSS.t438 46.8085
R5221 VSS.n18837 VSS.t183 46.8085
R5222 VSS.n736 VSS.t336 46.8085
R5223 VSS.n1431 VSS.t630 46.8085
R5224 VSS.n16911 VSS.t599 46.808
R5225 VSS.n17325 VSS.t121 46.808
R5226 VSS.n18507 VSS.t287 46.808
R5227 VSS.n9375 VSS.t36 46.808
R5228 VSS.n16317 VSS.t491 46.808
R5229 VSS.n1489 VSS.t562 46.808
R5230 VSS.n2120 VSS.t79 46.808
R5231 VSS.n2866 VSS.t465 46.808
R5232 VSS.n3458 VSS.t612 46.808
R5233 VSS.n4050 VSS.t517 46.808
R5234 VSS.n4642 VSS.t177 46.808
R5235 VSS.n2716 VSS.t215 46.808
R5236 VSS.n5677 VSS.t117 46.808
R5237 VSS.n6250 VSS.t619 46.808
R5238 VSS.n7599 VSS.t240 46.808
R5239 VSS.n8191 VSS.t500 46.808
R5240 VSS.n8783 VSS.t542 46.808
R5241 VSS.n9967 VSS.t277 46.808
R5242 VSS.n10559 VSS.t588 46.808
R5243 VSS.n11151 VSS.t225 46.808
R5244 VSS.n11743 VSS.t307 46.808
R5245 VSS.n12335 VSS.t28 46.808
R5246 VSS.n12927 VSS.t329 46.808
R5247 VSS.n13519 VSS.t538 46.808
R5248 VSS.n14111 VSS.t317 46.808
R5249 VSS.n14703 VSS.t581 46.808
R5250 VSS.n15295 VSS.t595 46.808
R5251 VSS.n6856 VSS.t291 46.808
R5252 VSS.n7006 VSS.t432 46.808
R5253 VSS.n104 VSS.t342 46.808
R5254 VSS.n679 VSS.t188 46.808
R5255 VSS.n1338 VSS.t199 46.808
R5256 VSS.n17995 VSS.n1156 44.8985
R5257 VSS.n17950 VSS.n1287 44.8985
R5258 VSS.n17124 VSS.n17105 44.7679
R5259 VSS.n17263 VSS.n25 44.7679
R5260 VSS.n17716 VSS.n17697 44.7679
R5261 VSS.n17855 VSS.n23 44.7679
R5262 VSS.n9766 VSS.n9747 44.7679
R5263 VSS.n9906 VSS.n32 44.7679
R5264 VSS.n16709 VSS.n16690 44.7679
R5265 VSS.n16849 VSS.n22 44.7679
R5266 VSS.n16116 VSS.n16097 44.7679
R5267 VSS.n16256 VSS.n26 44.7679
R5268 VSS.n2301 VSS.n2070 44.7679
R5269 VSS.n2203 VSS.n21 44.7679
R5270 VSS.n3257 VSS.n3238 44.7679
R5271 VSS.n3397 VSS.n27 44.7679
R5272 VSS.n3849 VSS.n3830 44.7679
R5273 VSS.n3989 VSS.n20 44.7679
R5274 VSS.n4441 VSS.n4422 44.7679
R5275 VSS.n4581 VSS.n28 44.7679
R5276 VSS.n5033 VSS.n5014 44.7679
R5277 VSS.n5173 VSS.n19 44.7679
R5278 VSS.n5266 VSS.n2666 44.7679
R5279 VSS.n2799 VSS.n29 44.7679
R5280 VSS.n5839 VSS.n5627 44.7679
R5281 VSS.n18879 VSS.n18878 44.7679
R5282 VSS.n6431 VSS.n6200 44.7679
R5283 VSS.n6333 VSS.n30 44.7679
R5284 VSS.n7990 VSS.n7971 44.7679
R5285 VSS.n8130 VSS.n18 44.7679
R5286 VSS.n8582 VSS.n8563 44.7679
R5287 VSS.n8722 VSS.n31 44.7679
R5288 VSS.n9174 VSS.n9155 44.7679
R5289 VSS.n9314 VSS.n17 44.7679
R5290 VSS.n10358 VSS.n10339 44.7679
R5291 VSS.n10498 VSS.n16 44.7679
R5292 VSS.n10950 VSS.n10931 44.7679
R5293 VSS.n11090 VSS.n33 44.7679
R5294 VSS.n11542 VSS.n11523 44.7679
R5295 VSS.n11682 VSS.n15 44.7679
R5296 VSS.n12134 VSS.n12115 44.7679
R5297 VSS.n12274 VSS.n34 44.7679
R5298 VSS.n12726 VSS.n12707 44.7679
R5299 VSS.n12866 VSS.n14 44.7679
R5300 VSS.n13318 VSS.n13299 44.7679
R5301 VSS.n13458 VSS.n35 44.7679
R5302 VSS.n13910 VSS.n13891 44.7679
R5303 VSS.n14050 VSS.n13 44.7679
R5304 VSS.n14502 VSS.n14483 44.7679
R5305 VSS.n14642 VSS.n36 44.7679
R5306 VSS.n15094 VSS.n15075 44.7679
R5307 VSS.n15234 VSS.n12 44.7679
R5308 VSS.n15686 VSS.n15667 44.7679
R5309 VSS.n15826 VSS.n37 44.7679
R5310 VSS.n15919 VSS.n6806 44.7679
R5311 VSS.n6939 VSS.n11 44.7679
R5312 VSS.n7398 VSS.n7379 44.7679
R5313 VSS.n7538 VSS.n38 44.7679
R5314 VSS.n18710 VSS.n18691 44.7679
R5315 VSS.n18850 VSS.n39 44.7679
R5316 VSS.n18536 VSS.n18305 44.7679
R5317 VSS.n18459 VSS.n10 44.7679
R5318 VSS.n833 VSS.n629 44.7679
R5319 VSS.n18876 VSS.n41 44.7679
R5320 VSS.n17942 VSS.n17941 38.0628
R5321 VSS.n17875 VSS.n17874 38.0628
R5322 VSS.n10140 VSS.n10138 37.3414
R5323 VSS.n10234 VSS.n6484 37.3414
R5324 VSS.n17003 VSS.n17001 37.2886
R5325 VSS.n17127 VSS.n17104 37.2886
R5326 VSS.n17417 VSS.n17415 37.2886
R5327 VSS.n17719 VSS.n17696 37.2886
R5328 VSS.n18075 VSS.n18073 37.2886
R5329 VSS.n18169 VSS.n208 37.2886
R5330 VSS.n9467 VSS.n9465 37.2886
R5331 VSS.n9769 VSS.n9746 37.2886
R5332 VSS.n16409 VSS.n16407 37.2886
R5333 VSS.n16712 VSS.n16689 37.2886
R5334 VSS.n16484 VSS.n16482 37.2886
R5335 VSS.n16586 VSS.n16585 37.2886
R5336 VSS.n1757 VSS.n1752 37.2886
R5337 VSS.n16119 VSS.n16096 37.2886
R5338 VSS.n1649 VSS.n1647 37.2886
R5339 VSS.n15993 VSS.n1750 37.2886
R5340 VSS.n2349 VSS.n1759 37.2886
R5341 VSS.n2304 VSS.n2069 37.2886
R5342 VSS.n1840 VSS.n1838 37.2886
R5343 VSS.n1934 VSS.n1758 37.2886
R5344 VSS.n2958 VSS.n2956 37.2886
R5345 VSS.n3260 VSS.n3237 37.2886
R5346 VSS.n3039 VSS.n3037 37.2886
R5347 VSS.n3133 VSS.n2350 37.2886
R5348 VSS.n3550 VSS.n3548 37.2886
R5349 VSS.n3852 VSS.n3829 37.2886
R5350 VSS.n3631 VSS.n3629 37.2886
R5351 VSS.n3725 VSS.n2351 37.2886
R5352 VSS.n4142 VSS.n4140 37.2886
R5353 VSS.n4444 VSS.n4421 37.2886
R5354 VSS.n4223 VSS.n4221 37.2886
R5355 VSS.n4317 VSS.n2352 37.2886
R5356 VSS.n4734 VSS.n4732 37.2886
R5357 VSS.n5036 VSS.n5013 37.2886
R5358 VSS.n4815 VSS.n4813 37.2886
R5359 VSS.n4909 VSS.n2353 37.2886
R5360 VSS.n5314 VSS.n2355 37.2886
R5361 VSS.n5269 VSS.n2665 37.2886
R5362 VSS.n2436 VSS.n2434 37.2886
R5363 VSS.n2530 VSS.n2354 37.2886
R5364 VSS.n5887 VSS.n5316 37.2886
R5365 VSS.n5842 VSS.n5626 37.2886
R5366 VSS.n5397 VSS.n5395 37.2886
R5367 VSS.n5491 VSS.n5315 37.2886
R5368 VSS.n6479 VSS.n5889 37.2886
R5369 VSS.n6434 VSS.n6199 37.2886
R5370 VSS.n5970 VSS.n5968 37.2886
R5371 VSS.n6064 VSS.n5888 37.2886
R5372 VSS.n7691 VSS.n7689 37.2886
R5373 VSS.n7993 VSS.n7970 37.2886
R5374 VSS.n7772 VSS.n7770 37.2886
R5375 VSS.n7866 VSS.n6480 37.2886
R5376 VSS.n8283 VSS.n8281 37.2886
R5377 VSS.n8585 VSS.n8562 37.2886
R5378 VSS.n8364 VSS.n8362 37.2886
R5379 VSS.n8458 VSS.n6481 37.2886
R5380 VSS.n8875 VSS.n8873 37.2886
R5381 VSS.n9177 VSS.n9154 37.2886
R5382 VSS.n8956 VSS.n8954 37.2886
R5383 VSS.n9050 VSS.n6482 37.2886
R5384 VSS.n10059 VSS.n10057 37.2886
R5385 VSS.n10361 VSS.n10338 37.2886
R5386 VSS.n10651 VSS.n10649 37.2886
R5387 VSS.n10953 VSS.n10930 37.2886
R5388 VSS.n10732 VSS.n10730 37.2886
R5389 VSS.n10826 VSS.n6485 37.2886
R5390 VSS.n11243 VSS.n11241 37.2886
R5391 VSS.n11545 VSS.n11522 37.2886
R5392 VSS.n11324 VSS.n11322 37.2886
R5393 VSS.n11418 VSS.n6486 37.2886
R5394 VSS.n11835 VSS.n11833 37.2886
R5395 VSS.n12137 VSS.n12114 37.2886
R5396 VSS.n11916 VSS.n11914 37.2886
R5397 VSS.n12010 VSS.n6487 37.2886
R5398 VSS.n12427 VSS.n12425 37.2886
R5399 VSS.n12729 VSS.n12706 37.2886
R5400 VSS.n12508 VSS.n12506 37.2886
R5401 VSS.n12602 VSS.n6488 37.2886
R5402 VSS.n13019 VSS.n13017 37.2886
R5403 VSS.n13321 VSS.n13298 37.2886
R5404 VSS.n13100 VSS.n13098 37.2886
R5405 VSS.n13194 VSS.n6489 37.2886
R5406 VSS.n13611 VSS.n13609 37.2886
R5407 VSS.n13913 VSS.n13890 37.2886
R5408 VSS.n13692 VSS.n13690 37.2886
R5409 VSS.n13786 VSS.n6490 37.2886
R5410 VSS.n14203 VSS.n14201 37.2886
R5411 VSS.n14505 VSS.n14482 37.2886
R5412 VSS.n14284 VSS.n14282 37.2886
R5413 VSS.n14378 VSS.n6491 37.2886
R5414 VSS.n14795 VSS.n14793 37.2886
R5415 VSS.n15097 VSS.n15074 37.2886
R5416 VSS.n14876 VSS.n14874 37.2886
R5417 VSS.n14970 VSS.n6492 37.2886
R5418 VSS.n15387 VSS.n15385 37.2886
R5419 VSS.n15689 VSS.n15666 37.2886
R5420 VSS.n15468 VSS.n15466 37.2886
R5421 VSS.n15562 VSS.n6493 37.2886
R5422 VSS.n15967 VSS.n6495 37.2886
R5423 VSS.n15922 VSS.n6805 37.2886
R5424 VSS.n6576 VSS.n6574 37.2886
R5425 VSS.n6670 VSS.n6494 37.2886
R5426 VSS.n7098 VSS.n7096 37.2886
R5427 VSS.n7401 VSS.n7378 37.2886
R5428 VSS.n7173 VSS.n7171 37.2886
R5429 VSS.n7275 VSS.n7274 37.2886
R5430 VSS.n206 VSS.n201 37.2886
R5431 VSS.n18713 VSS.n18690 37.2886
R5432 VSS.n453 VSS.n288 37.2886
R5433 VSS.n18587 VSS.n199 37.2886
R5434 VSS.n18584 VSS.n209 37.2886
R5435 VSS.n18539 VSS.n18304 37.2886
R5436 VSS.n561 VSS.n560 37.2886
R5437 VSS.n836 VSS.n628 37.2886
R5438 VSS.n1018 VSS.n454 37.2886
R5439 VSS.n973 VSS.n972 37.2886
R5440 VSS.n18044 VSS.n1021 37.2886
R5441 VSS.n17999 VSS.n1153 37.2886
R5442 VSS.n9548 VSS.n9546 37.236
R5443 VSS.n9642 VSS.n6483 37.236
R5444 VSS.n17528 VSS.n17527 36.3441
R5445 VSS.n17559 VSS.n17558 36.3441
R5446 VSS.n17949 VSS.n17948 33.5883
R5447 VSS.n17119 VSS.n17118 31.9772
R5448 VSS.n17262 VSS.n17261 31.9772
R5449 VSS.n17711 VSS.n17710 31.9772
R5450 VSS.n17854 VSS.n17853 31.9772
R5451 VSS.n9761 VSS.n9760 31.9772
R5452 VSS.n9905 VSS.n9904 31.9772
R5453 VSS.n16704 VSS.n16703 31.9772
R5454 VSS.n16848 VSS.n16847 31.9772
R5455 VSS.n16111 VSS.n16110 31.9772
R5456 VSS.n16255 VSS.n16254 31.9772
R5457 VSS.n2296 VSS.n2295 31.9772
R5458 VSS.n2229 VSS.n2228 31.9772
R5459 VSS.n3252 VSS.n3251 31.9772
R5460 VSS.n3396 VSS.n3395 31.9772
R5461 VSS.n3844 VSS.n3843 31.9772
R5462 VSS.n3988 VSS.n3987 31.9772
R5463 VSS.n4436 VSS.n4435 31.9772
R5464 VSS.n4580 VSS.n4579 31.9772
R5465 VSS.n5028 VSS.n5027 31.9772
R5466 VSS.n5172 VSS.n5171 31.9772
R5467 VSS.n5261 VSS.n5260 31.9772
R5468 VSS.n5194 VSS.n5193 31.9772
R5469 VSS.n5834 VSS.n5833 31.9772
R5470 VSS.n5767 VSS.n9 31.9772
R5471 VSS.n6426 VSS.n6425 31.9772
R5472 VSS.n6359 VSS.n6358 31.9772
R5473 VSS.n7985 VSS.n7984 31.9772
R5474 VSS.n8129 VSS.n8128 31.9772
R5475 VSS.n8577 VSS.n8576 31.9772
R5476 VSS.n8721 VSS.n8720 31.9772
R5477 VSS.n9169 VSS.n9168 31.9772
R5478 VSS.n9313 VSS.n9312 31.9772
R5479 VSS.n10353 VSS.n10352 31.9772
R5480 VSS.n10497 VSS.n10496 31.9772
R5481 VSS.n10945 VSS.n10944 31.9772
R5482 VSS.n11089 VSS.n11088 31.9772
R5483 VSS.n11537 VSS.n11536 31.9772
R5484 VSS.n11681 VSS.n11680 31.9772
R5485 VSS.n12129 VSS.n12128 31.9772
R5486 VSS.n12273 VSS.n12272 31.9772
R5487 VSS.n12721 VSS.n12720 31.9772
R5488 VSS.n12865 VSS.n12864 31.9772
R5489 VSS.n13313 VSS.n13312 31.9772
R5490 VSS.n13457 VSS.n13456 31.9772
R5491 VSS.n13905 VSS.n13904 31.9772
R5492 VSS.n14049 VSS.n14048 31.9772
R5493 VSS.n14497 VSS.n14496 31.9772
R5494 VSS.n14641 VSS.n14640 31.9772
R5495 VSS.n15089 VSS.n15088 31.9772
R5496 VSS.n15233 VSS.n15232 31.9772
R5497 VSS.n15681 VSS.n15680 31.9772
R5498 VSS.n15825 VSS.n15824 31.9772
R5499 VSS.n15914 VSS.n15913 31.9772
R5500 VSS.n15847 VSS.n15846 31.9772
R5501 VSS.n7393 VSS.n7392 31.9772
R5502 VSS.n7537 VSS.n7536 31.9772
R5503 VSS.n18705 VSS.n18704 31.9772
R5504 VSS.n18849 VSS.n18848 31.9772
R5505 VSS.n18531 VSS.n18530 31.9772
R5506 VSS.n18458 VSS.n18457 31.9772
R5507 VSS.n828 VSS.n827 31.9772
R5508 VSS.n18871 VSS.n18870 31.9772
R5509 VSS.n17525 VSS.n17524 31.4983
R5510 VSS.n17561 VSS.n17560 31.4983
R5511 VSS.n1245 VSS.n1217 29.9325
R5512 VSS.t584 VSS.n1199 29.9325
R5513 VSS.n18877 VSS.t12 27.9932
R5514 VSS.n15980 VSS.n15979 27.5867
R5515 VSS.n17498 VSS.n17497 26.6525
R5516 VSS.n17592 VSS.n17591 26.6525
R5517 VSS.n10166 VSS.n10123 24.8944
R5518 VSS.n17029 VSS.n17028 24.8593
R5519 VSS.t247 VSS.n16938 24.8593
R5520 VSS.n17621 VSS.n17620 24.8593
R5521 VSS.t46 VSS.n17352 24.8593
R5522 VSS.n18101 VSS.n273 24.8593
R5523 VSS.n9671 VSS.n9670 24.8593
R5524 VSS.t65 VSS.n9402 24.8593
R5525 VSS.n16614 VSS.n16613 24.8593
R5526 VSS.t143 VSS.n16344 24.8593
R5527 VSS.n16509 VSS.n16508 24.8593
R5528 VSS.n16021 VSS.n16020 24.8593
R5529 VSS.t455 VSS.n1516 24.8593
R5530 VSS.n1674 VSS.n1673 24.8593
R5531 VSS.n2027 VSS.n1999 24.8593
R5532 VSS.t284 VSS.n1981 24.8593
R5533 VSS.n1866 VSS.n1823 24.8593
R5534 VSS.n3162 VSS.n3161 24.8593
R5535 VSS.t313 VSS.n2893 24.8593
R5536 VSS.n3065 VSS.n3022 24.8593
R5537 VSS.n3754 VSS.n3753 24.8593
R5538 VSS.t294 VSS.n3485 24.8593
R5539 VSS.n3657 VSS.n3614 24.8593
R5540 VSS.n4346 VSS.n4345 24.8593
R5541 VSS.t75 VSS.n4077 24.8593
R5542 VSS.n4249 VSS.n4206 24.8593
R5543 VSS.n4938 VSS.n4937 24.8593
R5544 VSS.t364 VSS.n4669 24.8593
R5545 VSS.n4841 VSS.n4798 24.8593
R5546 VSS.n2623 VSS.n2595 24.8593
R5547 VSS.t549 VSS.n2577 24.8593
R5548 VSS.n2462 VSS.n2419 24.8593
R5549 VSS.n5584 VSS.n5556 24.8593
R5550 VSS.t418 VSS.n5538 24.8593
R5551 VSS.n5423 VSS.n5380 24.8593
R5552 VSS.n6157 VSS.n6129 24.8593
R5553 VSS.t81 VSS.n6111 24.8593
R5554 VSS.n5996 VSS.n5953 24.8593
R5555 VSS.n7895 VSS.n7894 24.8593
R5556 VSS.t72 VSS.n7626 24.8593
R5557 VSS.n7798 VSS.n7755 24.8593
R5558 VSS.n8487 VSS.n8486 24.8593
R5559 VSS.t93 VSS.n8218 24.8593
R5560 VSS.n8390 VSS.n8347 24.8593
R5561 VSS.n9079 VSS.n9078 24.8593
R5562 VSS.t85 VSS.n8810 24.8593
R5563 VSS.n8982 VSS.n8939 24.8593
R5564 VSS.n10263 VSS.n10262 24.8593
R5565 VSS.t100 VSS.n9994 24.8593
R5566 VSS.n10855 VSS.n10854 24.8593
R5567 VSS.t519 VSS.n10586 24.8593
R5568 VSS.n10758 VSS.n10715 24.8593
R5569 VSS.n11447 VSS.n11446 24.8593
R5570 VSS.t395 VSS.n11178 24.8593
R5571 VSS.n11350 VSS.n11307 24.8593
R5572 VSS.n12039 VSS.n12038 24.8593
R5573 VSS.t244 VSS.n11770 24.8593
R5574 VSS.n11942 VSS.n11899 24.8593
R5575 VSS.n12631 VSS.n12630 24.8593
R5576 VSS.t221 VSS.n12362 24.8593
R5577 VSS.n12534 VSS.n12491 24.8593
R5578 VSS.n13223 VSS.n13222 24.8593
R5579 VSS.t168 VSS.n12954 24.8593
R5580 VSS.n13126 VSS.n13083 24.8593
R5581 VSS.n13815 VSS.n13814 24.8593
R5582 VSS.t43 VSS.n13546 24.8593
R5583 VSS.n13718 VSS.n13675 24.8593
R5584 VSS.n14407 VSS.n14406 24.8593
R5585 VSS.t161 VSS.n14138 24.8593
R5586 VSS.n14310 VSS.n14267 24.8593
R5587 VSS.n14999 VSS.n14998 24.8593
R5588 VSS.t525 VSS.n14730 24.8593
R5589 VSS.n14902 VSS.n14859 24.8593
R5590 VSS.n15591 VSS.n15590 24.8593
R5591 VSS.t179 VSS.n15322 24.8593
R5592 VSS.n15494 VSS.n15451 24.8593
R5593 VSS.n6763 VSS.n6735 24.8593
R5594 VSS.t413 VSS.n6717 24.8593
R5595 VSS.n6602 VSS.n6559 24.8593
R5596 VSS.n7303 VSS.n7302 24.8593
R5597 VSS.t385 VSS.n7033 24.8593
R5598 VSS.n7198 VSS.n7197 24.8593
R5599 VSS.n18615 VSS.n18614 24.8593
R5600 VSS.t129 VSS.n131 24.8593
R5601 VSS.n361 VSS.n360 24.8593
R5602 VSS.n18262 VSS.n18234 24.8593
R5603 VSS.t69 VSS.n18216 24.8593
R5604 VSS.n586 VSS.n555 24.8593
R5605 VSS.t126 VSS.n537 24.8593
R5606 VSS.n929 VSS.n903 24.8593
R5607 VSS.n1110 VSS.n1084 24.8593
R5608 VSS.n9574 VSS.n9531 24.8242
R5609 VSS.n16914 VSS.n16894 24.6255
R5610 VSS.n17218 VSS.n16892 24.6255
R5611 VSS.n17328 VSS.n17308 24.6255
R5612 VSS.n17810 VSS.n17306 24.6255
R5613 VSS.n18381 VSS.n18359 24.6255
R5614 VSS.n18493 VSS.n18360 24.6255
R5615 VSS.n9378 VSS.n9358 24.6255
R5616 VSS.n9860 VSS.n9356 24.6255
R5617 VSS.n16320 VSS.n16300 24.6255
R5618 VSS.n16803 VSS.n16298 24.6255
R5619 VSS.n1492 VSS.n1472 24.6255
R5620 VSS.n16210 VSS.n1470 24.6255
R5621 VSS.n2266 VSS.n2122 24.6255
R5622 VSS.n2187 VSS.n2124 24.6255
R5623 VSS.n2869 VSS.n2849 24.6255
R5624 VSS.n3351 VSS.n2847 24.6255
R5625 VSS.n3461 VSS.n3441 24.6255
R5626 VSS.n3943 VSS.n3439 24.6255
R5627 VSS.n4053 VSS.n4033 24.6255
R5628 VSS.n4535 VSS.n4031 24.6255
R5629 VSS.n4645 VSS.n4625 24.6255
R5630 VSS.n5127 VSS.n4623 24.6255
R5631 VSS.n5231 VSS.n2718 24.6255
R5632 VSS.n2783 VSS.n2720 24.6255
R5633 VSS.n5804 VSS.n5679 24.6255
R5634 VSS.n5757 VSS.n5681 24.6255
R5635 VSS.n6396 VSS.n6252 24.6255
R5636 VSS.n6317 VSS.n6254 24.6255
R5637 VSS.n7602 VSS.n7582 24.6255
R5638 VSS.n8084 VSS.n7580 24.6255
R5639 VSS.n8194 VSS.n8174 24.6255
R5640 VSS.n8676 VSS.n8172 24.6255
R5641 VSS.n8786 VSS.n8766 24.6255
R5642 VSS.n9268 VSS.n8764 24.6255
R5643 VSS.n9970 VSS.n9950 24.6255
R5644 VSS.n10452 VSS.n9948 24.6255
R5645 VSS.n10562 VSS.n10542 24.6255
R5646 VSS.n11044 VSS.n10540 24.6255
R5647 VSS.n11154 VSS.n11134 24.6255
R5648 VSS.n11636 VSS.n11132 24.6255
R5649 VSS.n11746 VSS.n11726 24.6255
R5650 VSS.n12228 VSS.n11724 24.6255
R5651 VSS.n12338 VSS.n12318 24.6255
R5652 VSS.n12820 VSS.n12316 24.6255
R5653 VSS.n12930 VSS.n12910 24.6255
R5654 VSS.n13412 VSS.n12908 24.6255
R5655 VSS.n13522 VSS.n13502 24.6255
R5656 VSS.n14004 VSS.n13500 24.6255
R5657 VSS.n14114 VSS.n14094 24.6255
R5658 VSS.n14596 VSS.n14092 24.6255
R5659 VSS.n14706 VSS.n14686 24.6255
R5660 VSS.n15188 VSS.n14684 24.6255
R5661 VSS.n15298 VSS.n15278 24.6255
R5662 VSS.n15780 VSS.n15276 24.6255
R5663 VSS.n15884 VSS.n6858 24.6255
R5664 VSS.n6923 VSS.n6860 24.6255
R5665 VSS.n7009 VSS.n6989 24.6255
R5666 VSS.n7492 VSS.n6987 24.6255
R5667 VSS.n107 VSS.n87 24.6255
R5668 VSS.n18804 VSS.n85 24.6255
R5669 VSS.n798 VSS.n681 24.6255
R5670 VSS.n756 VSS.n683 24.6255
R5671 VSS.n17912 VSS.n1340 24.6255
R5672 VSS.n1405 VSS.n1342 24.6255
R5673 VSS.n17927 VSS.n17926 22.8379
R5674 VSS.n1414 VSS.t629 22.8379
R5675 VSS.n17163 VSS.n16913 21.5474
R5676 VSS.n17235 VSS.n16880 21.5474
R5677 VSS.n17755 VSS.n17327 21.5474
R5678 VSS.n17827 VSS.n17294 21.5474
R5679 VSS.n18372 VSS.n18362 21.5474
R5680 VSS.n18449 VSS.n18440 21.5474
R5681 VSS.n9805 VSS.n9377 21.5474
R5682 VSS.n9877 VSS.n9344 21.5474
R5683 VSS.n16748 VSS.n16319 21.5474
R5684 VSS.n16820 VSS.n16286 21.5474
R5685 VSS.n16155 VSS.n1491 21.5474
R5686 VSS.n16227 VSS.n1458 21.5474
R5687 VSS.n2278 VSS.n2104 21.5474
R5688 VSS.n2195 VSS.n2191 21.5474
R5689 VSS.n3296 VSS.n2868 21.5474
R5690 VSS.n3368 VSS.n2835 21.5474
R5691 VSS.n3888 VSS.n3460 21.5474
R5692 VSS.n3960 VSS.n3427 21.5474
R5693 VSS.n4480 VSS.n4052 21.5474
R5694 VSS.n4552 VSS.n4019 21.5474
R5695 VSS.n5072 VSS.n4644 21.5474
R5696 VSS.n5144 VSS.n4611 21.5474
R5697 VSS.n5243 VSS.n2700 21.5474
R5698 VSS.n2791 VSS.n2787 21.5474
R5699 VSS.n5816 VSS.n5661 21.5474
R5700 VSS.n5765 VSS.n5761 21.5474
R5701 VSS.n6408 VSS.n6234 21.5474
R5702 VSS.n6325 VSS.n6321 21.5474
R5703 VSS.n8029 VSS.n7601 21.5474
R5704 VSS.n8101 VSS.n7568 21.5474
R5705 VSS.n8621 VSS.n8193 21.5474
R5706 VSS.n8693 VSS.n8160 21.5474
R5707 VSS.n9213 VSS.n8785 21.5474
R5708 VSS.n9285 VSS.n8752 21.5474
R5709 VSS.n10397 VSS.n9969 21.5474
R5710 VSS.n10469 VSS.n9936 21.5474
R5711 VSS.n10989 VSS.n10561 21.5474
R5712 VSS.n11061 VSS.n10528 21.5474
R5713 VSS.n11581 VSS.n11153 21.5474
R5714 VSS.n11653 VSS.n11120 21.5474
R5715 VSS.n12173 VSS.n11745 21.5474
R5716 VSS.n12245 VSS.n11712 21.5474
R5717 VSS.n12765 VSS.n12337 21.5474
R5718 VSS.n12837 VSS.n12304 21.5474
R5719 VSS.n13357 VSS.n12929 21.5474
R5720 VSS.n13429 VSS.n12896 21.5474
R5721 VSS.n13949 VSS.n13521 21.5474
R5722 VSS.n14021 VSS.n13488 21.5474
R5723 VSS.n14541 VSS.n14113 21.5474
R5724 VSS.n14613 VSS.n14080 21.5474
R5725 VSS.n15133 VSS.n14705 21.5474
R5726 VSS.n15205 VSS.n14672 21.5474
R5727 VSS.n15725 VSS.n15297 21.5474
R5728 VSS.n15797 VSS.n15264 21.5474
R5729 VSS.n15896 VSS.n6840 21.5474
R5730 VSS.n6931 VSS.n6927 21.5474
R5731 VSS.n7437 VSS.n7008 21.5474
R5732 VSS.n7509 VSS.n6975 21.5474
R5733 VSS.n18749 VSS.n106 21.5474
R5734 VSS.n18821 VSS.n73 21.5474
R5735 VSS.n810 VSS.n663 21.5474
R5736 VSS.n758 VSS.n744 21.5474
R5737 VSS.n17924 VSS.n1322 21.5474
R5738 VSS.n1413 VSS.n1409 21.5474
R5739 VSS.n1252 VSS.n1213 21.1076
R5740 VSS.n1256 VSS.n1209 21.1076
R5741 VSS.n17526 VSS.n17480 21.1076
R5742 VSS.n17557 VSS.n17450 21.1076
R5743 VSS.n1117 VSS.n1080 21.1076
R5744 VSS.n1121 VSS.n1075 21.1076
R5745 VSS.n936 VSS.n899 21.1076
R5746 VSS.n940 VSS.n894 21.1076
R5747 VSS.n17049 VSS.n16972 21.1076
R5748 VSS.n16973 VSS.n16954 21.1076
R5749 VSS.n17641 VSS.n17386 21.1076
R5750 VSS.n17387 VSS.n17368 21.1076
R5751 VSS.n18269 VSS.n18230 21.1076
R5752 VSS.n18273 VSS.n18226 21.1076
R5753 VSS.n18103 VSS.n272 21.1076
R5754 VSS.n18134 VSS.n242 21.1076
R5755 VSS.n9576 VSS.n9530 21.1076
R5756 VSS.n9607 VSS.n9500 21.1076
R5757 VSS.n9691 VSS.n9436 21.1076
R5758 VSS.n9437 VSS.n9418 21.1076
R5759 VSS.n16529 VSS.n16455 21.1076
R5760 VSS.n16456 VSS.n16435 21.1076
R5761 VSS.n16634 VSS.n16378 21.1076
R5762 VSS.n16379 VSS.n16360 21.1076
R5763 VSS.n1694 VSS.n1620 21.1076
R5764 VSS.n1621 VSS.n1600 21.1076
R5765 VSS.n16041 VSS.n1550 21.1076
R5766 VSS.n1551 VSS.n1532 21.1076
R5767 VSS.n1868 VSS.n1822 21.1076
R5768 VSS.n1899 VSS.n1792 21.1076
R5769 VSS.n2034 VSS.n1995 21.1076
R5770 VSS.n2038 VSS.n1991 21.1076
R5771 VSS.n3067 VSS.n3021 21.1076
R5772 VSS.n3098 VSS.n2991 21.1076
R5773 VSS.n3182 VSS.n2927 21.1076
R5774 VSS.n2928 VSS.n2909 21.1076
R5775 VSS.n3659 VSS.n3613 21.1076
R5776 VSS.n3690 VSS.n3583 21.1076
R5777 VSS.n3774 VSS.n3519 21.1076
R5778 VSS.n3520 VSS.n3501 21.1076
R5779 VSS.n4251 VSS.n4205 21.1076
R5780 VSS.n4282 VSS.n4175 21.1076
R5781 VSS.n4366 VSS.n4111 21.1076
R5782 VSS.n4112 VSS.n4093 21.1076
R5783 VSS.n4843 VSS.n4797 21.1076
R5784 VSS.n4874 VSS.n4767 21.1076
R5785 VSS.n4958 VSS.n4703 21.1076
R5786 VSS.n4704 VSS.n4685 21.1076
R5787 VSS.n2464 VSS.n2418 21.1076
R5788 VSS.n2495 VSS.n2388 21.1076
R5789 VSS.n2630 VSS.n2591 21.1076
R5790 VSS.n2634 VSS.n2587 21.1076
R5791 VSS.n5425 VSS.n5379 21.1076
R5792 VSS.n5456 VSS.n5349 21.1076
R5793 VSS.n5591 VSS.n5552 21.1076
R5794 VSS.n5595 VSS.n5548 21.1076
R5795 VSS.n5998 VSS.n5952 21.1076
R5796 VSS.n6029 VSS.n5922 21.1076
R5797 VSS.n6164 VSS.n6125 21.1076
R5798 VSS.n6168 VSS.n6121 21.1076
R5799 VSS.n7800 VSS.n7754 21.1076
R5800 VSS.n7831 VSS.n7724 21.1076
R5801 VSS.n7915 VSS.n7660 21.1076
R5802 VSS.n7661 VSS.n7642 21.1076
R5803 VSS.n8392 VSS.n8346 21.1076
R5804 VSS.n8423 VSS.n8316 21.1076
R5805 VSS.n8507 VSS.n8252 21.1076
R5806 VSS.n8253 VSS.n8234 21.1076
R5807 VSS.n8984 VSS.n8938 21.1076
R5808 VSS.n9015 VSS.n8908 21.1076
R5809 VSS.n9099 VSS.n8844 21.1076
R5810 VSS.n8845 VSS.n8826 21.1076
R5811 VSS.n10168 VSS.n10122 21.1076
R5812 VSS.n10199 VSS.n10092 21.1076
R5813 VSS.n10283 VSS.n10028 21.1076
R5814 VSS.n10029 VSS.n10010 21.1076
R5815 VSS.n10760 VSS.n10714 21.1076
R5816 VSS.n10791 VSS.n10684 21.1076
R5817 VSS.n10875 VSS.n10620 21.1076
R5818 VSS.n10621 VSS.n10602 21.1076
R5819 VSS.n11352 VSS.n11306 21.1076
R5820 VSS.n11383 VSS.n11276 21.1076
R5821 VSS.n11467 VSS.n11212 21.1076
R5822 VSS.n11213 VSS.n11194 21.1076
R5823 VSS.n11944 VSS.n11898 21.1076
R5824 VSS.n11975 VSS.n11868 21.1076
R5825 VSS.n12059 VSS.n11804 21.1076
R5826 VSS.n11805 VSS.n11786 21.1076
R5827 VSS.n12536 VSS.n12490 21.1076
R5828 VSS.n12567 VSS.n12460 21.1076
R5829 VSS.n12651 VSS.n12396 21.1076
R5830 VSS.n12397 VSS.n12378 21.1076
R5831 VSS.n13128 VSS.n13082 21.1076
R5832 VSS.n13159 VSS.n13052 21.1076
R5833 VSS.n13243 VSS.n12988 21.1076
R5834 VSS.n12989 VSS.n12970 21.1076
R5835 VSS.n13720 VSS.n13674 21.1076
R5836 VSS.n13751 VSS.n13644 21.1076
R5837 VSS.n13835 VSS.n13580 21.1076
R5838 VSS.n13581 VSS.n13562 21.1076
R5839 VSS.n14312 VSS.n14266 21.1076
R5840 VSS.n14343 VSS.n14236 21.1076
R5841 VSS.n14427 VSS.n14172 21.1076
R5842 VSS.n14173 VSS.n14154 21.1076
R5843 VSS.n14904 VSS.n14858 21.1076
R5844 VSS.n14935 VSS.n14828 21.1076
R5845 VSS.n15019 VSS.n14764 21.1076
R5846 VSS.n14765 VSS.n14746 21.1076
R5847 VSS.n15496 VSS.n15450 21.1076
R5848 VSS.n15527 VSS.n15420 21.1076
R5849 VSS.n15611 VSS.n15356 21.1076
R5850 VSS.n15357 VSS.n15338 21.1076
R5851 VSS.n6604 VSS.n6558 21.1076
R5852 VSS.n6635 VSS.n6528 21.1076
R5853 VSS.n6770 VSS.n6731 21.1076
R5854 VSS.n6774 VSS.n6727 21.1076
R5855 VSS.n7218 VSS.n7144 21.1076
R5856 VSS.n7145 VSS.n7124 21.1076
R5857 VSS.n7323 VSS.n7067 21.1076
R5858 VSS.n7068 VSS.n7049 21.1076
R5859 VSS.n376 VSS.n339 21.1076
R5860 VSS.n381 VSS.n335 21.1076
R5861 VSS.n18635 VSS.n165 21.1076
R5862 VSS.n166 VSS.n147 21.1076
R5863 VSS.n593 VSS.n551 21.1076
R5864 VSS.n597 VSS.n547 21.1076
R5865 VSS.n17164 VSS.n16915 19.1865
R5866 VSS.n17237 VSS.t173 19.1865
R5867 VSS.n17756 VSS.n17329 19.1865
R5868 VSS.n17829 VSS.t568 19.1865
R5869 VSS.n9806 VSS.n9379 19.1865
R5870 VSS.n9879 VSS.t449 19.1865
R5871 VSS.n16749 VSS.n16321 19.1865
R5872 VSS.n16822 VSS.t62 19.1865
R5873 VSS.n16156 VSS.n1493 19.1865
R5874 VSS.n16229 VSS.t512 19.1865
R5875 VSS.n2281 VSS.n2280 19.1865
R5876 VSS.n2196 VSS.t473 19.1865
R5877 VSS.n3297 VSS.n2870 19.1865
R5878 VSS.n3370 VSS.t575 19.1865
R5879 VSS.n3889 VSS.n3462 19.1865
R5880 VSS.n3962 VSS.t134 19.1865
R5881 VSS.n4481 VSS.n4054 19.1865
R5882 VSS.n4554 VSS.t269 19.1865
R5883 VSS.n5073 VSS.n4646 19.1865
R5884 VSS.n5146 VSS.t399 19.1865
R5885 VSS.n5246 VSS.n5245 19.1865
R5886 VSS.n2792 VSS.t505 19.1865
R5887 VSS.n5819 VSS.n5818 19.1865
R5888 VSS.n5766 VSS.t17 19.1865
R5889 VSS.n6411 VSS.n6410 19.1865
R5890 VSS.n6326 VSS.t31 19.1865
R5891 VSS.n8030 VSS.n7603 19.1865
R5892 VSS.n8103 VSS.t361 19.1865
R5893 VSS.n8622 VSS.n8195 19.1865
R5894 VSS.n8695 VSS.t494 19.1865
R5895 VSS.n9214 VSS.n8787 19.1865
R5896 VSS.n9287 VSS.t406 19.1865
R5897 VSS.n10398 VSS.n9971 19.1865
R5898 VSS.n10471 VSS.t378 19.1865
R5899 VSS.n10990 VSS.n10563 19.1865
R5900 VSS.n11063 VSS.t164 19.1865
R5901 VSS.n11582 VSS.n11155 19.1865
R5902 VSS.n11655 VSS.t58 19.1865
R5903 VSS.n12174 VSS.n11747 19.1865
R5904 VSS.n12247 VSS.t259 19.1865
R5905 VSS.n12766 VSS.n12339 19.1865
R5906 VSS.n12839 VSS.t441 19.1865
R5907 VSS.n13358 VSS.n12931 19.1865
R5908 VSS.n13431 VSS.t3 19.1865
R5909 VSS.n13950 VSS.n13523 19.1865
R5910 VSS.n14023 VSS.t460 19.1865
R5911 VSS.n14542 VSS.n14115 19.1865
R5912 VSS.n14615 VSS.t39 19.1865
R5913 VSS.n15134 VSS.n14707 19.1865
R5914 VSS.n15207 VSS.t152 19.1865
R5915 VSS.n15726 VSS.n15299 19.1865
R5916 VSS.n15799 VSS.t374 19.1865
R5917 VSS.n15899 VSS.n15898 19.1865
R5918 VSS.n6932 VSS.t113 19.1865
R5919 VSS.n7438 VSS.n7010 19.1865
R5920 VSS.n7511 VSS.t437 19.1865
R5921 VSS.n18750 VSS.n108 19.1865
R5922 VSS.n18823 VSS.t182 19.1865
R5923 VSS.n18370 VSS.n18369 19.1865
R5924 VSS.n18451 VSS.t349 19.1865
R5925 VSS.n813 VSS.n812 19.1865
R5926 VSS.n760 VSS.t335 19.1865
R5927 VSS.n10232 VSS.t635 18.6709
R5928 VSS.n18167 VSS.t466 18.6446
R5929 VSS.t528 VSS.n16419 18.6446
R5930 VSS.t323 VSS.n1584 18.6446
R5931 VSS.n1932 VSS.t206 18.6446
R5932 VSS.n3131 VSS.t281 18.6446
R5933 VSS.n3723 VSS.t264 18.6446
R5934 VSS.n4315 VSS.t320 18.6446
R5935 VSS.n4907 VSS.t191 18.6446
R5936 VSS.n2528 VSS.t148 18.6446
R5937 VSS.n5489 VSS.t383 18.6446
R5938 VSS.n6062 VSS.t55 18.6446
R5939 VSS.n7864 VSS.t427 18.6446
R5940 VSS.n8456 VSS.t200 18.6446
R5941 VSS.n9048 VSS.t108 18.6446
R5942 VSS.n10824 VSS.t303 18.6446
R5943 VSS.n11416 VSS.t534 18.6446
R5944 VSS.n12008 VSS.t602 18.6446
R5945 VSS.n12600 VSS.t623 18.6446
R5946 VSS.n13192 VSS.t193 18.6446
R5947 VSS.n13784 VSS.t367 18.6446
R5948 VSS.n14376 VSS.t300 18.6446
R5949 VSS.n14968 VSS.t403 18.6446
R5950 VSS.n15560 VSS.t470 18.6446
R5951 VSS.n6668 VSS.t435 18.6446
R5952 VSS.t502 VSS.n7108 18.6446
R5953 VSS.n400 VSS.t13 18.6446
R5954 VSS.t234 VSS.n884 18.6446
R5955 VSS.t255 VSS.n1065 18.6446
R5956 VSS.n9640 VSS.t249 18.6183
R5957 VSS.n17117 VSS.n17113 18.4693
R5958 VSS.n17260 VSS.n16869 18.4693
R5959 VSS.n17709 VSS.n17705 18.4693
R5960 VSS.n17852 VSS.n17283 18.4693
R5961 VSS.n18529 VSS.n18311 18.4693
R5962 VSS.n18456 VSS.n18453 18.4693
R5963 VSS.n9759 VSS.n9755 18.4693
R5964 VSS.n9903 VSS.n9334 18.4693
R5965 VSS.n16702 VSS.n16698 18.4693
R5966 VSS.n16846 VSS.n16276 18.4693
R5967 VSS.n16109 VSS.n16105 18.4693
R5968 VSS.n16253 VSS.n1448 18.4693
R5969 VSS.n2294 VSS.n2076 18.4693
R5970 VSS.n2231 VSS.n2176 18.4693
R5971 VSS.n3250 VSS.n3246 18.4693
R5972 VSS.n3394 VSS.n2825 18.4693
R5973 VSS.n3842 VSS.n3838 18.4693
R5974 VSS.n3986 VSS.n3417 18.4693
R5975 VSS.n4434 VSS.n4430 18.4693
R5976 VSS.n4578 VSS.n4009 18.4693
R5977 VSS.n5026 VSS.n5022 18.4693
R5978 VSS.n5170 VSS.n4601 18.4693
R5979 VSS.n5259 VSS.n2672 18.4693
R5980 VSS.n5196 VSS.n2772 18.4693
R5981 VSS.n5832 VSS.n5633 18.4693
R5982 VSS.n5769 VSS.n5746 18.4693
R5983 VSS.n6424 VSS.n6206 18.4693
R5984 VSS.n6361 VSS.n6306 18.4693
R5985 VSS.n7983 VSS.n7979 18.4693
R5986 VSS.n8127 VSS.n7558 18.4693
R5987 VSS.n8575 VSS.n8571 18.4693
R5988 VSS.n8719 VSS.n8150 18.4693
R5989 VSS.n9167 VSS.n9163 18.4693
R5990 VSS.n9311 VSS.n8742 18.4693
R5991 VSS.n10351 VSS.n10347 18.4693
R5992 VSS.n10495 VSS.n9926 18.4693
R5993 VSS.n10943 VSS.n10939 18.4693
R5994 VSS.n11087 VSS.n10518 18.4693
R5995 VSS.n11535 VSS.n11531 18.4693
R5996 VSS.n11679 VSS.n11110 18.4693
R5997 VSS.n12127 VSS.n12123 18.4693
R5998 VSS.n12271 VSS.n11702 18.4693
R5999 VSS.n12719 VSS.n12715 18.4693
R6000 VSS.n12863 VSS.n12294 18.4693
R6001 VSS.n13311 VSS.n13307 18.4693
R6002 VSS.n13455 VSS.n12886 18.4693
R6003 VSS.n13903 VSS.n13899 18.4693
R6004 VSS.n14047 VSS.n13478 18.4693
R6005 VSS.n14495 VSS.n14491 18.4693
R6006 VSS.n14639 VSS.n14070 18.4693
R6007 VSS.n15087 VSS.n15083 18.4693
R6008 VSS.n15231 VSS.n14662 18.4693
R6009 VSS.n15679 VSS.n15675 18.4693
R6010 VSS.n15823 VSS.n15254 18.4693
R6011 VSS.n15912 VSS.n6812 18.4693
R6012 VSS.n15849 VSS.n6912 18.4693
R6013 VSS.n7391 VSS.n7387 18.4693
R6014 VSS.n7535 VSS.n6965 18.4693
R6015 VSS.n18703 VSS.n18699 18.4693
R6016 VSS.n18847 VSS.n63 18.4693
R6017 VSS.n826 VSS.n635 18.4693
R6018 VSS.n18869 VSS.n47 18.4693
R6019 VSS.n17940 VSS.n1294 18.4693
R6020 VSS.n17877 VSS.n1394 18.4693
R6021 VSS.n1244 VSS.n1216 18.2934
R6022 VSS.n1272 VSS.n1207 18.2934
R6023 VSS.n17523 VSS.n17479 18.2934
R6024 VSS.n17457 VSS.n17427 18.2934
R6025 VSS.n1109 VSS.n1083 18.2934
R6026 VSS.n1138 VSS.n1073 18.2934
R6027 VSS.n928 VSS.n902 18.2934
R6028 VSS.n957 VSS.n892 18.2934
R6029 VSS.n17031 VSS.n16988 18.2934
R6030 VSS.n17083 VSS.n16952 18.2934
R6031 VSS.n17623 VSS.n17402 18.2934
R6032 VSS.n17675 VSS.n17366 18.2934
R6033 VSS.n18261 VSS.n18233 18.2934
R6034 VSS.n18289 VSS.n18224 18.2934
R6035 VSS.n18100 VSS.n271 18.2934
R6036 VSS.n249 VSS.n219 18.2934
R6037 VSS.n9573 VSS.n9529 18.2934
R6038 VSS.n9507 VSS.n9477 18.2934
R6039 VSS.n9673 VSS.n9452 18.2934
R6040 VSS.n9725 VSS.n9416 18.2934
R6041 VSS.n16511 VSS.n16469 18.2934
R6042 VSS.n16564 VSS.n16433 18.2934
R6043 VSS.n16616 VSS.n16394 18.2934
R6044 VSS.n16668 VSS.n16358 18.2934
R6045 VSS.n1676 VSS.n1634 18.2934
R6046 VSS.n1729 VSS.n1598 18.2934
R6047 VSS.n16023 VSS.n1566 18.2934
R6048 VSS.n16075 VSS.n1530 18.2934
R6049 VSS.n1865 VSS.n1821 18.2934
R6050 VSS.n1799 VSS.n1769 18.2934
R6051 VSS.n2026 VSS.n1998 18.2934
R6052 VSS.n2054 VSS.n1989 18.2934
R6053 VSS.n3064 VSS.n3020 18.2934
R6054 VSS.n2998 VSS.n2968 18.2934
R6055 VSS.n3164 VSS.n2943 18.2934
R6056 VSS.n3216 VSS.n2907 18.2934
R6057 VSS.n3656 VSS.n3612 18.2934
R6058 VSS.n3590 VSS.n3560 18.2934
R6059 VSS.n3756 VSS.n3535 18.2934
R6060 VSS.n3808 VSS.n3499 18.2934
R6061 VSS.n4248 VSS.n4204 18.2934
R6062 VSS.n4182 VSS.n4152 18.2934
R6063 VSS.n4348 VSS.n4127 18.2934
R6064 VSS.n4400 VSS.n4091 18.2934
R6065 VSS.n4840 VSS.n4796 18.2934
R6066 VSS.n4774 VSS.n4744 18.2934
R6067 VSS.n4940 VSS.n4719 18.2934
R6068 VSS.n4992 VSS.n4683 18.2934
R6069 VSS.n2461 VSS.n2417 18.2934
R6070 VSS.n2395 VSS.n2365 18.2934
R6071 VSS.n2622 VSS.n2594 18.2934
R6072 VSS.n2650 VSS.n2585 18.2934
R6073 VSS.n5422 VSS.n5378 18.2934
R6074 VSS.n5356 VSS.n5326 18.2934
R6075 VSS.n5583 VSS.n5555 18.2934
R6076 VSS.n5611 VSS.n5546 18.2934
R6077 VSS.n5995 VSS.n5951 18.2934
R6078 VSS.n5929 VSS.n5899 18.2934
R6079 VSS.n6156 VSS.n6128 18.2934
R6080 VSS.n6184 VSS.n6119 18.2934
R6081 VSS.n7797 VSS.n7753 18.2934
R6082 VSS.n7731 VSS.n7701 18.2934
R6083 VSS.n7897 VSS.n7676 18.2934
R6084 VSS.n7949 VSS.n7640 18.2934
R6085 VSS.n8389 VSS.n8345 18.2934
R6086 VSS.n8323 VSS.n8293 18.2934
R6087 VSS.n8489 VSS.n8268 18.2934
R6088 VSS.n8541 VSS.n8232 18.2934
R6089 VSS.n8981 VSS.n8937 18.2934
R6090 VSS.n8915 VSS.n8885 18.2934
R6091 VSS.n9081 VSS.n8860 18.2934
R6092 VSS.n9133 VSS.n8824 18.2934
R6093 VSS.n10165 VSS.n10121 18.2934
R6094 VSS.n10099 VSS.n10069 18.2934
R6095 VSS.n10265 VSS.n10044 18.2934
R6096 VSS.n10317 VSS.n10008 18.2934
R6097 VSS.n10757 VSS.n10713 18.2934
R6098 VSS.n10691 VSS.n10661 18.2934
R6099 VSS.n10857 VSS.n10636 18.2934
R6100 VSS.n10909 VSS.n10600 18.2934
R6101 VSS.n11349 VSS.n11305 18.2934
R6102 VSS.n11283 VSS.n11253 18.2934
R6103 VSS.n11449 VSS.n11228 18.2934
R6104 VSS.n11501 VSS.n11192 18.2934
R6105 VSS.n11941 VSS.n11897 18.2934
R6106 VSS.n11875 VSS.n11845 18.2934
R6107 VSS.n12041 VSS.n11820 18.2934
R6108 VSS.n12093 VSS.n11784 18.2934
R6109 VSS.n12533 VSS.n12489 18.2934
R6110 VSS.n12467 VSS.n12437 18.2934
R6111 VSS.n12633 VSS.n12412 18.2934
R6112 VSS.n12685 VSS.n12376 18.2934
R6113 VSS.n13125 VSS.n13081 18.2934
R6114 VSS.n13059 VSS.n13029 18.2934
R6115 VSS.n13225 VSS.n13004 18.2934
R6116 VSS.n13277 VSS.n12968 18.2934
R6117 VSS.n13717 VSS.n13673 18.2934
R6118 VSS.n13651 VSS.n13621 18.2934
R6119 VSS.n13817 VSS.n13596 18.2934
R6120 VSS.n13869 VSS.n13560 18.2934
R6121 VSS.n14309 VSS.n14265 18.2934
R6122 VSS.n14243 VSS.n14213 18.2934
R6123 VSS.n14409 VSS.n14188 18.2934
R6124 VSS.n14461 VSS.n14152 18.2934
R6125 VSS.n14901 VSS.n14857 18.2934
R6126 VSS.n14835 VSS.n14805 18.2934
R6127 VSS.n15001 VSS.n14780 18.2934
R6128 VSS.n15053 VSS.n14744 18.2934
R6129 VSS.n15493 VSS.n15449 18.2934
R6130 VSS.n15427 VSS.n15397 18.2934
R6131 VSS.n15593 VSS.n15372 18.2934
R6132 VSS.n15645 VSS.n15336 18.2934
R6133 VSS.n6601 VSS.n6557 18.2934
R6134 VSS.n6535 VSS.n6505 18.2934
R6135 VSS.n6762 VSS.n6734 18.2934
R6136 VSS.n6790 VSS.n6725 18.2934
R6137 VSS.n7200 VSS.n7158 18.2934
R6138 VSS.n7253 VSS.n7122 18.2934
R6139 VSS.n7305 VSS.n7083 18.2934
R6140 VSS.n7357 VSS.n7047 18.2934
R6141 VSS.n362 VSS.n341 18.2934
R6142 VSS.n398 VSS.n331 18.2934
R6143 VSS.n18617 VSS.n181 18.2934
R6144 VSS.n18669 VSS.n145 18.2934
R6145 VSS.n585 VSS.n554 18.2934
R6146 VSS.n613 VSS.n545 18.2934
R6147 VSS.t12 VSS.t51 17.244
R6148 VSS.t0 VSS.t1 16.3482
R6149 VSS.t51 VSS.t0 16.1243
R6150 VSS.n1220 VSS.n1157 15.4791
R6151 VSS.n1285 VSS.n1198 15.4791
R6152 VSS.n17499 VSS.n17495 15.4791
R6153 VSS.n17593 VSS.n17426 15.4791
R6154 VSS.n1087 VSS.n1022 15.4791
R6155 VSS.n1151 VSS.n1064 15.4791
R6156 VSS.n906 VSS.n455 15.4791
R6157 VSS.n970 VSS.n883 15.4791
R6158 VSS.n17004 VSS.n16989 15.4791
R6159 VSS.n17102 VSS.n16937 15.4791
R6160 VSS.n17418 VSS.n17403 15.4791
R6161 VSS.n17694 VSS.n17351 15.4791
R6162 VSS.n18237 VSS.n210 15.4791
R6163 VSS.n18302 VSS.n18215 15.4791
R6164 VSS.n18076 VSS.n287 15.4791
R6165 VSS.n18170 VSS.n218 15.4791
R6166 VSS.n9549 VSS.n9545 15.4791
R6167 VSS.n9643 VSS.n9476 15.4791
R6168 VSS.n9468 VSS.n9453 15.4791
R6169 VSS.n9744 VSS.n9401 15.4791
R6170 VSS.n16485 VSS.n16470 15.4791
R6171 VSS.n16583 VSS.n16418 15.4791
R6172 VSS.n16410 VSS.n16395 15.4791
R6173 VSS.n16687 VSS.n16343 15.4791
R6174 VSS.n1650 VSS.n1635 15.4791
R6175 VSS.n1748 VSS.n1583 15.4791
R6176 VSS.n1755 VSS.n1567 15.4791
R6177 VSS.n16094 VSS.n1515 15.4791
R6178 VSS.n1841 VSS.n1837 15.4791
R6179 VSS.n1935 VSS.n1768 15.4791
R6180 VSS.n2002 VSS.n1760 15.4791
R6181 VSS.n2067 VSS.n1980 15.4791
R6182 VSS.n3040 VSS.n3036 15.4791
R6183 VSS.n3134 VSS.n2967 15.4791
R6184 VSS.n2959 VSS.n2944 15.4791
R6185 VSS.n3235 VSS.n2892 15.4791
R6186 VSS.n3632 VSS.n3628 15.4791
R6187 VSS.n3726 VSS.n3559 15.4791
R6188 VSS.n3551 VSS.n3536 15.4791
R6189 VSS.n3827 VSS.n3484 15.4791
R6190 VSS.n4224 VSS.n4220 15.4791
R6191 VSS.n4318 VSS.n4151 15.4791
R6192 VSS.n4143 VSS.n4128 15.4791
R6193 VSS.n4419 VSS.n4076 15.4791
R6194 VSS.n4816 VSS.n4812 15.4791
R6195 VSS.n4910 VSS.n4743 15.4791
R6196 VSS.n4735 VSS.n4720 15.4791
R6197 VSS.n5011 VSS.n4668 15.4791
R6198 VSS.n2437 VSS.n2433 15.4791
R6199 VSS.n2531 VSS.n2364 15.4791
R6200 VSS.n2598 VSS.n2356 15.4791
R6201 VSS.n2663 VSS.n2576 15.4791
R6202 VSS.n5398 VSS.n5394 15.4791
R6203 VSS.n5492 VSS.n5325 15.4791
R6204 VSS.n5559 VSS.n5317 15.4791
R6205 VSS.n5624 VSS.n5537 15.4791
R6206 VSS.n5971 VSS.n5967 15.4791
R6207 VSS.n6065 VSS.n5898 15.4791
R6208 VSS.n6132 VSS.n5890 15.4791
R6209 VSS.n6197 VSS.n6110 15.4791
R6210 VSS.n7773 VSS.n7769 15.4791
R6211 VSS.n7867 VSS.n7700 15.4791
R6212 VSS.n7692 VSS.n7677 15.4791
R6213 VSS.n7968 VSS.n7625 15.4791
R6214 VSS.n8365 VSS.n8361 15.4791
R6215 VSS.n8459 VSS.n8292 15.4791
R6216 VSS.n8284 VSS.n8269 15.4791
R6217 VSS.n8560 VSS.n8217 15.4791
R6218 VSS.n8957 VSS.n8953 15.4791
R6219 VSS.n9051 VSS.n8884 15.4791
R6220 VSS.n8876 VSS.n8861 15.4791
R6221 VSS.n9152 VSS.n8809 15.4791
R6222 VSS.n10141 VSS.n10137 15.4791
R6223 VSS.n10235 VSS.n10068 15.4791
R6224 VSS.n10060 VSS.n10045 15.4791
R6225 VSS.n10336 VSS.n9993 15.4791
R6226 VSS.n10733 VSS.n10729 15.4791
R6227 VSS.n10827 VSS.n10660 15.4791
R6228 VSS.n10652 VSS.n10637 15.4791
R6229 VSS.n10928 VSS.n10585 15.4791
R6230 VSS.n11325 VSS.n11321 15.4791
R6231 VSS.n11419 VSS.n11252 15.4791
R6232 VSS.n11244 VSS.n11229 15.4791
R6233 VSS.n11520 VSS.n11177 15.4791
R6234 VSS.n11917 VSS.n11913 15.4791
R6235 VSS.n12011 VSS.n11844 15.4791
R6236 VSS.n11836 VSS.n11821 15.4791
R6237 VSS.n12112 VSS.n11769 15.4791
R6238 VSS.n12509 VSS.n12505 15.4791
R6239 VSS.n12603 VSS.n12436 15.4791
R6240 VSS.n12428 VSS.n12413 15.4791
R6241 VSS.n12704 VSS.n12361 15.4791
R6242 VSS.n13101 VSS.n13097 15.4791
R6243 VSS.n13195 VSS.n13028 15.4791
R6244 VSS.n13020 VSS.n13005 15.4791
R6245 VSS.n13296 VSS.n12953 15.4791
R6246 VSS.n13693 VSS.n13689 15.4791
R6247 VSS.n13787 VSS.n13620 15.4791
R6248 VSS.n13612 VSS.n13597 15.4791
R6249 VSS.n13888 VSS.n13545 15.4791
R6250 VSS.n14285 VSS.n14281 15.4791
R6251 VSS.n14379 VSS.n14212 15.4791
R6252 VSS.n14204 VSS.n14189 15.4791
R6253 VSS.n14480 VSS.n14137 15.4791
R6254 VSS.n14877 VSS.n14873 15.4791
R6255 VSS.n14971 VSS.n14804 15.4791
R6256 VSS.n14796 VSS.n14781 15.4791
R6257 VSS.n15072 VSS.n14729 15.4791
R6258 VSS.n15469 VSS.n15465 15.4791
R6259 VSS.n15563 VSS.n15396 15.4791
R6260 VSS.n15388 VSS.n15373 15.4791
R6261 VSS.n15664 VSS.n15321 15.4791
R6262 VSS.n6577 VSS.n6573 15.4791
R6263 VSS.n6671 VSS.n6504 15.4791
R6264 VSS.n6738 VSS.n6496 15.4791
R6265 VSS.n6803 VSS.n6716 15.4791
R6266 VSS.n7174 VSS.n7159 15.4791
R6267 VSS.n7272 VSS.n7107 15.4791
R6268 VSS.n7099 VSS.n7084 15.4791
R6269 VSS.n7376 VSS.n7032 15.4791
R6270 VSS.n358 VSS.n289 15.4791
R6271 VSS.n402 VSS.n198 15.4791
R6272 VSS.n204 VSS.n182 15.4791
R6273 VSS.n18688 VSS.n130 15.4791
R6274 VSS.n563 VSS.n558 15.4791
R6275 VSS.n626 VSS.n536 15.4791
R6276 VSS.n17121 VSS.n17106 15.3911
R6277 VSS.n17265 VSS.n16867 15.3911
R6278 VSS.n17713 VSS.n17698 15.3911
R6279 VSS.n17857 VSS.n17281 15.3911
R6280 VSS.n18533 VSS.n18306 15.3911
R6281 VSS.n18461 VSS.n18438 15.3911
R6282 VSS.n9763 VSS.n9748 15.3911
R6283 VSS.n9908 VSS.n9332 15.3911
R6284 VSS.n16706 VSS.n16691 15.3911
R6285 VSS.n16851 VSS.n16274 15.3911
R6286 VSS.n16113 VSS.n16098 15.3911
R6287 VSS.n16258 VSS.n1446 15.3911
R6288 VSS.n2298 VSS.n2071 15.3911
R6289 VSS.n2204 VSS.n2198 15.3911
R6290 VSS.n3254 VSS.n3239 15.3911
R6291 VSS.n3399 VSS.n2823 15.3911
R6292 VSS.n3846 VSS.n3831 15.3911
R6293 VSS.n3991 VSS.n3415 15.3911
R6294 VSS.n4438 VSS.n4423 15.3911
R6295 VSS.n4583 VSS.n4007 15.3911
R6296 VSS.n5030 VSS.n5015 15.3911
R6297 VSS.n5175 VSS.n4599 15.3911
R6298 VSS.n5263 VSS.n2667 15.3911
R6299 VSS.n2800 VSS.n2794 15.3911
R6300 VSS.n5836 VSS.n5628 15.3911
R6301 VSS.n18881 VSS.n8 15.3911
R6302 VSS.n6428 VSS.n6201 15.3911
R6303 VSS.n6334 VSS.n6328 15.3911
R6304 VSS.n7987 VSS.n7972 15.3911
R6305 VSS.n8132 VSS.n7556 15.3911
R6306 VSS.n8579 VSS.n8564 15.3911
R6307 VSS.n8724 VSS.n8148 15.3911
R6308 VSS.n9171 VSS.n9156 15.3911
R6309 VSS.n9316 VSS.n8740 15.3911
R6310 VSS.n10355 VSS.n10340 15.3911
R6311 VSS.n10500 VSS.n9924 15.3911
R6312 VSS.n10947 VSS.n10932 15.3911
R6313 VSS.n11092 VSS.n10516 15.3911
R6314 VSS.n11539 VSS.n11524 15.3911
R6315 VSS.n11684 VSS.n11108 15.3911
R6316 VSS.n12131 VSS.n12116 15.3911
R6317 VSS.n12276 VSS.n11700 15.3911
R6318 VSS.n12723 VSS.n12708 15.3911
R6319 VSS.n12868 VSS.n12292 15.3911
R6320 VSS.n13315 VSS.n13300 15.3911
R6321 VSS.n13460 VSS.n12884 15.3911
R6322 VSS.n13907 VSS.n13892 15.3911
R6323 VSS.n14052 VSS.n13476 15.3911
R6324 VSS.n14499 VSS.n14484 15.3911
R6325 VSS.n14644 VSS.n14068 15.3911
R6326 VSS.n15091 VSS.n15076 15.3911
R6327 VSS.n15236 VSS.n14660 15.3911
R6328 VSS.n15683 VSS.n15668 15.3911
R6329 VSS.n15828 VSS.n15252 15.3911
R6330 VSS.n15916 VSS.n6807 15.3911
R6331 VSS.n6940 VSS.n6934 15.3911
R6332 VSS.n7395 VSS.n7380 15.3911
R6333 VSS.n7540 VSS.n6963 15.3911
R6334 VSS.n18707 VSS.n18692 15.3911
R6335 VSS.n18852 VSS.n61 15.3911
R6336 VSS.n830 VSS.n630 15.3911
R6337 VSS.n18873 VSS.n42 15.3911
R6338 VSS.n17944 VSS.n1289 15.3911
R6339 VSS.n1422 VSS.n1416 15.3911
R6340 VSS.n1247 VSS.n1212 14.9665
R6341 VSS.n1270 VSS.n1208 14.9665
R6342 VSS.n17498 VSS.n17496 14.5379
R6343 VSS.n17592 VSS.n1155 14.5379
R6344 VSS.n10171 VSS.n10170 12.4475
R6345 VSS.n10204 VSS.n10201 12.4475
R6346 VSS.n17050 VSS.n16974 12.4299
R6347 VSS.n17081 VSS.n16953 12.4299
R6348 VSS.n17642 VSS.n17388 12.4299
R6349 VSS.n17673 VSS.n17367 12.4299
R6350 VSS.n18106 VSS.n18105 12.4299
R6351 VSS.n18139 VSS.n18136 12.4299
R6352 VSS.n9692 VSS.n9438 12.4299
R6353 VSS.n9723 VSS.n9417 12.4299
R6354 VSS.n16635 VSS.n16380 12.4299
R6355 VSS.n16666 VSS.n16359 12.4299
R6356 VSS.n16530 VSS.n16457 12.4299
R6357 VSS.n16561 VSS.n16434 12.4299
R6358 VSS.n16042 VSS.n1552 12.4299
R6359 VSS.n16073 VSS.n1531 12.4299
R6360 VSS.n1695 VSS.n1622 12.4299
R6361 VSS.n1726 VSS.n1599 12.4299
R6362 VSS.n2029 VSS.n1994 12.4299
R6363 VSS.n2052 VSS.n1990 12.4299
R6364 VSS.n1871 VSS.n1870 12.4299
R6365 VSS.n1904 VSS.n1901 12.4299
R6366 VSS.n3183 VSS.n2929 12.4299
R6367 VSS.n3214 VSS.n2908 12.4299
R6368 VSS.n3070 VSS.n3069 12.4299
R6369 VSS.n3103 VSS.n3100 12.4299
R6370 VSS.n3775 VSS.n3521 12.4299
R6371 VSS.n3806 VSS.n3500 12.4299
R6372 VSS.n3662 VSS.n3661 12.4299
R6373 VSS.n3695 VSS.n3692 12.4299
R6374 VSS.n4367 VSS.n4113 12.4299
R6375 VSS.n4398 VSS.n4092 12.4299
R6376 VSS.n4254 VSS.n4253 12.4299
R6377 VSS.n4287 VSS.n4284 12.4299
R6378 VSS.n4959 VSS.n4705 12.4299
R6379 VSS.n4990 VSS.n4684 12.4299
R6380 VSS.n4846 VSS.n4845 12.4299
R6381 VSS.n4879 VSS.n4876 12.4299
R6382 VSS.n2625 VSS.n2590 12.4299
R6383 VSS.n2648 VSS.n2586 12.4299
R6384 VSS.n2467 VSS.n2466 12.4299
R6385 VSS.n2500 VSS.n2497 12.4299
R6386 VSS.n5586 VSS.n5551 12.4299
R6387 VSS.n5609 VSS.n5547 12.4299
R6388 VSS.n5428 VSS.n5427 12.4299
R6389 VSS.n5461 VSS.n5458 12.4299
R6390 VSS.n6159 VSS.n6124 12.4299
R6391 VSS.n6182 VSS.n6120 12.4299
R6392 VSS.n6001 VSS.n6000 12.4299
R6393 VSS.n6034 VSS.n6031 12.4299
R6394 VSS.n7916 VSS.n7662 12.4299
R6395 VSS.n7947 VSS.n7641 12.4299
R6396 VSS.n7803 VSS.n7802 12.4299
R6397 VSS.n7836 VSS.n7833 12.4299
R6398 VSS.n8508 VSS.n8254 12.4299
R6399 VSS.n8539 VSS.n8233 12.4299
R6400 VSS.n8395 VSS.n8394 12.4299
R6401 VSS.n8428 VSS.n8425 12.4299
R6402 VSS.n9100 VSS.n8846 12.4299
R6403 VSS.n9131 VSS.n8825 12.4299
R6404 VSS.n8987 VSS.n8986 12.4299
R6405 VSS.n9020 VSS.n9017 12.4299
R6406 VSS.n10284 VSS.n10030 12.4299
R6407 VSS.n10315 VSS.n10009 12.4299
R6408 VSS.n10876 VSS.n10622 12.4299
R6409 VSS.n10907 VSS.n10601 12.4299
R6410 VSS.n10763 VSS.n10762 12.4299
R6411 VSS.n10796 VSS.n10793 12.4299
R6412 VSS.n11468 VSS.n11214 12.4299
R6413 VSS.n11499 VSS.n11193 12.4299
R6414 VSS.n11355 VSS.n11354 12.4299
R6415 VSS.n11388 VSS.n11385 12.4299
R6416 VSS.n12060 VSS.n11806 12.4299
R6417 VSS.n12091 VSS.n11785 12.4299
R6418 VSS.n11947 VSS.n11946 12.4299
R6419 VSS.n11980 VSS.n11977 12.4299
R6420 VSS.n12652 VSS.n12398 12.4299
R6421 VSS.n12683 VSS.n12377 12.4299
R6422 VSS.n12539 VSS.n12538 12.4299
R6423 VSS.n12572 VSS.n12569 12.4299
R6424 VSS.n13244 VSS.n12990 12.4299
R6425 VSS.n13275 VSS.n12969 12.4299
R6426 VSS.n13131 VSS.n13130 12.4299
R6427 VSS.n13164 VSS.n13161 12.4299
R6428 VSS.n13836 VSS.n13582 12.4299
R6429 VSS.n13867 VSS.n13561 12.4299
R6430 VSS.n13723 VSS.n13722 12.4299
R6431 VSS.n13756 VSS.n13753 12.4299
R6432 VSS.n14428 VSS.n14174 12.4299
R6433 VSS.n14459 VSS.n14153 12.4299
R6434 VSS.n14315 VSS.n14314 12.4299
R6435 VSS.n14348 VSS.n14345 12.4299
R6436 VSS.n15020 VSS.n14766 12.4299
R6437 VSS.n15051 VSS.n14745 12.4299
R6438 VSS.n14907 VSS.n14906 12.4299
R6439 VSS.n14940 VSS.n14937 12.4299
R6440 VSS.n15612 VSS.n15358 12.4299
R6441 VSS.n15643 VSS.n15337 12.4299
R6442 VSS.n15499 VSS.n15498 12.4299
R6443 VSS.n15532 VSS.n15529 12.4299
R6444 VSS.n6765 VSS.n6730 12.4299
R6445 VSS.n6788 VSS.n6726 12.4299
R6446 VSS.n6607 VSS.n6606 12.4299
R6447 VSS.n6640 VSS.n6637 12.4299
R6448 VSS.n7324 VSS.n7069 12.4299
R6449 VSS.n7355 VSS.n7048 12.4299
R6450 VSS.n7219 VSS.n7146 12.4299
R6451 VSS.n7250 VSS.n7123 12.4299
R6452 VSS.n18636 VSS.n167 12.4299
R6453 VSS.n18667 VSS.n146 12.4299
R6454 VSS.n374 VSS.n373 12.4299
R6455 VSS.n384 VSS.n383 12.4299
R6456 VSS.n18264 VSS.n18229 12.4299
R6457 VSS.n18287 VSS.n18225 12.4299
R6458 VSS.n588 VSS.n550 12.4299
R6459 VSS.n611 VSS.n546 12.4299
R6460 VSS.n931 VSS.n898 12.4299
R6461 VSS.n954 VSS.n893 12.4299
R6462 VSS.n1112 VSS.n1079 12.4299
R6463 VSS.n1135 VSS.n1074 12.4299
R6464 VSS.n9579 VSS.n9578 12.4123
R6465 VSS.n9612 VSS.n9609 12.4123
R6466 VSS.n17524 VSS.n17481 9.69213
R6467 VSS.n17994 VSS.n17993 9.38145
R6468 VSS.n18043 VSS.n18042 9.38145
R6469 VSS.n17006 VSS.n16999 9.38145
R6470 VSS.n17501 VSS.n17493 9.38145
R6471 VSS.n17420 VSS.n17413 9.38145
R6472 VSS.n18583 VSS.n18582 9.38145
R6473 VSS.n18078 VSS.n285 9.38145
R6474 VSS.n9470 VSS.n9463 9.38145
R6475 VSS.n9551 VSS.n9543 9.38145
R6476 VSS.n16412 VSS.n16405 9.38145
R6477 VSS.n16487 VSS.n16480 9.38145
R6478 VSS.n1756 VSS.n1577 9.38145
R6479 VSS.n1652 VSS.n1645 9.38145
R6480 VSS.n2348 VSS.n2347 9.38145
R6481 VSS.n1843 VSS.n1835 9.38145
R6482 VSS.n2961 VSS.n2954 9.38145
R6483 VSS.n3042 VSS.n3034 9.38145
R6484 VSS.n3553 VSS.n3546 9.38145
R6485 VSS.n3634 VSS.n3626 9.38145
R6486 VSS.n4145 VSS.n4138 9.38145
R6487 VSS.n4226 VSS.n4218 9.38145
R6488 VSS.n4737 VSS.n4730 9.38145
R6489 VSS.n4818 VSS.n4810 9.38145
R6490 VSS.n5313 VSS.n5312 9.38145
R6491 VSS.n2439 VSS.n2431 9.38145
R6492 VSS.n5886 VSS.n5885 9.38145
R6493 VSS.n5400 VSS.n5392 9.38145
R6494 VSS.n6478 VSS.n6477 9.38145
R6495 VSS.n5973 VSS.n5965 9.38145
R6496 VSS.n7694 VSS.n7687 9.38145
R6497 VSS.n7775 VSS.n7767 9.38145
R6498 VSS.n8286 VSS.n8279 9.38145
R6499 VSS.n8367 VSS.n8359 9.38145
R6500 VSS.n8878 VSS.n8871 9.38145
R6501 VSS.n8959 VSS.n8951 9.38145
R6502 VSS.n10062 VSS.n10055 9.38145
R6503 VSS.n10143 VSS.n10135 9.38145
R6504 VSS.n10654 VSS.n10647 9.38145
R6505 VSS.n10735 VSS.n10727 9.38145
R6506 VSS.n11246 VSS.n11239 9.38145
R6507 VSS.n11327 VSS.n11319 9.38145
R6508 VSS.n11838 VSS.n11831 9.38145
R6509 VSS.n11919 VSS.n11911 9.38145
R6510 VSS.n12430 VSS.n12423 9.38145
R6511 VSS.n12511 VSS.n12503 9.38145
R6512 VSS.n13022 VSS.n13015 9.38145
R6513 VSS.n13103 VSS.n13095 9.38145
R6514 VSS.n13614 VSS.n13607 9.38145
R6515 VSS.n13695 VSS.n13687 9.38145
R6516 VSS.n14206 VSS.n14199 9.38145
R6517 VSS.n14287 VSS.n14279 9.38145
R6518 VSS.n14798 VSS.n14791 9.38145
R6519 VSS.n14879 VSS.n14871 9.38145
R6520 VSS.n15390 VSS.n15383 9.38145
R6521 VSS.n15471 VSS.n15463 9.38145
R6522 VSS.n15966 VSS.n15965 9.38145
R6523 VSS.n6579 VSS.n6571 9.38145
R6524 VSS.n7101 VSS.n7094 9.38145
R6525 VSS.n7176 VSS.n7169 9.38145
R6526 VSS.n205 VSS.n192 9.38145
R6527 VSS.n452 VSS.n451 9.38145
R6528 VSS.n559 VSS.n497 9.38145
R6529 VSS.n1017 VSS.n1016 9.38145
R6530 VSS.n17266 VSS.n16862 9.30555
R6531 VSS.n17122 VSS.n17110 9.30555
R6532 VSS.n17858 VSS.n17276 9.30555
R6533 VSS.n17714 VSS.n17702 9.30555
R6534 VSS.n18462 VSS.n18432 9.30555
R6535 VSS.n18534 VSS.n18308 9.30555
R6536 VSS.n9909 VSS.n9327 9.30555
R6537 VSS.n9764 VSS.n9752 9.30555
R6538 VSS.n16852 VSS.n16269 9.30555
R6539 VSS.n16707 VSS.n16695 9.30555
R6540 VSS.n16259 VSS.n1441 9.30555
R6541 VSS.n16114 VSS.n16102 9.30555
R6542 VSS.n2207 VSS.n2206 9.30555
R6543 VSS.n2299 VSS.n2073 9.30555
R6544 VSS.n3400 VSS.n2818 9.30555
R6545 VSS.n3255 VSS.n3243 9.30555
R6546 VSS.n3992 VSS.n3410 9.30555
R6547 VSS.n3847 VSS.n3835 9.30555
R6548 VSS.n4584 VSS.n4002 9.30555
R6549 VSS.n4439 VSS.n4427 9.30555
R6550 VSS.n5176 VSS.n4594 9.30555
R6551 VSS.n5031 VSS.n5019 9.30555
R6552 VSS.n2803 VSS.n2802 9.30555
R6553 VSS.n5264 VSS.n2669 9.30555
R6554 VSS.n18882 VSS.n3 9.30555
R6555 VSS.n5837 VSS.n5630 9.30555
R6556 VSS.n6337 VSS.n6336 9.30555
R6557 VSS.n6429 VSS.n6203 9.30555
R6558 VSS.n8133 VSS.n7551 9.30555
R6559 VSS.n7988 VSS.n7976 9.30555
R6560 VSS.n8725 VSS.n8143 9.30555
R6561 VSS.n8580 VSS.n8568 9.30555
R6562 VSS.n9317 VSS.n8735 9.30555
R6563 VSS.n9172 VSS.n9160 9.30555
R6564 VSS.n10501 VSS.n9919 9.30555
R6565 VSS.n10356 VSS.n10344 9.30555
R6566 VSS.n11093 VSS.n10511 9.30555
R6567 VSS.n10948 VSS.n10936 9.30555
R6568 VSS.n11685 VSS.n11103 9.30555
R6569 VSS.n11540 VSS.n11528 9.30555
R6570 VSS.n12277 VSS.n11695 9.30555
R6571 VSS.n12132 VSS.n12120 9.30555
R6572 VSS.n12869 VSS.n12287 9.30555
R6573 VSS.n12724 VSS.n12712 9.30555
R6574 VSS.n13461 VSS.n12879 9.30555
R6575 VSS.n13316 VSS.n13304 9.30555
R6576 VSS.n14053 VSS.n13471 9.30555
R6577 VSS.n13908 VSS.n13896 9.30555
R6578 VSS.n14645 VSS.n14063 9.30555
R6579 VSS.n14500 VSS.n14488 9.30555
R6580 VSS.n15237 VSS.n14655 9.30555
R6581 VSS.n15092 VSS.n15080 9.30555
R6582 VSS.n15829 VSS.n15247 9.30555
R6583 VSS.n15684 VSS.n15672 9.30555
R6584 VSS.n6943 VSS.n6942 9.30555
R6585 VSS.n15917 VSS.n6809 9.30555
R6586 VSS.n7541 VSS.n6958 9.30555
R6587 VSS.n7396 VSS.n7384 9.30555
R6588 VSS.n18853 VSS.n56 9.30555
R6589 VSS.n18708 VSS.n18696 9.30555
R6590 VSS.n18874 VSS.n44 9.30555
R6591 VSS.n831 VSS.n632 9.30555
R6592 VSS.n1425 VSS.n1424 9.30555
R6593 VSS.n17945 VSS.n1291 9.30555
R6594 VSS.n1241 VSS.n1240 9.3005
R6595 VSS.n1262 VSS.n1261 9.3005
R6596 VSS.n1202 VSS.n1201 9.3005
R6597 VSS.n1283 VSS.n1282 9.3005
R6598 VSS.n1106 VSS.n1105 9.3005
R6599 VSS.n1127 VSS.n1126 9.3005
R6600 VSS.n1068 VSS.n1067 9.3005
R6601 VSS.n1149 VSS.n1148 9.3005
R6602 VSS.n17171 VSS.n17170 9.3005
R6603 VSS.n16864 VSS.n16863 9.3005
R6604 VSS.n17221 VSS.n16890 9.3005
R6605 VSS.n16898 VSS.n16896 9.3005
R6606 VSS.n17186 VSS.n17185 9.3005
R6607 VSS.n17240 VSS.n16878 9.3005
R6608 VSS.n17242 VSS.n17241 9.3005
R6609 VSS.n17224 VSS.n17222 9.3005
R6610 VSS.n17172 VSS.n16910 9.3005
R6611 VSS.n17184 VSS.n16903 9.3005
R6612 VSS.n17199 VSS.n17198 9.3005
R6613 VSS.n17114 VSS.n16930 9.3005
R6614 VSS.n17151 VSS.n16921 9.3005
R6615 VSS.n17153 VSS.n17152 9.3005
R6616 VSS.n17034 VSS.n17033 9.3005
R6617 VSS.n17072 VSS.n17071 9.3005
R6618 VSS.n16941 VSS.n16940 9.3005
R6619 VSS.n17100 VSS.n17099 9.3005
R6620 VSS.n17079 VSS.n17078 9.3005
R6621 VSS.n17080 VSS.n17079 9.3005
R6622 VSS.n17081 VSS.n17080 9.3005
R6623 VSS.n17047 VSS.n17046 9.3005
R6624 VSS.n17047 VSS.n16975 9.3005
R6625 VSS.n16975 VSS.n16974 9.3005
R6626 VSS.n17027 VSS.n17026 9.3005
R6627 VSS.n17028 VSS.n17027 9.3005
R6628 VSS.n17087 VSS.n17086 9.3005
R6629 VSS.n17086 VSS.n16939 9.3005
R6630 VSS.n16939 VSS.n16938 9.3005
R6631 VSS.n17129 VSS.n17128 9.3005
R6632 VSS.n17128 VSS.n17127 9.3005
R6633 VSS.n17001 VSS.n16999 9.3005
R6634 VSS.n17257 VSS.n17256 9.3005
R6635 VSS.n17257 VSS.n16869 9.3005
R6636 VSS.n16869 VSS.n16868 9.3005
R6637 VSS.n17234 VSS.n17233 9.3005
R6638 VSS.n17235 VSS.n17234 9.3005
R6639 VSS.n17236 VSS.n17235 9.3005
R6640 VSS.n17202 VSS.n16891 9.3005
R6641 VSS.n16892 VSS.n16891 9.3005
R6642 VSS.n17216 VSS.n16892 9.3005
R6643 VSS.n17161 VSS.n17160 9.3005
R6644 VSS.n17161 VSS.n16913 9.3005
R6645 VSS.n17165 VSS.n16913 9.3005
R6646 VSS.n17181 VSS.n16904 9.3005
R6647 VSS.n16904 VSS.n16894 9.3005
R6648 VSS.n16894 VSS.n16893 9.3005
R6649 VSS.n17266 VSS.n17265 9.3005
R6650 VSS.n17265 VSS.n17264 9.3005
R6651 VSS.n17122 VSS.n17121 9.3005
R6652 VSS.n17121 VSS.n17120 9.3005
R6653 VSS.n16923 VSS.n16922 9.3005
R6654 VSS.n17113 VSS.n16922 9.3005
R6655 VSS.n17113 VSS.n17112 9.3005
R6656 VSS.n17477 VSS.n17473 9.3005
R6657 VSS.n17455 VSS.n17454 9.3005
R6658 VSS.n17435 VSS.n17434 9.3005
R6659 VSS.n17438 VSS.n17437 9.3005
R6660 VSS.n17763 VSS.n17762 9.3005
R6661 VSS.n17278 VSS.n17277 9.3005
R6662 VSS.n17813 VSS.n17304 9.3005
R6663 VSS.n17312 VSS.n17310 9.3005
R6664 VSS.n17778 VSS.n17777 9.3005
R6665 VSS.n17832 VSS.n17292 9.3005
R6666 VSS.n17834 VSS.n17833 9.3005
R6667 VSS.n17816 VSS.n17814 9.3005
R6668 VSS.n17764 VSS.n17324 9.3005
R6669 VSS.n17776 VSS.n17317 9.3005
R6670 VSS.n17791 VSS.n17790 9.3005
R6671 VSS.n17706 VSS.n17344 9.3005
R6672 VSS.n17743 VSS.n17335 9.3005
R6673 VSS.n17745 VSS.n17744 9.3005
R6674 VSS.n17626 VSS.n17625 9.3005
R6675 VSS.n17664 VSS.n17663 9.3005
R6676 VSS.n17355 VSS.n17354 9.3005
R6677 VSS.n17692 VSS.n17691 9.3005
R6678 VSS.n17671 VSS.n17670 9.3005
R6679 VSS.n17672 VSS.n17671 9.3005
R6680 VSS.n17673 VSS.n17672 9.3005
R6681 VSS.n17639 VSS.n17638 9.3005
R6682 VSS.n17639 VSS.n17389 9.3005
R6683 VSS.n17389 VSS.n17388 9.3005
R6684 VSS.n17619 VSS.n17618 9.3005
R6685 VSS.n17620 VSS.n17619 9.3005
R6686 VSS.n17679 VSS.n17678 9.3005
R6687 VSS.n17678 VSS.n17353 9.3005
R6688 VSS.n17353 VSS.n17352 9.3005
R6689 VSS.n17721 VSS.n17720 9.3005
R6690 VSS.n17720 VSS.n17719 9.3005
R6691 VSS.n17415 VSS.n17413 9.3005
R6692 VSS.n17849 VSS.n17848 9.3005
R6693 VSS.n17849 VSS.n17283 9.3005
R6694 VSS.n17283 VSS.n17282 9.3005
R6695 VSS.n17826 VSS.n17825 9.3005
R6696 VSS.n17827 VSS.n17826 9.3005
R6697 VSS.n17828 VSS.n17827 9.3005
R6698 VSS.n17794 VSS.n17305 9.3005
R6699 VSS.n17306 VSS.n17305 9.3005
R6700 VSS.n17808 VSS.n17306 9.3005
R6701 VSS.n17753 VSS.n17752 9.3005
R6702 VSS.n17753 VSS.n17327 9.3005
R6703 VSS.n17757 VSS.n17327 9.3005
R6704 VSS.n17773 VSS.n17318 9.3005
R6705 VSS.n17318 VSS.n17308 9.3005
R6706 VSS.n17308 VSS.n17307 9.3005
R6707 VSS.n17858 VSS.n17857 9.3005
R6708 VSS.n17857 VSS.n17856 9.3005
R6709 VSS.n17714 VSS.n17713 9.3005
R6710 VSS.n17713 VSS.n17712 9.3005
R6711 VSS.n17337 VSS.n17336 9.3005
R6712 VSS.n17705 VSS.n17336 9.3005
R6713 VSS.n17705 VSS.n17704 9.3005
R6714 VSS.n18258 VSS.n18257 9.3005
R6715 VSS.n18279 VSS.n18278 9.3005
R6716 VSS.n18219 VSS.n18218 9.3005
R6717 VSS.n18300 VSS.n18299 9.3005
R6718 VSS.n18509 VSS.n18508 9.3005
R6719 VSS.n18435 VSS.n18434 9.3005
R6720 VSS.n18490 VSS.n18489 9.3005
R6721 VSS.n18402 VSS.n18396 9.3005
R6722 VSS.n18357 VSS.n18355 9.3005
R6723 VSS.n18482 VSS.n18481 9.3005
R6724 VSS.n18480 VSS.n18419 9.3005
R6725 VSS.n18488 VSS.n18387 9.3005
R6726 VSS.n18510 VSS.n18342 9.3005
R6727 VSS.n18376 VSS.n18375 9.3005
R6728 VSS.n18404 VSS.n18403 9.3005
R6729 VSS.n18323 VSS.n18322 9.3005
R6730 VSS.n18364 VSS.n18363 9.3005
R6731 VSS.n18365 VSS.n18339 9.3005
R6732 VSS.n269 VSS.n265 9.3005
R6733 VSS.n247 VSS.n246 9.3005
R6734 VSS.n227 VSS.n226 9.3005
R6735 VSS.n230 VSS.n229 9.3005
R6736 VSS.n18142 VSS.n18141 9.3005
R6737 VSS.n18141 VSS.n18140 9.3005
R6738 VSS.n18140 VSS.n18139 9.3005
R6739 VSS.n18108 VSS.n268 9.3005
R6740 VSS.n18108 VSS.n18107 9.3005
R6741 VSS.n18107 VSS.n18106 9.3005
R6742 VSS.n18097 VSS.n274 9.3005
R6743 VSS.n274 VSS.n273 9.3005
R6744 VSS.n18165 VSS.n18164 9.3005
R6745 VSS.n18166 VSS.n18165 9.3005
R6746 VSS.n18167 VSS.n18166 9.3005
R6747 VSS.n18172 VSS.n18171 9.3005
R6748 VSS.n18171 VSS.n208 9.3005
R6749 VSS.n18073 VSS.n285 9.3005
R6750 VSS.n9676 VSS.n9675 9.3005
R6751 VSS.n9714 VSS.n9713 9.3005
R6752 VSS.n9405 VSS.n9404 9.3005
R6753 VSS.n9742 VSS.n9741 9.3005
R6754 VSS.n9721 VSS.n9720 9.3005
R6755 VSS.n9722 VSS.n9721 9.3005
R6756 VSS.n9723 VSS.n9722 9.3005
R6757 VSS.n9689 VSS.n9688 9.3005
R6758 VSS.n9689 VSS.n9439 9.3005
R6759 VSS.n9439 VSS.n9438 9.3005
R6760 VSS.n9669 VSS.n9668 9.3005
R6761 VSS.n9670 VSS.n9669 9.3005
R6762 VSS.n9729 VSS.n9728 9.3005
R6763 VSS.n9728 VSS.n9403 9.3005
R6764 VSS.n9403 VSS.n9402 9.3005
R6765 VSS.n9771 VSS.n9770 9.3005
R6766 VSS.n9770 VSS.n9769 9.3005
R6767 VSS.n9465 VSS.n9463 9.3005
R6768 VSS.n9813 VSS.n9812 9.3005
R6769 VSS.n9329 VSS.n9328 9.3005
R6770 VSS.n9863 VSS.n9354 9.3005
R6771 VSS.n9362 VSS.n9360 9.3005
R6772 VSS.n9828 VSS.n9827 9.3005
R6773 VSS.n9900 VSS.n9899 9.3005
R6774 VSS.n9900 VSS.n9334 9.3005
R6775 VSS.n9334 VSS.n9333 9.3005
R6776 VSS.n9882 VSS.n9342 9.3005
R6777 VSS.n9884 VSS.n9883 9.3005
R6778 VSS.n9876 VSS.n9875 9.3005
R6779 VSS.n9877 VSS.n9876 9.3005
R6780 VSS.n9878 VSS.n9877 9.3005
R6781 VSS.n9866 VSS.n9864 9.3005
R6782 VSS.n9844 VSS.n9355 9.3005
R6783 VSS.n9356 VSS.n9355 9.3005
R6784 VSS.n9858 VSS.n9356 9.3005
R6785 VSS.n9803 VSS.n9802 9.3005
R6786 VSS.n9803 VSS.n9377 9.3005
R6787 VSS.n9807 VSS.n9377 9.3005
R6788 VSS.n9814 VSS.n9374 9.3005
R6789 VSS.n9823 VSS.n9368 9.3005
R6790 VSS.n9368 VSS.n9358 9.3005
R6791 VSS.n9358 VSS.n9357 9.3005
R6792 VSS.n9826 VSS.n9367 9.3005
R6793 VSS.n9841 VSS.n9840 9.3005
R6794 VSS.n9909 VSS.n9908 9.3005
R6795 VSS.n9908 VSS.n9907 9.3005
R6796 VSS.n9756 VSS.n9394 9.3005
R6797 VSS.n9764 VSS.n9763 9.3005
R6798 VSS.n9763 VSS.n9762 9.3005
R6799 VSS.n9387 VSS.n9386 9.3005
R6800 VSS.n9755 VSS.n9386 9.3005
R6801 VSS.n9755 VSS.n9754 9.3005
R6802 VSS.n9793 VSS.n9385 9.3005
R6803 VSS.n9795 VSS.n9794 9.3005
R6804 VSS.n9527 VSS.n9523 9.3005
R6805 VSS.n9505 VSS.n9504 9.3005
R6806 VSS.n9485 VSS.n9484 9.3005
R6807 VSS.n9488 VSS.n9487 9.3005
R6808 VSS.n9615 VSS.n9614 9.3005
R6809 VSS.n9614 VSS.n9613 9.3005
R6810 VSS.n9613 VSS.n9612 9.3005
R6811 VSS.n9570 VSS.n9532 9.3005
R6812 VSS.n9532 VSS.n9531 9.3005
R6813 VSS.n9581 VSS.n9526 9.3005
R6814 VSS.n9581 VSS.n9580 9.3005
R6815 VSS.n9580 VSS.n9579 9.3005
R6816 VSS.n9638 VSS.n9637 9.3005
R6817 VSS.n9639 VSS.n9638 9.3005
R6818 VSS.n9640 VSS.n9639 9.3005
R6819 VSS.n9645 VSS.n9644 9.3005
R6820 VSS.n9644 VSS.n6483 9.3005
R6821 VSS.n9546 VSS.n9543 9.3005
R6822 VSS.n16619 VSS.n16618 9.3005
R6823 VSS.n16657 VSS.n16656 9.3005
R6824 VSS.n16347 VSS.n16346 9.3005
R6825 VSS.n16685 VSS.n16684 9.3005
R6826 VSS.n16664 VSS.n16663 9.3005
R6827 VSS.n16665 VSS.n16664 9.3005
R6828 VSS.n16666 VSS.n16665 9.3005
R6829 VSS.n16632 VSS.n16631 9.3005
R6830 VSS.n16632 VSS.n16381 9.3005
R6831 VSS.n16381 VSS.n16380 9.3005
R6832 VSS.n16612 VSS.n16611 9.3005
R6833 VSS.n16613 VSS.n16612 9.3005
R6834 VSS.n16672 VSS.n16671 9.3005
R6835 VSS.n16671 VSS.n16345 9.3005
R6836 VSS.n16345 VSS.n16344 9.3005
R6837 VSS.n16714 VSS.n16713 9.3005
R6838 VSS.n16713 VSS.n16712 9.3005
R6839 VSS.n16407 VSS.n16405 9.3005
R6840 VSS.n16756 VSS.n16755 9.3005
R6841 VSS.n16271 VSS.n16270 9.3005
R6842 VSS.n16806 VSS.n16296 9.3005
R6843 VSS.n16304 VSS.n16302 9.3005
R6844 VSS.n16771 VSS.n16770 9.3005
R6845 VSS.n16843 VSS.n16842 9.3005
R6846 VSS.n16843 VSS.n16276 9.3005
R6847 VSS.n16276 VSS.n16275 9.3005
R6848 VSS.n16825 VSS.n16284 9.3005
R6849 VSS.n16827 VSS.n16826 9.3005
R6850 VSS.n16819 VSS.n16818 9.3005
R6851 VSS.n16820 VSS.n16819 9.3005
R6852 VSS.n16821 VSS.n16820 9.3005
R6853 VSS.n16809 VSS.n16807 9.3005
R6854 VSS.n16787 VSS.n16297 9.3005
R6855 VSS.n16298 VSS.n16297 9.3005
R6856 VSS.n16801 VSS.n16298 9.3005
R6857 VSS.n16746 VSS.n16745 9.3005
R6858 VSS.n16746 VSS.n16319 9.3005
R6859 VSS.n16750 VSS.n16319 9.3005
R6860 VSS.n16757 VSS.n16316 9.3005
R6861 VSS.n16766 VSS.n16310 9.3005
R6862 VSS.n16310 VSS.n16300 9.3005
R6863 VSS.n16300 VSS.n16299 9.3005
R6864 VSS.n16769 VSS.n16309 9.3005
R6865 VSS.n16784 VSS.n16783 9.3005
R6866 VSS.n16852 VSS.n16851 9.3005
R6867 VSS.n16851 VSS.n16850 9.3005
R6868 VSS.n16699 VSS.n16336 9.3005
R6869 VSS.n16707 VSS.n16706 9.3005
R6870 VSS.n16706 VSS.n16705 9.3005
R6871 VSS.n16329 VSS.n16328 9.3005
R6872 VSS.n16698 VSS.n16328 9.3005
R6873 VSS.n16698 VSS.n16697 9.3005
R6874 VSS.n16736 VSS.n16327 9.3005
R6875 VSS.n16738 VSS.n16737 9.3005
R6876 VSS.n16514 VSS.n16513 9.3005
R6877 VSS.n16552 VSS.n16551 9.3005
R6878 VSS.n16422 VSS.n16421 9.3005
R6879 VSS.n16581 VSS.n16580 9.3005
R6880 VSS.n16559 VSS.n16558 9.3005
R6881 VSS.n16560 VSS.n16559 9.3005
R6882 VSS.n16561 VSS.n16560 9.3005
R6883 VSS.n16527 VSS.n16526 9.3005
R6884 VSS.n16527 VSS.n16458 9.3005
R6885 VSS.n16458 VSS.n16457 9.3005
R6886 VSS.n16507 VSS.n16506 9.3005
R6887 VSS.n16508 VSS.n16507 9.3005
R6888 VSS.n16568 VSS.n16567 9.3005
R6889 VSS.n16567 VSS.n16420 9.3005
R6890 VSS.n16420 VSS.n16419 9.3005
R6891 VSS.n16588 VSS.n16587 9.3005
R6892 VSS.n16587 VSS.n16586 9.3005
R6893 VSS.n16482 VSS.n16480 9.3005
R6894 VSS.n16026 VSS.n16025 9.3005
R6895 VSS.n16064 VSS.n16063 9.3005
R6896 VSS.n1519 VSS.n1518 9.3005
R6897 VSS.n16092 VSS.n16091 9.3005
R6898 VSS.n16071 VSS.n16070 9.3005
R6899 VSS.n16072 VSS.n16071 9.3005
R6900 VSS.n16073 VSS.n16072 9.3005
R6901 VSS.n16039 VSS.n16038 9.3005
R6902 VSS.n16039 VSS.n1553 9.3005
R6903 VSS.n1553 VSS.n1552 9.3005
R6904 VSS.n16019 VSS.n16018 9.3005
R6905 VSS.n16020 VSS.n16019 9.3005
R6906 VSS.n16079 VSS.n16078 9.3005
R6907 VSS.n16078 VSS.n1517 9.3005
R6908 VSS.n1517 VSS.n1516 9.3005
R6909 VSS.n16121 VSS.n16120 9.3005
R6910 VSS.n16120 VSS.n16119 9.3005
R6911 VSS.n1757 VSS.n1756 9.3005
R6912 VSS.n16163 VSS.n16162 9.3005
R6913 VSS.n1443 VSS.n1442 9.3005
R6914 VSS.n16213 VSS.n1468 9.3005
R6915 VSS.n1476 VSS.n1474 9.3005
R6916 VSS.n16178 VSS.n16177 9.3005
R6917 VSS.n16250 VSS.n16249 9.3005
R6918 VSS.n16250 VSS.n1448 9.3005
R6919 VSS.n1448 VSS.n1447 9.3005
R6920 VSS.n16232 VSS.n1456 9.3005
R6921 VSS.n16234 VSS.n16233 9.3005
R6922 VSS.n16226 VSS.n16225 9.3005
R6923 VSS.n16227 VSS.n16226 9.3005
R6924 VSS.n16228 VSS.n16227 9.3005
R6925 VSS.n16216 VSS.n16214 9.3005
R6926 VSS.n16194 VSS.n1469 9.3005
R6927 VSS.n1470 VSS.n1469 9.3005
R6928 VSS.n16208 VSS.n1470 9.3005
R6929 VSS.n16153 VSS.n16152 9.3005
R6930 VSS.n16153 VSS.n1491 9.3005
R6931 VSS.n16157 VSS.n1491 9.3005
R6932 VSS.n16164 VSS.n1488 9.3005
R6933 VSS.n16173 VSS.n1482 9.3005
R6934 VSS.n1482 VSS.n1472 9.3005
R6935 VSS.n1472 VSS.n1471 9.3005
R6936 VSS.n16176 VSS.n1481 9.3005
R6937 VSS.n16191 VSS.n16190 9.3005
R6938 VSS.n16259 VSS.n16258 9.3005
R6939 VSS.n16258 VSS.n16257 9.3005
R6940 VSS.n16106 VSS.n1508 9.3005
R6941 VSS.n16114 VSS.n16113 9.3005
R6942 VSS.n16113 VSS.n16112 9.3005
R6943 VSS.n1501 VSS.n1500 9.3005
R6944 VSS.n16105 VSS.n1500 9.3005
R6945 VSS.n16105 VSS.n16104 9.3005
R6946 VSS.n16143 VSS.n1499 9.3005
R6947 VSS.n16145 VSS.n16144 9.3005
R6948 VSS.n1679 VSS.n1678 9.3005
R6949 VSS.n1717 VSS.n1716 9.3005
R6950 VSS.n1587 VSS.n1586 9.3005
R6951 VSS.n1746 VSS.n1745 9.3005
R6952 VSS.n1724 VSS.n1723 9.3005
R6953 VSS.n1725 VSS.n1724 9.3005
R6954 VSS.n1726 VSS.n1725 9.3005
R6955 VSS.n1692 VSS.n1691 9.3005
R6956 VSS.n1692 VSS.n1623 9.3005
R6957 VSS.n1623 VSS.n1622 9.3005
R6958 VSS.n1672 VSS.n1671 9.3005
R6959 VSS.n1673 VSS.n1672 9.3005
R6960 VSS.n1733 VSS.n1732 9.3005
R6961 VSS.n1732 VSS.n1585 9.3005
R6962 VSS.n1585 VSS.n1584 9.3005
R6963 VSS.n15995 VSS.n15994 9.3005
R6964 VSS.n15994 VSS.n15993 9.3005
R6965 VSS.n1647 VSS.n1645 9.3005
R6966 VSS.n2023 VSS.n2022 9.3005
R6967 VSS.n2044 VSS.n2043 9.3005
R6968 VSS.n1984 VSS.n1983 9.3005
R6969 VSS.n2065 VSS.n2064 9.3005
R6970 VSS.n2050 VSS.n2049 9.3005
R6971 VSS.n2051 VSS.n2050 9.3005
R6972 VSS.n2052 VSS.n2051 9.3005
R6973 VSS.n2031 VSS.n1997 9.3005
R6974 VSS.n2031 VSS.n2030 9.3005
R6975 VSS.n2030 VSS.n2029 9.3005
R6976 VSS.n2016 VSS.n2000 9.3005
R6977 VSS.n2000 VSS.n1999 9.3005
R6978 VSS.n2056 VSS.n1987 9.3005
R6979 VSS.n2056 VSS.n1982 9.3005
R6980 VSS.n1982 VSS.n1981 9.3005
R6981 VSS.n2306 VSS.n2305 9.3005
R6982 VSS.n2305 VSS.n2304 9.3005
R6983 VSS.n2349 VSS.n2348 9.3005
R6984 VSS.n2270 VSS.n2269 9.3005
R6985 VSS.n2225 VSS.n2224 9.3005
R6986 VSS.n2251 VSS.n2250 9.3005
R6987 VSS.n2128 VSS.n2126 9.3005
R6988 VSS.n2146 VSS.n2145 9.3005
R6989 VSS.n2232 VSS.n2172 9.3005
R6990 VSS.n2232 VSS.n2231 9.3005
R6991 VSS.n2231 VSS.n2230 9.3005
R6992 VSS.n2192 VSS.n2163 9.3005
R6993 VSS.n2173 VSS.n2171 9.3005
R6994 VSS.n2162 VSS.n2158 9.3005
R6995 VSS.n2191 VSS.n2158 9.3005
R6996 VSS.n2191 VSS.n2177 9.3005
R6997 VSS.n2249 VSS.n2156 9.3005
R6998 VSS.n2185 VSS.n2184 9.3005
R6999 VSS.n2185 VSS.n2124 9.3005
R7000 VSS.n2124 VSS.n2123 9.3005
R7001 VSS.n2277 VSS.n2276 9.3005
R7002 VSS.n2278 VSS.n2277 9.3005
R7003 VSS.n2279 VSS.n2278 9.3005
R7004 VSS.n2271 VSS.n2119 9.3005
R7005 VSS.n2141 VSS.n2121 9.3005
R7006 VSS.n2122 VSS.n2121 9.3005
R7007 VSS.n2264 VSS.n2122 9.3005
R7008 VSS.n2144 VSS.n2133 9.3005
R7009 VSS.n2180 VSS.n2179 9.3005
R7010 VSS.n2206 VSS.n2198 9.3005
R7011 VSS.n2198 VSS.n2197 9.3005
R7012 VSS.n2087 VSS.n2086 9.3005
R7013 VSS.n2299 VSS.n2298 9.3005
R7014 VSS.n2298 VSS.n2297 9.3005
R7015 VSS.n2292 VSS.n2291 9.3005
R7016 VSS.n2292 VSS.n2076 9.3005
R7017 VSS.n2076 VSS.n2075 9.3005
R7018 VSS.n2286 VSS.n2285 9.3005
R7019 VSS.n2284 VSS.n2102 9.3005
R7020 VSS.n1819 VSS.n1815 9.3005
R7021 VSS.n1797 VSS.n1796 9.3005
R7022 VSS.n1777 VSS.n1776 9.3005
R7023 VSS.n1780 VSS.n1779 9.3005
R7024 VSS.n1907 VSS.n1906 9.3005
R7025 VSS.n1906 VSS.n1905 9.3005
R7026 VSS.n1905 VSS.n1904 9.3005
R7027 VSS.n1873 VSS.n1818 9.3005
R7028 VSS.n1873 VSS.n1872 9.3005
R7029 VSS.n1872 VSS.n1871 9.3005
R7030 VSS.n1862 VSS.n1824 9.3005
R7031 VSS.n1824 VSS.n1823 9.3005
R7032 VSS.n1930 VSS.n1929 9.3005
R7033 VSS.n1931 VSS.n1930 9.3005
R7034 VSS.n1932 VSS.n1931 9.3005
R7035 VSS.n1937 VSS.n1936 9.3005
R7036 VSS.n1936 VSS.n1758 9.3005
R7037 VSS.n1838 VSS.n1835 9.3005
R7038 VSS.n3167 VSS.n3166 9.3005
R7039 VSS.n3205 VSS.n3204 9.3005
R7040 VSS.n2896 VSS.n2895 9.3005
R7041 VSS.n3233 VSS.n3232 9.3005
R7042 VSS.n3212 VSS.n3211 9.3005
R7043 VSS.n3213 VSS.n3212 9.3005
R7044 VSS.n3214 VSS.n3213 9.3005
R7045 VSS.n3180 VSS.n3179 9.3005
R7046 VSS.n3180 VSS.n2930 9.3005
R7047 VSS.n2930 VSS.n2929 9.3005
R7048 VSS.n3160 VSS.n3159 9.3005
R7049 VSS.n3161 VSS.n3160 9.3005
R7050 VSS.n3220 VSS.n3219 9.3005
R7051 VSS.n3219 VSS.n2894 9.3005
R7052 VSS.n2894 VSS.n2893 9.3005
R7053 VSS.n3262 VSS.n3261 9.3005
R7054 VSS.n3261 VSS.n3260 9.3005
R7055 VSS.n2956 VSS.n2954 9.3005
R7056 VSS.n3304 VSS.n3303 9.3005
R7057 VSS.n2820 VSS.n2819 9.3005
R7058 VSS.n3354 VSS.n2845 9.3005
R7059 VSS.n2853 VSS.n2851 9.3005
R7060 VSS.n3319 VSS.n3318 9.3005
R7061 VSS.n3391 VSS.n3390 9.3005
R7062 VSS.n3391 VSS.n2825 9.3005
R7063 VSS.n2825 VSS.n2824 9.3005
R7064 VSS.n3373 VSS.n2833 9.3005
R7065 VSS.n3375 VSS.n3374 9.3005
R7066 VSS.n3367 VSS.n3366 9.3005
R7067 VSS.n3368 VSS.n3367 9.3005
R7068 VSS.n3369 VSS.n3368 9.3005
R7069 VSS.n3357 VSS.n3355 9.3005
R7070 VSS.n3335 VSS.n2846 9.3005
R7071 VSS.n2847 VSS.n2846 9.3005
R7072 VSS.n3349 VSS.n2847 9.3005
R7073 VSS.n3294 VSS.n3293 9.3005
R7074 VSS.n3294 VSS.n2868 9.3005
R7075 VSS.n3298 VSS.n2868 9.3005
R7076 VSS.n3305 VSS.n2865 9.3005
R7077 VSS.n3314 VSS.n2859 9.3005
R7078 VSS.n2859 VSS.n2849 9.3005
R7079 VSS.n2849 VSS.n2848 9.3005
R7080 VSS.n3317 VSS.n2858 9.3005
R7081 VSS.n3332 VSS.n3331 9.3005
R7082 VSS.n3400 VSS.n3399 9.3005
R7083 VSS.n3399 VSS.n3398 9.3005
R7084 VSS.n3247 VSS.n2885 9.3005
R7085 VSS.n3255 VSS.n3254 9.3005
R7086 VSS.n3254 VSS.n3253 9.3005
R7087 VSS.n2878 VSS.n2877 9.3005
R7088 VSS.n3246 VSS.n2877 9.3005
R7089 VSS.n3246 VSS.n3245 9.3005
R7090 VSS.n3284 VSS.n2876 9.3005
R7091 VSS.n3286 VSS.n3285 9.3005
R7092 VSS.n3018 VSS.n3014 9.3005
R7093 VSS.n2996 VSS.n2995 9.3005
R7094 VSS.n2976 VSS.n2975 9.3005
R7095 VSS.n2979 VSS.n2978 9.3005
R7096 VSS.n3106 VSS.n3105 9.3005
R7097 VSS.n3105 VSS.n3104 9.3005
R7098 VSS.n3104 VSS.n3103 9.3005
R7099 VSS.n3072 VSS.n3017 9.3005
R7100 VSS.n3072 VSS.n3071 9.3005
R7101 VSS.n3071 VSS.n3070 9.3005
R7102 VSS.n3061 VSS.n3023 9.3005
R7103 VSS.n3023 VSS.n3022 9.3005
R7104 VSS.n3129 VSS.n3128 9.3005
R7105 VSS.n3130 VSS.n3129 9.3005
R7106 VSS.n3131 VSS.n3130 9.3005
R7107 VSS.n3136 VSS.n3135 9.3005
R7108 VSS.n3135 VSS.n2350 9.3005
R7109 VSS.n3037 VSS.n3034 9.3005
R7110 VSS.n3759 VSS.n3758 9.3005
R7111 VSS.n3797 VSS.n3796 9.3005
R7112 VSS.n3488 VSS.n3487 9.3005
R7113 VSS.n3825 VSS.n3824 9.3005
R7114 VSS.n3804 VSS.n3803 9.3005
R7115 VSS.n3805 VSS.n3804 9.3005
R7116 VSS.n3806 VSS.n3805 9.3005
R7117 VSS.n3772 VSS.n3771 9.3005
R7118 VSS.n3772 VSS.n3522 9.3005
R7119 VSS.n3522 VSS.n3521 9.3005
R7120 VSS.n3752 VSS.n3751 9.3005
R7121 VSS.n3753 VSS.n3752 9.3005
R7122 VSS.n3812 VSS.n3811 9.3005
R7123 VSS.n3811 VSS.n3486 9.3005
R7124 VSS.n3486 VSS.n3485 9.3005
R7125 VSS.n3854 VSS.n3853 9.3005
R7126 VSS.n3853 VSS.n3852 9.3005
R7127 VSS.n3548 VSS.n3546 9.3005
R7128 VSS.n3896 VSS.n3895 9.3005
R7129 VSS.n3412 VSS.n3411 9.3005
R7130 VSS.n3946 VSS.n3437 9.3005
R7131 VSS.n3445 VSS.n3443 9.3005
R7132 VSS.n3911 VSS.n3910 9.3005
R7133 VSS.n3983 VSS.n3982 9.3005
R7134 VSS.n3983 VSS.n3417 9.3005
R7135 VSS.n3417 VSS.n3416 9.3005
R7136 VSS.n3965 VSS.n3425 9.3005
R7137 VSS.n3967 VSS.n3966 9.3005
R7138 VSS.n3959 VSS.n3958 9.3005
R7139 VSS.n3960 VSS.n3959 9.3005
R7140 VSS.n3961 VSS.n3960 9.3005
R7141 VSS.n3949 VSS.n3947 9.3005
R7142 VSS.n3927 VSS.n3438 9.3005
R7143 VSS.n3439 VSS.n3438 9.3005
R7144 VSS.n3941 VSS.n3439 9.3005
R7145 VSS.n3886 VSS.n3885 9.3005
R7146 VSS.n3886 VSS.n3460 9.3005
R7147 VSS.n3890 VSS.n3460 9.3005
R7148 VSS.n3897 VSS.n3457 9.3005
R7149 VSS.n3906 VSS.n3451 9.3005
R7150 VSS.n3451 VSS.n3441 9.3005
R7151 VSS.n3441 VSS.n3440 9.3005
R7152 VSS.n3909 VSS.n3450 9.3005
R7153 VSS.n3924 VSS.n3923 9.3005
R7154 VSS.n3992 VSS.n3991 9.3005
R7155 VSS.n3991 VSS.n3990 9.3005
R7156 VSS.n3839 VSS.n3477 9.3005
R7157 VSS.n3847 VSS.n3846 9.3005
R7158 VSS.n3846 VSS.n3845 9.3005
R7159 VSS.n3470 VSS.n3469 9.3005
R7160 VSS.n3838 VSS.n3469 9.3005
R7161 VSS.n3838 VSS.n3837 9.3005
R7162 VSS.n3876 VSS.n3468 9.3005
R7163 VSS.n3878 VSS.n3877 9.3005
R7164 VSS.n3610 VSS.n3606 9.3005
R7165 VSS.n3588 VSS.n3587 9.3005
R7166 VSS.n3568 VSS.n3567 9.3005
R7167 VSS.n3571 VSS.n3570 9.3005
R7168 VSS.n3698 VSS.n3697 9.3005
R7169 VSS.n3697 VSS.n3696 9.3005
R7170 VSS.n3696 VSS.n3695 9.3005
R7171 VSS.n3664 VSS.n3609 9.3005
R7172 VSS.n3664 VSS.n3663 9.3005
R7173 VSS.n3663 VSS.n3662 9.3005
R7174 VSS.n3653 VSS.n3615 9.3005
R7175 VSS.n3615 VSS.n3614 9.3005
R7176 VSS.n3721 VSS.n3720 9.3005
R7177 VSS.n3722 VSS.n3721 9.3005
R7178 VSS.n3723 VSS.n3722 9.3005
R7179 VSS.n3728 VSS.n3727 9.3005
R7180 VSS.n3727 VSS.n2351 9.3005
R7181 VSS.n3629 VSS.n3626 9.3005
R7182 VSS.n4351 VSS.n4350 9.3005
R7183 VSS.n4389 VSS.n4388 9.3005
R7184 VSS.n4080 VSS.n4079 9.3005
R7185 VSS.n4417 VSS.n4416 9.3005
R7186 VSS.n4396 VSS.n4395 9.3005
R7187 VSS.n4397 VSS.n4396 9.3005
R7188 VSS.n4398 VSS.n4397 9.3005
R7189 VSS.n4364 VSS.n4363 9.3005
R7190 VSS.n4364 VSS.n4114 9.3005
R7191 VSS.n4114 VSS.n4113 9.3005
R7192 VSS.n4344 VSS.n4343 9.3005
R7193 VSS.n4345 VSS.n4344 9.3005
R7194 VSS.n4404 VSS.n4403 9.3005
R7195 VSS.n4403 VSS.n4078 9.3005
R7196 VSS.n4078 VSS.n4077 9.3005
R7197 VSS.n4446 VSS.n4445 9.3005
R7198 VSS.n4445 VSS.n4444 9.3005
R7199 VSS.n4140 VSS.n4138 9.3005
R7200 VSS.n4488 VSS.n4487 9.3005
R7201 VSS.n4004 VSS.n4003 9.3005
R7202 VSS.n4538 VSS.n4029 9.3005
R7203 VSS.n4037 VSS.n4035 9.3005
R7204 VSS.n4503 VSS.n4502 9.3005
R7205 VSS.n4575 VSS.n4574 9.3005
R7206 VSS.n4575 VSS.n4009 9.3005
R7207 VSS.n4009 VSS.n4008 9.3005
R7208 VSS.n4557 VSS.n4017 9.3005
R7209 VSS.n4559 VSS.n4558 9.3005
R7210 VSS.n4551 VSS.n4550 9.3005
R7211 VSS.n4552 VSS.n4551 9.3005
R7212 VSS.n4553 VSS.n4552 9.3005
R7213 VSS.n4541 VSS.n4539 9.3005
R7214 VSS.n4519 VSS.n4030 9.3005
R7215 VSS.n4031 VSS.n4030 9.3005
R7216 VSS.n4533 VSS.n4031 9.3005
R7217 VSS.n4478 VSS.n4477 9.3005
R7218 VSS.n4478 VSS.n4052 9.3005
R7219 VSS.n4482 VSS.n4052 9.3005
R7220 VSS.n4489 VSS.n4049 9.3005
R7221 VSS.n4498 VSS.n4043 9.3005
R7222 VSS.n4043 VSS.n4033 9.3005
R7223 VSS.n4033 VSS.n4032 9.3005
R7224 VSS.n4501 VSS.n4042 9.3005
R7225 VSS.n4516 VSS.n4515 9.3005
R7226 VSS.n4584 VSS.n4583 9.3005
R7227 VSS.n4583 VSS.n4582 9.3005
R7228 VSS.n4431 VSS.n4069 9.3005
R7229 VSS.n4439 VSS.n4438 9.3005
R7230 VSS.n4438 VSS.n4437 9.3005
R7231 VSS.n4062 VSS.n4061 9.3005
R7232 VSS.n4430 VSS.n4061 9.3005
R7233 VSS.n4430 VSS.n4429 9.3005
R7234 VSS.n4468 VSS.n4060 9.3005
R7235 VSS.n4470 VSS.n4469 9.3005
R7236 VSS.n4202 VSS.n4198 9.3005
R7237 VSS.n4180 VSS.n4179 9.3005
R7238 VSS.n4160 VSS.n4159 9.3005
R7239 VSS.n4163 VSS.n4162 9.3005
R7240 VSS.n4290 VSS.n4289 9.3005
R7241 VSS.n4289 VSS.n4288 9.3005
R7242 VSS.n4288 VSS.n4287 9.3005
R7243 VSS.n4256 VSS.n4201 9.3005
R7244 VSS.n4256 VSS.n4255 9.3005
R7245 VSS.n4255 VSS.n4254 9.3005
R7246 VSS.n4245 VSS.n4207 9.3005
R7247 VSS.n4207 VSS.n4206 9.3005
R7248 VSS.n4313 VSS.n4312 9.3005
R7249 VSS.n4314 VSS.n4313 9.3005
R7250 VSS.n4315 VSS.n4314 9.3005
R7251 VSS.n4320 VSS.n4319 9.3005
R7252 VSS.n4319 VSS.n2352 9.3005
R7253 VSS.n4221 VSS.n4218 9.3005
R7254 VSS.n4943 VSS.n4942 9.3005
R7255 VSS.n4981 VSS.n4980 9.3005
R7256 VSS.n4672 VSS.n4671 9.3005
R7257 VSS.n5009 VSS.n5008 9.3005
R7258 VSS.n4988 VSS.n4987 9.3005
R7259 VSS.n4989 VSS.n4988 9.3005
R7260 VSS.n4990 VSS.n4989 9.3005
R7261 VSS.n4956 VSS.n4955 9.3005
R7262 VSS.n4956 VSS.n4706 9.3005
R7263 VSS.n4706 VSS.n4705 9.3005
R7264 VSS.n4936 VSS.n4935 9.3005
R7265 VSS.n4937 VSS.n4936 9.3005
R7266 VSS.n4996 VSS.n4995 9.3005
R7267 VSS.n4995 VSS.n4670 9.3005
R7268 VSS.n4670 VSS.n4669 9.3005
R7269 VSS.n5038 VSS.n5037 9.3005
R7270 VSS.n5037 VSS.n5036 9.3005
R7271 VSS.n4732 VSS.n4730 9.3005
R7272 VSS.n5080 VSS.n5079 9.3005
R7273 VSS.n4596 VSS.n4595 9.3005
R7274 VSS.n5130 VSS.n4621 9.3005
R7275 VSS.n4629 VSS.n4627 9.3005
R7276 VSS.n5095 VSS.n5094 9.3005
R7277 VSS.n5167 VSS.n5166 9.3005
R7278 VSS.n5167 VSS.n4601 9.3005
R7279 VSS.n4601 VSS.n4600 9.3005
R7280 VSS.n5149 VSS.n4609 9.3005
R7281 VSS.n5151 VSS.n5150 9.3005
R7282 VSS.n5143 VSS.n5142 9.3005
R7283 VSS.n5144 VSS.n5143 9.3005
R7284 VSS.n5145 VSS.n5144 9.3005
R7285 VSS.n5133 VSS.n5131 9.3005
R7286 VSS.n5111 VSS.n4622 9.3005
R7287 VSS.n4623 VSS.n4622 9.3005
R7288 VSS.n5125 VSS.n4623 9.3005
R7289 VSS.n5070 VSS.n5069 9.3005
R7290 VSS.n5070 VSS.n4644 9.3005
R7291 VSS.n5074 VSS.n4644 9.3005
R7292 VSS.n5081 VSS.n4641 9.3005
R7293 VSS.n5090 VSS.n4635 9.3005
R7294 VSS.n4635 VSS.n4625 9.3005
R7295 VSS.n4625 VSS.n4624 9.3005
R7296 VSS.n5093 VSS.n4634 9.3005
R7297 VSS.n5108 VSS.n5107 9.3005
R7298 VSS.n5176 VSS.n5175 9.3005
R7299 VSS.n5175 VSS.n5174 9.3005
R7300 VSS.n5023 VSS.n4661 9.3005
R7301 VSS.n5031 VSS.n5030 9.3005
R7302 VSS.n5030 VSS.n5029 9.3005
R7303 VSS.n4654 VSS.n4653 9.3005
R7304 VSS.n5022 VSS.n4653 9.3005
R7305 VSS.n5022 VSS.n5021 9.3005
R7306 VSS.n5060 VSS.n4652 9.3005
R7307 VSS.n5062 VSS.n5061 9.3005
R7308 VSS.n4794 VSS.n4790 9.3005
R7309 VSS.n4772 VSS.n4771 9.3005
R7310 VSS.n4752 VSS.n4751 9.3005
R7311 VSS.n4755 VSS.n4754 9.3005
R7312 VSS.n4882 VSS.n4881 9.3005
R7313 VSS.n4881 VSS.n4880 9.3005
R7314 VSS.n4880 VSS.n4879 9.3005
R7315 VSS.n4848 VSS.n4793 9.3005
R7316 VSS.n4848 VSS.n4847 9.3005
R7317 VSS.n4847 VSS.n4846 9.3005
R7318 VSS.n4837 VSS.n4799 9.3005
R7319 VSS.n4799 VSS.n4798 9.3005
R7320 VSS.n4905 VSS.n4904 9.3005
R7321 VSS.n4906 VSS.n4905 9.3005
R7322 VSS.n4907 VSS.n4906 9.3005
R7323 VSS.n4912 VSS.n4911 9.3005
R7324 VSS.n4911 VSS.n2353 9.3005
R7325 VSS.n4813 VSS.n4810 9.3005
R7326 VSS.n2619 VSS.n2618 9.3005
R7327 VSS.n2640 VSS.n2639 9.3005
R7328 VSS.n2580 VSS.n2579 9.3005
R7329 VSS.n2661 VSS.n2660 9.3005
R7330 VSS.n2646 VSS.n2645 9.3005
R7331 VSS.n2647 VSS.n2646 9.3005
R7332 VSS.n2648 VSS.n2647 9.3005
R7333 VSS.n2627 VSS.n2593 9.3005
R7334 VSS.n2627 VSS.n2626 9.3005
R7335 VSS.n2626 VSS.n2625 9.3005
R7336 VSS.n2612 VSS.n2596 9.3005
R7337 VSS.n2596 VSS.n2595 9.3005
R7338 VSS.n2652 VSS.n2583 9.3005
R7339 VSS.n2652 VSS.n2578 9.3005
R7340 VSS.n2578 VSS.n2577 9.3005
R7341 VSS.n5271 VSS.n5270 9.3005
R7342 VSS.n5270 VSS.n5269 9.3005
R7343 VSS.n5314 VSS.n5313 9.3005
R7344 VSS.n5235 VSS.n5234 9.3005
R7345 VSS.n5190 VSS.n5189 9.3005
R7346 VSS.n5216 VSS.n5215 9.3005
R7347 VSS.n2724 VSS.n2722 9.3005
R7348 VSS.n2742 VSS.n2741 9.3005
R7349 VSS.n5197 VSS.n2768 9.3005
R7350 VSS.n5197 VSS.n5196 9.3005
R7351 VSS.n5196 VSS.n5195 9.3005
R7352 VSS.n2788 VSS.n2759 9.3005
R7353 VSS.n2769 VSS.n2767 9.3005
R7354 VSS.n2758 VSS.n2754 9.3005
R7355 VSS.n2787 VSS.n2754 9.3005
R7356 VSS.n2787 VSS.n2773 9.3005
R7357 VSS.n5214 VSS.n2752 9.3005
R7358 VSS.n2781 VSS.n2780 9.3005
R7359 VSS.n2781 VSS.n2720 9.3005
R7360 VSS.n2720 VSS.n2719 9.3005
R7361 VSS.n5242 VSS.n5241 9.3005
R7362 VSS.n5243 VSS.n5242 9.3005
R7363 VSS.n5244 VSS.n5243 9.3005
R7364 VSS.n5236 VSS.n2715 9.3005
R7365 VSS.n2737 VSS.n2717 9.3005
R7366 VSS.n2718 VSS.n2717 9.3005
R7367 VSS.n5229 VSS.n2718 9.3005
R7368 VSS.n2740 VSS.n2729 9.3005
R7369 VSS.n2776 VSS.n2775 9.3005
R7370 VSS.n2802 VSS.n2794 9.3005
R7371 VSS.n2794 VSS.n2793 9.3005
R7372 VSS.n2683 VSS.n2682 9.3005
R7373 VSS.n5264 VSS.n5263 9.3005
R7374 VSS.n5263 VSS.n5262 9.3005
R7375 VSS.n5257 VSS.n5256 9.3005
R7376 VSS.n5257 VSS.n2672 9.3005
R7377 VSS.n2672 VSS.n2671 9.3005
R7378 VSS.n5251 VSS.n5250 9.3005
R7379 VSS.n5249 VSS.n2698 9.3005
R7380 VSS.n2415 VSS.n2411 9.3005
R7381 VSS.n2393 VSS.n2392 9.3005
R7382 VSS.n2373 VSS.n2372 9.3005
R7383 VSS.n2376 VSS.n2375 9.3005
R7384 VSS.n2503 VSS.n2502 9.3005
R7385 VSS.n2502 VSS.n2501 9.3005
R7386 VSS.n2501 VSS.n2500 9.3005
R7387 VSS.n2469 VSS.n2414 9.3005
R7388 VSS.n2469 VSS.n2468 9.3005
R7389 VSS.n2468 VSS.n2467 9.3005
R7390 VSS.n2458 VSS.n2420 9.3005
R7391 VSS.n2420 VSS.n2419 9.3005
R7392 VSS.n2526 VSS.n2525 9.3005
R7393 VSS.n2527 VSS.n2526 9.3005
R7394 VSS.n2528 VSS.n2527 9.3005
R7395 VSS.n2533 VSS.n2532 9.3005
R7396 VSS.n2532 VSS.n2354 9.3005
R7397 VSS.n2434 VSS.n2431 9.3005
R7398 VSS.n5580 VSS.n5579 9.3005
R7399 VSS.n5601 VSS.n5600 9.3005
R7400 VSS.n5541 VSS.n5540 9.3005
R7401 VSS.n5622 VSS.n5621 9.3005
R7402 VSS.n5607 VSS.n5606 9.3005
R7403 VSS.n5608 VSS.n5607 9.3005
R7404 VSS.n5609 VSS.n5608 9.3005
R7405 VSS.n5588 VSS.n5554 9.3005
R7406 VSS.n5588 VSS.n5587 9.3005
R7407 VSS.n5587 VSS.n5586 9.3005
R7408 VSS.n5573 VSS.n5557 9.3005
R7409 VSS.n5557 VSS.n5556 9.3005
R7410 VSS.n5613 VSS.n5544 9.3005
R7411 VSS.n5613 VSS.n5539 9.3005
R7412 VSS.n5539 VSS.n5538 9.3005
R7413 VSS.n5844 VSS.n5843 9.3005
R7414 VSS.n5843 VSS.n5842 9.3005
R7415 VSS.n5887 VSS.n5886 9.3005
R7416 VSS.n5808 VSS.n5807 9.3005
R7417 VSS.n5 VSS.n4 9.3005
R7418 VSS.n5789 VSS.n5788 9.3005
R7419 VSS.n5685 VSS.n5683 9.3005
R7420 VSS.n5703 VSS.n5702 9.3005
R7421 VSS.n5770 VSS.n5741 9.3005
R7422 VSS.n5770 VSS.n5769 9.3005
R7423 VSS.n5769 VSS.n5768 9.3005
R7424 VSS.n5762 VSS.n5720 9.3005
R7425 VSS.n5742 VSS.n5728 9.3005
R7426 VSS.n5719 VSS.n5715 9.3005
R7427 VSS.n5761 VSS.n5715 9.3005
R7428 VSS.n5761 VSS.n5747 9.3005
R7429 VSS.n5787 VSS.n5713 9.3005
R7430 VSS.n5755 VSS.n5754 9.3005
R7431 VSS.n5755 VSS.n5681 9.3005
R7432 VSS.n5681 VSS.n5680 9.3005
R7433 VSS.n5815 VSS.n5814 9.3005
R7434 VSS.n5816 VSS.n5815 9.3005
R7435 VSS.n5817 VSS.n5816 9.3005
R7436 VSS.n5809 VSS.n5676 9.3005
R7437 VSS.n5698 VSS.n5678 9.3005
R7438 VSS.n5679 VSS.n5678 9.3005
R7439 VSS.n5802 VSS.n5679 9.3005
R7440 VSS.n5701 VSS.n5690 9.3005
R7441 VSS.n5750 VSS.n5749 9.3005
R7442 VSS.n18882 VSS.n18881 9.3005
R7443 VSS.n18881 VSS.n18880 9.3005
R7444 VSS.n5644 VSS.n5643 9.3005
R7445 VSS.n5837 VSS.n5836 9.3005
R7446 VSS.n5836 VSS.n5835 9.3005
R7447 VSS.n5830 VSS.n5829 9.3005
R7448 VSS.n5830 VSS.n5633 9.3005
R7449 VSS.n5633 VSS.n5632 9.3005
R7450 VSS.n5824 VSS.n5823 9.3005
R7451 VSS.n5822 VSS.n5659 9.3005
R7452 VSS.n5376 VSS.n5372 9.3005
R7453 VSS.n5354 VSS.n5353 9.3005
R7454 VSS.n5334 VSS.n5333 9.3005
R7455 VSS.n5337 VSS.n5336 9.3005
R7456 VSS.n5464 VSS.n5463 9.3005
R7457 VSS.n5463 VSS.n5462 9.3005
R7458 VSS.n5462 VSS.n5461 9.3005
R7459 VSS.n5430 VSS.n5375 9.3005
R7460 VSS.n5430 VSS.n5429 9.3005
R7461 VSS.n5429 VSS.n5428 9.3005
R7462 VSS.n5419 VSS.n5381 9.3005
R7463 VSS.n5381 VSS.n5380 9.3005
R7464 VSS.n5487 VSS.n5486 9.3005
R7465 VSS.n5488 VSS.n5487 9.3005
R7466 VSS.n5489 VSS.n5488 9.3005
R7467 VSS.n5494 VSS.n5493 9.3005
R7468 VSS.n5493 VSS.n5315 9.3005
R7469 VSS.n5395 VSS.n5392 9.3005
R7470 VSS.n6153 VSS.n6152 9.3005
R7471 VSS.n6174 VSS.n6173 9.3005
R7472 VSS.n6114 VSS.n6113 9.3005
R7473 VSS.n6195 VSS.n6194 9.3005
R7474 VSS.n6180 VSS.n6179 9.3005
R7475 VSS.n6181 VSS.n6180 9.3005
R7476 VSS.n6182 VSS.n6181 9.3005
R7477 VSS.n6161 VSS.n6127 9.3005
R7478 VSS.n6161 VSS.n6160 9.3005
R7479 VSS.n6160 VSS.n6159 9.3005
R7480 VSS.n6146 VSS.n6130 9.3005
R7481 VSS.n6130 VSS.n6129 9.3005
R7482 VSS.n6186 VSS.n6117 9.3005
R7483 VSS.n6186 VSS.n6112 9.3005
R7484 VSS.n6112 VSS.n6111 9.3005
R7485 VSS.n6436 VSS.n6435 9.3005
R7486 VSS.n6435 VSS.n6434 9.3005
R7487 VSS.n6479 VSS.n6478 9.3005
R7488 VSS.n6400 VSS.n6399 9.3005
R7489 VSS.n6355 VSS.n6354 9.3005
R7490 VSS.n6381 VSS.n6380 9.3005
R7491 VSS.n6258 VSS.n6256 9.3005
R7492 VSS.n6276 VSS.n6275 9.3005
R7493 VSS.n6362 VSS.n6302 9.3005
R7494 VSS.n6362 VSS.n6361 9.3005
R7495 VSS.n6361 VSS.n6360 9.3005
R7496 VSS.n6322 VSS.n6293 9.3005
R7497 VSS.n6303 VSS.n6301 9.3005
R7498 VSS.n6292 VSS.n6288 9.3005
R7499 VSS.n6321 VSS.n6288 9.3005
R7500 VSS.n6321 VSS.n6307 9.3005
R7501 VSS.n6379 VSS.n6286 9.3005
R7502 VSS.n6315 VSS.n6314 9.3005
R7503 VSS.n6315 VSS.n6254 9.3005
R7504 VSS.n6254 VSS.n6253 9.3005
R7505 VSS.n6407 VSS.n6406 9.3005
R7506 VSS.n6408 VSS.n6407 9.3005
R7507 VSS.n6409 VSS.n6408 9.3005
R7508 VSS.n6401 VSS.n6249 9.3005
R7509 VSS.n6271 VSS.n6251 9.3005
R7510 VSS.n6252 VSS.n6251 9.3005
R7511 VSS.n6394 VSS.n6252 9.3005
R7512 VSS.n6274 VSS.n6263 9.3005
R7513 VSS.n6310 VSS.n6309 9.3005
R7514 VSS.n6336 VSS.n6328 9.3005
R7515 VSS.n6328 VSS.n6327 9.3005
R7516 VSS.n6217 VSS.n6216 9.3005
R7517 VSS.n6429 VSS.n6428 9.3005
R7518 VSS.n6428 VSS.n6427 9.3005
R7519 VSS.n6422 VSS.n6421 9.3005
R7520 VSS.n6422 VSS.n6206 9.3005
R7521 VSS.n6206 VSS.n6205 9.3005
R7522 VSS.n6416 VSS.n6415 9.3005
R7523 VSS.n6414 VSS.n6232 9.3005
R7524 VSS.n5949 VSS.n5945 9.3005
R7525 VSS.n5927 VSS.n5926 9.3005
R7526 VSS.n5907 VSS.n5906 9.3005
R7527 VSS.n5910 VSS.n5909 9.3005
R7528 VSS.n6037 VSS.n6036 9.3005
R7529 VSS.n6036 VSS.n6035 9.3005
R7530 VSS.n6035 VSS.n6034 9.3005
R7531 VSS.n6003 VSS.n5948 9.3005
R7532 VSS.n6003 VSS.n6002 9.3005
R7533 VSS.n6002 VSS.n6001 9.3005
R7534 VSS.n5992 VSS.n5954 9.3005
R7535 VSS.n5954 VSS.n5953 9.3005
R7536 VSS.n6060 VSS.n6059 9.3005
R7537 VSS.n6061 VSS.n6060 9.3005
R7538 VSS.n6062 VSS.n6061 9.3005
R7539 VSS.n6067 VSS.n6066 9.3005
R7540 VSS.n6066 VSS.n5888 9.3005
R7541 VSS.n5968 VSS.n5965 9.3005
R7542 VSS.n7900 VSS.n7899 9.3005
R7543 VSS.n7938 VSS.n7937 9.3005
R7544 VSS.n7629 VSS.n7628 9.3005
R7545 VSS.n7966 VSS.n7965 9.3005
R7546 VSS.n7945 VSS.n7944 9.3005
R7547 VSS.n7946 VSS.n7945 9.3005
R7548 VSS.n7947 VSS.n7946 9.3005
R7549 VSS.n7913 VSS.n7912 9.3005
R7550 VSS.n7913 VSS.n7663 9.3005
R7551 VSS.n7663 VSS.n7662 9.3005
R7552 VSS.n7893 VSS.n7892 9.3005
R7553 VSS.n7894 VSS.n7893 9.3005
R7554 VSS.n7953 VSS.n7952 9.3005
R7555 VSS.n7952 VSS.n7627 9.3005
R7556 VSS.n7627 VSS.n7626 9.3005
R7557 VSS.n7995 VSS.n7994 9.3005
R7558 VSS.n7994 VSS.n7993 9.3005
R7559 VSS.n7689 VSS.n7687 9.3005
R7560 VSS.n8037 VSS.n8036 9.3005
R7561 VSS.n7553 VSS.n7552 9.3005
R7562 VSS.n8087 VSS.n7578 9.3005
R7563 VSS.n7586 VSS.n7584 9.3005
R7564 VSS.n8052 VSS.n8051 9.3005
R7565 VSS.n8124 VSS.n8123 9.3005
R7566 VSS.n8124 VSS.n7558 9.3005
R7567 VSS.n7558 VSS.n7557 9.3005
R7568 VSS.n8106 VSS.n7566 9.3005
R7569 VSS.n8108 VSS.n8107 9.3005
R7570 VSS.n8100 VSS.n8099 9.3005
R7571 VSS.n8101 VSS.n8100 9.3005
R7572 VSS.n8102 VSS.n8101 9.3005
R7573 VSS.n8090 VSS.n8088 9.3005
R7574 VSS.n8068 VSS.n7579 9.3005
R7575 VSS.n7580 VSS.n7579 9.3005
R7576 VSS.n8082 VSS.n7580 9.3005
R7577 VSS.n8027 VSS.n8026 9.3005
R7578 VSS.n8027 VSS.n7601 9.3005
R7579 VSS.n8031 VSS.n7601 9.3005
R7580 VSS.n8038 VSS.n7598 9.3005
R7581 VSS.n8047 VSS.n7592 9.3005
R7582 VSS.n7592 VSS.n7582 9.3005
R7583 VSS.n7582 VSS.n7581 9.3005
R7584 VSS.n8050 VSS.n7591 9.3005
R7585 VSS.n8065 VSS.n8064 9.3005
R7586 VSS.n8133 VSS.n8132 9.3005
R7587 VSS.n8132 VSS.n8131 9.3005
R7588 VSS.n7980 VSS.n7618 9.3005
R7589 VSS.n7988 VSS.n7987 9.3005
R7590 VSS.n7987 VSS.n7986 9.3005
R7591 VSS.n7611 VSS.n7610 9.3005
R7592 VSS.n7979 VSS.n7610 9.3005
R7593 VSS.n7979 VSS.n7978 9.3005
R7594 VSS.n8017 VSS.n7609 9.3005
R7595 VSS.n8019 VSS.n8018 9.3005
R7596 VSS.n7751 VSS.n7747 9.3005
R7597 VSS.n7729 VSS.n7728 9.3005
R7598 VSS.n7709 VSS.n7708 9.3005
R7599 VSS.n7712 VSS.n7711 9.3005
R7600 VSS.n7839 VSS.n7838 9.3005
R7601 VSS.n7838 VSS.n7837 9.3005
R7602 VSS.n7837 VSS.n7836 9.3005
R7603 VSS.n7805 VSS.n7750 9.3005
R7604 VSS.n7805 VSS.n7804 9.3005
R7605 VSS.n7804 VSS.n7803 9.3005
R7606 VSS.n7794 VSS.n7756 9.3005
R7607 VSS.n7756 VSS.n7755 9.3005
R7608 VSS.n7862 VSS.n7861 9.3005
R7609 VSS.n7863 VSS.n7862 9.3005
R7610 VSS.n7864 VSS.n7863 9.3005
R7611 VSS.n7869 VSS.n7868 9.3005
R7612 VSS.n7868 VSS.n6480 9.3005
R7613 VSS.n7770 VSS.n7767 9.3005
R7614 VSS.n8492 VSS.n8491 9.3005
R7615 VSS.n8530 VSS.n8529 9.3005
R7616 VSS.n8221 VSS.n8220 9.3005
R7617 VSS.n8558 VSS.n8557 9.3005
R7618 VSS.n8537 VSS.n8536 9.3005
R7619 VSS.n8538 VSS.n8537 9.3005
R7620 VSS.n8539 VSS.n8538 9.3005
R7621 VSS.n8505 VSS.n8504 9.3005
R7622 VSS.n8505 VSS.n8255 9.3005
R7623 VSS.n8255 VSS.n8254 9.3005
R7624 VSS.n8485 VSS.n8484 9.3005
R7625 VSS.n8486 VSS.n8485 9.3005
R7626 VSS.n8545 VSS.n8544 9.3005
R7627 VSS.n8544 VSS.n8219 9.3005
R7628 VSS.n8219 VSS.n8218 9.3005
R7629 VSS.n8587 VSS.n8586 9.3005
R7630 VSS.n8586 VSS.n8585 9.3005
R7631 VSS.n8281 VSS.n8279 9.3005
R7632 VSS.n8629 VSS.n8628 9.3005
R7633 VSS.n8145 VSS.n8144 9.3005
R7634 VSS.n8679 VSS.n8170 9.3005
R7635 VSS.n8178 VSS.n8176 9.3005
R7636 VSS.n8644 VSS.n8643 9.3005
R7637 VSS.n8716 VSS.n8715 9.3005
R7638 VSS.n8716 VSS.n8150 9.3005
R7639 VSS.n8150 VSS.n8149 9.3005
R7640 VSS.n8698 VSS.n8158 9.3005
R7641 VSS.n8700 VSS.n8699 9.3005
R7642 VSS.n8692 VSS.n8691 9.3005
R7643 VSS.n8693 VSS.n8692 9.3005
R7644 VSS.n8694 VSS.n8693 9.3005
R7645 VSS.n8682 VSS.n8680 9.3005
R7646 VSS.n8660 VSS.n8171 9.3005
R7647 VSS.n8172 VSS.n8171 9.3005
R7648 VSS.n8674 VSS.n8172 9.3005
R7649 VSS.n8619 VSS.n8618 9.3005
R7650 VSS.n8619 VSS.n8193 9.3005
R7651 VSS.n8623 VSS.n8193 9.3005
R7652 VSS.n8630 VSS.n8190 9.3005
R7653 VSS.n8639 VSS.n8184 9.3005
R7654 VSS.n8184 VSS.n8174 9.3005
R7655 VSS.n8174 VSS.n8173 9.3005
R7656 VSS.n8642 VSS.n8183 9.3005
R7657 VSS.n8657 VSS.n8656 9.3005
R7658 VSS.n8725 VSS.n8724 9.3005
R7659 VSS.n8724 VSS.n8723 9.3005
R7660 VSS.n8572 VSS.n8210 9.3005
R7661 VSS.n8580 VSS.n8579 9.3005
R7662 VSS.n8579 VSS.n8578 9.3005
R7663 VSS.n8203 VSS.n8202 9.3005
R7664 VSS.n8571 VSS.n8202 9.3005
R7665 VSS.n8571 VSS.n8570 9.3005
R7666 VSS.n8609 VSS.n8201 9.3005
R7667 VSS.n8611 VSS.n8610 9.3005
R7668 VSS.n8343 VSS.n8339 9.3005
R7669 VSS.n8321 VSS.n8320 9.3005
R7670 VSS.n8301 VSS.n8300 9.3005
R7671 VSS.n8304 VSS.n8303 9.3005
R7672 VSS.n8431 VSS.n8430 9.3005
R7673 VSS.n8430 VSS.n8429 9.3005
R7674 VSS.n8429 VSS.n8428 9.3005
R7675 VSS.n8397 VSS.n8342 9.3005
R7676 VSS.n8397 VSS.n8396 9.3005
R7677 VSS.n8396 VSS.n8395 9.3005
R7678 VSS.n8386 VSS.n8348 9.3005
R7679 VSS.n8348 VSS.n8347 9.3005
R7680 VSS.n8454 VSS.n8453 9.3005
R7681 VSS.n8455 VSS.n8454 9.3005
R7682 VSS.n8456 VSS.n8455 9.3005
R7683 VSS.n8461 VSS.n8460 9.3005
R7684 VSS.n8460 VSS.n6481 9.3005
R7685 VSS.n8362 VSS.n8359 9.3005
R7686 VSS.n9084 VSS.n9083 9.3005
R7687 VSS.n9122 VSS.n9121 9.3005
R7688 VSS.n8813 VSS.n8812 9.3005
R7689 VSS.n9150 VSS.n9149 9.3005
R7690 VSS.n9129 VSS.n9128 9.3005
R7691 VSS.n9130 VSS.n9129 9.3005
R7692 VSS.n9131 VSS.n9130 9.3005
R7693 VSS.n9097 VSS.n9096 9.3005
R7694 VSS.n9097 VSS.n8847 9.3005
R7695 VSS.n8847 VSS.n8846 9.3005
R7696 VSS.n9077 VSS.n9076 9.3005
R7697 VSS.n9078 VSS.n9077 9.3005
R7698 VSS.n9137 VSS.n9136 9.3005
R7699 VSS.n9136 VSS.n8811 9.3005
R7700 VSS.n8811 VSS.n8810 9.3005
R7701 VSS.n9179 VSS.n9178 9.3005
R7702 VSS.n9178 VSS.n9177 9.3005
R7703 VSS.n8873 VSS.n8871 9.3005
R7704 VSS.n9221 VSS.n9220 9.3005
R7705 VSS.n8737 VSS.n8736 9.3005
R7706 VSS.n9271 VSS.n8762 9.3005
R7707 VSS.n8770 VSS.n8768 9.3005
R7708 VSS.n9236 VSS.n9235 9.3005
R7709 VSS.n9308 VSS.n9307 9.3005
R7710 VSS.n9308 VSS.n8742 9.3005
R7711 VSS.n8742 VSS.n8741 9.3005
R7712 VSS.n9290 VSS.n8750 9.3005
R7713 VSS.n9292 VSS.n9291 9.3005
R7714 VSS.n9284 VSS.n9283 9.3005
R7715 VSS.n9285 VSS.n9284 9.3005
R7716 VSS.n9286 VSS.n9285 9.3005
R7717 VSS.n9274 VSS.n9272 9.3005
R7718 VSS.n9252 VSS.n8763 9.3005
R7719 VSS.n8764 VSS.n8763 9.3005
R7720 VSS.n9266 VSS.n8764 9.3005
R7721 VSS.n9211 VSS.n9210 9.3005
R7722 VSS.n9211 VSS.n8785 9.3005
R7723 VSS.n9215 VSS.n8785 9.3005
R7724 VSS.n9222 VSS.n8782 9.3005
R7725 VSS.n9231 VSS.n8776 9.3005
R7726 VSS.n8776 VSS.n8766 9.3005
R7727 VSS.n8766 VSS.n8765 9.3005
R7728 VSS.n9234 VSS.n8775 9.3005
R7729 VSS.n9249 VSS.n9248 9.3005
R7730 VSS.n9317 VSS.n9316 9.3005
R7731 VSS.n9316 VSS.n9315 9.3005
R7732 VSS.n9164 VSS.n8802 9.3005
R7733 VSS.n9172 VSS.n9171 9.3005
R7734 VSS.n9171 VSS.n9170 9.3005
R7735 VSS.n8795 VSS.n8794 9.3005
R7736 VSS.n9163 VSS.n8794 9.3005
R7737 VSS.n9163 VSS.n9162 9.3005
R7738 VSS.n9201 VSS.n8793 9.3005
R7739 VSS.n9203 VSS.n9202 9.3005
R7740 VSS.n8935 VSS.n8931 9.3005
R7741 VSS.n8913 VSS.n8912 9.3005
R7742 VSS.n8893 VSS.n8892 9.3005
R7743 VSS.n8896 VSS.n8895 9.3005
R7744 VSS.n9023 VSS.n9022 9.3005
R7745 VSS.n9022 VSS.n9021 9.3005
R7746 VSS.n9021 VSS.n9020 9.3005
R7747 VSS.n8989 VSS.n8934 9.3005
R7748 VSS.n8989 VSS.n8988 9.3005
R7749 VSS.n8988 VSS.n8987 9.3005
R7750 VSS.n8978 VSS.n8940 9.3005
R7751 VSS.n8940 VSS.n8939 9.3005
R7752 VSS.n9046 VSS.n9045 9.3005
R7753 VSS.n9047 VSS.n9046 9.3005
R7754 VSS.n9048 VSS.n9047 9.3005
R7755 VSS.n9053 VSS.n9052 9.3005
R7756 VSS.n9052 VSS.n6482 9.3005
R7757 VSS.n8954 VSS.n8951 9.3005
R7758 VSS.n10268 VSS.n10267 9.3005
R7759 VSS.n10306 VSS.n10305 9.3005
R7760 VSS.n9997 VSS.n9996 9.3005
R7761 VSS.n10334 VSS.n10333 9.3005
R7762 VSS.n10313 VSS.n10312 9.3005
R7763 VSS.n10314 VSS.n10313 9.3005
R7764 VSS.n10315 VSS.n10314 9.3005
R7765 VSS.n10281 VSS.n10280 9.3005
R7766 VSS.n10281 VSS.n10031 9.3005
R7767 VSS.n10031 VSS.n10030 9.3005
R7768 VSS.n10261 VSS.n10260 9.3005
R7769 VSS.n10262 VSS.n10261 9.3005
R7770 VSS.n10321 VSS.n10320 9.3005
R7771 VSS.n10320 VSS.n9995 9.3005
R7772 VSS.n9995 VSS.n9994 9.3005
R7773 VSS.n10363 VSS.n10362 9.3005
R7774 VSS.n10362 VSS.n10361 9.3005
R7775 VSS.n10057 VSS.n10055 9.3005
R7776 VSS.n10405 VSS.n10404 9.3005
R7777 VSS.n9921 VSS.n9920 9.3005
R7778 VSS.n10455 VSS.n9946 9.3005
R7779 VSS.n9954 VSS.n9952 9.3005
R7780 VSS.n10420 VSS.n10419 9.3005
R7781 VSS.n10492 VSS.n10491 9.3005
R7782 VSS.n10492 VSS.n9926 9.3005
R7783 VSS.n9926 VSS.n9925 9.3005
R7784 VSS.n10474 VSS.n9934 9.3005
R7785 VSS.n10476 VSS.n10475 9.3005
R7786 VSS.n10468 VSS.n10467 9.3005
R7787 VSS.n10469 VSS.n10468 9.3005
R7788 VSS.n10470 VSS.n10469 9.3005
R7789 VSS.n10458 VSS.n10456 9.3005
R7790 VSS.n10436 VSS.n9947 9.3005
R7791 VSS.n9948 VSS.n9947 9.3005
R7792 VSS.n10450 VSS.n9948 9.3005
R7793 VSS.n10395 VSS.n10394 9.3005
R7794 VSS.n10395 VSS.n9969 9.3005
R7795 VSS.n10399 VSS.n9969 9.3005
R7796 VSS.n10406 VSS.n9966 9.3005
R7797 VSS.n10415 VSS.n9960 9.3005
R7798 VSS.n9960 VSS.n9950 9.3005
R7799 VSS.n9950 VSS.n9949 9.3005
R7800 VSS.n10418 VSS.n9959 9.3005
R7801 VSS.n10433 VSS.n10432 9.3005
R7802 VSS.n10501 VSS.n10500 9.3005
R7803 VSS.n10500 VSS.n10499 9.3005
R7804 VSS.n10348 VSS.n9986 9.3005
R7805 VSS.n10356 VSS.n10355 9.3005
R7806 VSS.n10355 VSS.n10354 9.3005
R7807 VSS.n9979 VSS.n9978 9.3005
R7808 VSS.n10347 VSS.n9978 9.3005
R7809 VSS.n10347 VSS.n10346 9.3005
R7810 VSS.n10385 VSS.n9977 9.3005
R7811 VSS.n10387 VSS.n10386 9.3005
R7812 VSS.n10119 VSS.n10115 9.3005
R7813 VSS.n10097 VSS.n10096 9.3005
R7814 VSS.n10077 VSS.n10076 9.3005
R7815 VSS.n10080 VSS.n10079 9.3005
R7816 VSS.n10207 VSS.n10206 9.3005
R7817 VSS.n10206 VSS.n10205 9.3005
R7818 VSS.n10205 VSS.n10204 9.3005
R7819 VSS.n10173 VSS.n10118 9.3005
R7820 VSS.n10173 VSS.n10172 9.3005
R7821 VSS.n10172 VSS.n10171 9.3005
R7822 VSS.n10162 VSS.n10124 9.3005
R7823 VSS.n10124 VSS.n10123 9.3005
R7824 VSS.n10230 VSS.n10229 9.3005
R7825 VSS.n10231 VSS.n10230 9.3005
R7826 VSS.n10232 VSS.n10231 9.3005
R7827 VSS.n10237 VSS.n10236 9.3005
R7828 VSS.n10236 VSS.n6484 9.3005
R7829 VSS.n10138 VSS.n10135 9.3005
R7830 VSS.n10860 VSS.n10859 9.3005
R7831 VSS.n10898 VSS.n10897 9.3005
R7832 VSS.n10589 VSS.n10588 9.3005
R7833 VSS.n10926 VSS.n10925 9.3005
R7834 VSS.n10905 VSS.n10904 9.3005
R7835 VSS.n10906 VSS.n10905 9.3005
R7836 VSS.n10907 VSS.n10906 9.3005
R7837 VSS.n10873 VSS.n10872 9.3005
R7838 VSS.n10873 VSS.n10623 9.3005
R7839 VSS.n10623 VSS.n10622 9.3005
R7840 VSS.n10853 VSS.n10852 9.3005
R7841 VSS.n10854 VSS.n10853 9.3005
R7842 VSS.n10913 VSS.n10912 9.3005
R7843 VSS.n10912 VSS.n10587 9.3005
R7844 VSS.n10587 VSS.n10586 9.3005
R7845 VSS.n10955 VSS.n10954 9.3005
R7846 VSS.n10954 VSS.n10953 9.3005
R7847 VSS.n10649 VSS.n10647 9.3005
R7848 VSS.n10997 VSS.n10996 9.3005
R7849 VSS.n10513 VSS.n10512 9.3005
R7850 VSS.n11047 VSS.n10538 9.3005
R7851 VSS.n10546 VSS.n10544 9.3005
R7852 VSS.n11012 VSS.n11011 9.3005
R7853 VSS.n11084 VSS.n11083 9.3005
R7854 VSS.n11084 VSS.n10518 9.3005
R7855 VSS.n10518 VSS.n10517 9.3005
R7856 VSS.n11066 VSS.n10526 9.3005
R7857 VSS.n11068 VSS.n11067 9.3005
R7858 VSS.n11060 VSS.n11059 9.3005
R7859 VSS.n11061 VSS.n11060 9.3005
R7860 VSS.n11062 VSS.n11061 9.3005
R7861 VSS.n11050 VSS.n11048 9.3005
R7862 VSS.n11028 VSS.n10539 9.3005
R7863 VSS.n10540 VSS.n10539 9.3005
R7864 VSS.n11042 VSS.n10540 9.3005
R7865 VSS.n10987 VSS.n10986 9.3005
R7866 VSS.n10987 VSS.n10561 9.3005
R7867 VSS.n10991 VSS.n10561 9.3005
R7868 VSS.n10998 VSS.n10558 9.3005
R7869 VSS.n11007 VSS.n10552 9.3005
R7870 VSS.n10552 VSS.n10542 9.3005
R7871 VSS.n10542 VSS.n10541 9.3005
R7872 VSS.n11010 VSS.n10551 9.3005
R7873 VSS.n11025 VSS.n11024 9.3005
R7874 VSS.n11093 VSS.n11092 9.3005
R7875 VSS.n11092 VSS.n11091 9.3005
R7876 VSS.n10940 VSS.n10578 9.3005
R7877 VSS.n10948 VSS.n10947 9.3005
R7878 VSS.n10947 VSS.n10946 9.3005
R7879 VSS.n10571 VSS.n10570 9.3005
R7880 VSS.n10939 VSS.n10570 9.3005
R7881 VSS.n10939 VSS.n10938 9.3005
R7882 VSS.n10977 VSS.n10569 9.3005
R7883 VSS.n10979 VSS.n10978 9.3005
R7884 VSS.n10711 VSS.n10707 9.3005
R7885 VSS.n10689 VSS.n10688 9.3005
R7886 VSS.n10669 VSS.n10668 9.3005
R7887 VSS.n10672 VSS.n10671 9.3005
R7888 VSS.n10799 VSS.n10798 9.3005
R7889 VSS.n10798 VSS.n10797 9.3005
R7890 VSS.n10797 VSS.n10796 9.3005
R7891 VSS.n10765 VSS.n10710 9.3005
R7892 VSS.n10765 VSS.n10764 9.3005
R7893 VSS.n10764 VSS.n10763 9.3005
R7894 VSS.n10754 VSS.n10716 9.3005
R7895 VSS.n10716 VSS.n10715 9.3005
R7896 VSS.n10822 VSS.n10821 9.3005
R7897 VSS.n10823 VSS.n10822 9.3005
R7898 VSS.n10824 VSS.n10823 9.3005
R7899 VSS.n10829 VSS.n10828 9.3005
R7900 VSS.n10828 VSS.n6485 9.3005
R7901 VSS.n10730 VSS.n10727 9.3005
R7902 VSS.n11452 VSS.n11451 9.3005
R7903 VSS.n11490 VSS.n11489 9.3005
R7904 VSS.n11181 VSS.n11180 9.3005
R7905 VSS.n11518 VSS.n11517 9.3005
R7906 VSS.n11497 VSS.n11496 9.3005
R7907 VSS.n11498 VSS.n11497 9.3005
R7908 VSS.n11499 VSS.n11498 9.3005
R7909 VSS.n11465 VSS.n11464 9.3005
R7910 VSS.n11465 VSS.n11215 9.3005
R7911 VSS.n11215 VSS.n11214 9.3005
R7912 VSS.n11445 VSS.n11444 9.3005
R7913 VSS.n11446 VSS.n11445 9.3005
R7914 VSS.n11505 VSS.n11504 9.3005
R7915 VSS.n11504 VSS.n11179 9.3005
R7916 VSS.n11179 VSS.n11178 9.3005
R7917 VSS.n11547 VSS.n11546 9.3005
R7918 VSS.n11546 VSS.n11545 9.3005
R7919 VSS.n11241 VSS.n11239 9.3005
R7920 VSS.n11589 VSS.n11588 9.3005
R7921 VSS.n11105 VSS.n11104 9.3005
R7922 VSS.n11639 VSS.n11130 9.3005
R7923 VSS.n11138 VSS.n11136 9.3005
R7924 VSS.n11604 VSS.n11603 9.3005
R7925 VSS.n11676 VSS.n11675 9.3005
R7926 VSS.n11676 VSS.n11110 9.3005
R7927 VSS.n11110 VSS.n11109 9.3005
R7928 VSS.n11658 VSS.n11118 9.3005
R7929 VSS.n11660 VSS.n11659 9.3005
R7930 VSS.n11652 VSS.n11651 9.3005
R7931 VSS.n11653 VSS.n11652 9.3005
R7932 VSS.n11654 VSS.n11653 9.3005
R7933 VSS.n11642 VSS.n11640 9.3005
R7934 VSS.n11620 VSS.n11131 9.3005
R7935 VSS.n11132 VSS.n11131 9.3005
R7936 VSS.n11634 VSS.n11132 9.3005
R7937 VSS.n11579 VSS.n11578 9.3005
R7938 VSS.n11579 VSS.n11153 9.3005
R7939 VSS.n11583 VSS.n11153 9.3005
R7940 VSS.n11590 VSS.n11150 9.3005
R7941 VSS.n11599 VSS.n11144 9.3005
R7942 VSS.n11144 VSS.n11134 9.3005
R7943 VSS.n11134 VSS.n11133 9.3005
R7944 VSS.n11602 VSS.n11143 9.3005
R7945 VSS.n11617 VSS.n11616 9.3005
R7946 VSS.n11685 VSS.n11684 9.3005
R7947 VSS.n11684 VSS.n11683 9.3005
R7948 VSS.n11532 VSS.n11170 9.3005
R7949 VSS.n11540 VSS.n11539 9.3005
R7950 VSS.n11539 VSS.n11538 9.3005
R7951 VSS.n11163 VSS.n11162 9.3005
R7952 VSS.n11531 VSS.n11162 9.3005
R7953 VSS.n11531 VSS.n11530 9.3005
R7954 VSS.n11569 VSS.n11161 9.3005
R7955 VSS.n11571 VSS.n11570 9.3005
R7956 VSS.n11303 VSS.n11299 9.3005
R7957 VSS.n11281 VSS.n11280 9.3005
R7958 VSS.n11261 VSS.n11260 9.3005
R7959 VSS.n11264 VSS.n11263 9.3005
R7960 VSS.n11391 VSS.n11390 9.3005
R7961 VSS.n11390 VSS.n11389 9.3005
R7962 VSS.n11389 VSS.n11388 9.3005
R7963 VSS.n11357 VSS.n11302 9.3005
R7964 VSS.n11357 VSS.n11356 9.3005
R7965 VSS.n11356 VSS.n11355 9.3005
R7966 VSS.n11346 VSS.n11308 9.3005
R7967 VSS.n11308 VSS.n11307 9.3005
R7968 VSS.n11414 VSS.n11413 9.3005
R7969 VSS.n11415 VSS.n11414 9.3005
R7970 VSS.n11416 VSS.n11415 9.3005
R7971 VSS.n11421 VSS.n11420 9.3005
R7972 VSS.n11420 VSS.n6486 9.3005
R7973 VSS.n11322 VSS.n11319 9.3005
R7974 VSS.n12044 VSS.n12043 9.3005
R7975 VSS.n12082 VSS.n12081 9.3005
R7976 VSS.n11773 VSS.n11772 9.3005
R7977 VSS.n12110 VSS.n12109 9.3005
R7978 VSS.n12089 VSS.n12088 9.3005
R7979 VSS.n12090 VSS.n12089 9.3005
R7980 VSS.n12091 VSS.n12090 9.3005
R7981 VSS.n12057 VSS.n12056 9.3005
R7982 VSS.n12057 VSS.n11807 9.3005
R7983 VSS.n11807 VSS.n11806 9.3005
R7984 VSS.n12037 VSS.n12036 9.3005
R7985 VSS.n12038 VSS.n12037 9.3005
R7986 VSS.n12097 VSS.n12096 9.3005
R7987 VSS.n12096 VSS.n11771 9.3005
R7988 VSS.n11771 VSS.n11770 9.3005
R7989 VSS.n12139 VSS.n12138 9.3005
R7990 VSS.n12138 VSS.n12137 9.3005
R7991 VSS.n11833 VSS.n11831 9.3005
R7992 VSS.n12181 VSS.n12180 9.3005
R7993 VSS.n11697 VSS.n11696 9.3005
R7994 VSS.n12231 VSS.n11722 9.3005
R7995 VSS.n11730 VSS.n11728 9.3005
R7996 VSS.n12196 VSS.n12195 9.3005
R7997 VSS.n12268 VSS.n12267 9.3005
R7998 VSS.n12268 VSS.n11702 9.3005
R7999 VSS.n11702 VSS.n11701 9.3005
R8000 VSS.n12250 VSS.n11710 9.3005
R8001 VSS.n12252 VSS.n12251 9.3005
R8002 VSS.n12244 VSS.n12243 9.3005
R8003 VSS.n12245 VSS.n12244 9.3005
R8004 VSS.n12246 VSS.n12245 9.3005
R8005 VSS.n12234 VSS.n12232 9.3005
R8006 VSS.n12212 VSS.n11723 9.3005
R8007 VSS.n11724 VSS.n11723 9.3005
R8008 VSS.n12226 VSS.n11724 9.3005
R8009 VSS.n12171 VSS.n12170 9.3005
R8010 VSS.n12171 VSS.n11745 9.3005
R8011 VSS.n12175 VSS.n11745 9.3005
R8012 VSS.n12182 VSS.n11742 9.3005
R8013 VSS.n12191 VSS.n11736 9.3005
R8014 VSS.n11736 VSS.n11726 9.3005
R8015 VSS.n11726 VSS.n11725 9.3005
R8016 VSS.n12194 VSS.n11735 9.3005
R8017 VSS.n12209 VSS.n12208 9.3005
R8018 VSS.n12277 VSS.n12276 9.3005
R8019 VSS.n12276 VSS.n12275 9.3005
R8020 VSS.n12124 VSS.n11762 9.3005
R8021 VSS.n12132 VSS.n12131 9.3005
R8022 VSS.n12131 VSS.n12130 9.3005
R8023 VSS.n11755 VSS.n11754 9.3005
R8024 VSS.n12123 VSS.n11754 9.3005
R8025 VSS.n12123 VSS.n12122 9.3005
R8026 VSS.n12161 VSS.n11753 9.3005
R8027 VSS.n12163 VSS.n12162 9.3005
R8028 VSS.n11895 VSS.n11891 9.3005
R8029 VSS.n11873 VSS.n11872 9.3005
R8030 VSS.n11853 VSS.n11852 9.3005
R8031 VSS.n11856 VSS.n11855 9.3005
R8032 VSS.n11983 VSS.n11982 9.3005
R8033 VSS.n11982 VSS.n11981 9.3005
R8034 VSS.n11981 VSS.n11980 9.3005
R8035 VSS.n11949 VSS.n11894 9.3005
R8036 VSS.n11949 VSS.n11948 9.3005
R8037 VSS.n11948 VSS.n11947 9.3005
R8038 VSS.n11938 VSS.n11900 9.3005
R8039 VSS.n11900 VSS.n11899 9.3005
R8040 VSS.n12006 VSS.n12005 9.3005
R8041 VSS.n12007 VSS.n12006 9.3005
R8042 VSS.n12008 VSS.n12007 9.3005
R8043 VSS.n12013 VSS.n12012 9.3005
R8044 VSS.n12012 VSS.n6487 9.3005
R8045 VSS.n11914 VSS.n11911 9.3005
R8046 VSS.n12636 VSS.n12635 9.3005
R8047 VSS.n12674 VSS.n12673 9.3005
R8048 VSS.n12365 VSS.n12364 9.3005
R8049 VSS.n12702 VSS.n12701 9.3005
R8050 VSS.n12681 VSS.n12680 9.3005
R8051 VSS.n12682 VSS.n12681 9.3005
R8052 VSS.n12683 VSS.n12682 9.3005
R8053 VSS.n12649 VSS.n12648 9.3005
R8054 VSS.n12649 VSS.n12399 9.3005
R8055 VSS.n12399 VSS.n12398 9.3005
R8056 VSS.n12629 VSS.n12628 9.3005
R8057 VSS.n12630 VSS.n12629 9.3005
R8058 VSS.n12689 VSS.n12688 9.3005
R8059 VSS.n12688 VSS.n12363 9.3005
R8060 VSS.n12363 VSS.n12362 9.3005
R8061 VSS.n12731 VSS.n12730 9.3005
R8062 VSS.n12730 VSS.n12729 9.3005
R8063 VSS.n12425 VSS.n12423 9.3005
R8064 VSS.n12773 VSS.n12772 9.3005
R8065 VSS.n12289 VSS.n12288 9.3005
R8066 VSS.n12823 VSS.n12314 9.3005
R8067 VSS.n12322 VSS.n12320 9.3005
R8068 VSS.n12788 VSS.n12787 9.3005
R8069 VSS.n12860 VSS.n12859 9.3005
R8070 VSS.n12860 VSS.n12294 9.3005
R8071 VSS.n12294 VSS.n12293 9.3005
R8072 VSS.n12842 VSS.n12302 9.3005
R8073 VSS.n12844 VSS.n12843 9.3005
R8074 VSS.n12836 VSS.n12835 9.3005
R8075 VSS.n12837 VSS.n12836 9.3005
R8076 VSS.n12838 VSS.n12837 9.3005
R8077 VSS.n12826 VSS.n12824 9.3005
R8078 VSS.n12804 VSS.n12315 9.3005
R8079 VSS.n12316 VSS.n12315 9.3005
R8080 VSS.n12818 VSS.n12316 9.3005
R8081 VSS.n12763 VSS.n12762 9.3005
R8082 VSS.n12763 VSS.n12337 9.3005
R8083 VSS.n12767 VSS.n12337 9.3005
R8084 VSS.n12774 VSS.n12334 9.3005
R8085 VSS.n12783 VSS.n12328 9.3005
R8086 VSS.n12328 VSS.n12318 9.3005
R8087 VSS.n12318 VSS.n12317 9.3005
R8088 VSS.n12786 VSS.n12327 9.3005
R8089 VSS.n12801 VSS.n12800 9.3005
R8090 VSS.n12869 VSS.n12868 9.3005
R8091 VSS.n12868 VSS.n12867 9.3005
R8092 VSS.n12716 VSS.n12354 9.3005
R8093 VSS.n12724 VSS.n12723 9.3005
R8094 VSS.n12723 VSS.n12722 9.3005
R8095 VSS.n12347 VSS.n12346 9.3005
R8096 VSS.n12715 VSS.n12346 9.3005
R8097 VSS.n12715 VSS.n12714 9.3005
R8098 VSS.n12753 VSS.n12345 9.3005
R8099 VSS.n12755 VSS.n12754 9.3005
R8100 VSS.n12487 VSS.n12483 9.3005
R8101 VSS.n12465 VSS.n12464 9.3005
R8102 VSS.n12445 VSS.n12444 9.3005
R8103 VSS.n12448 VSS.n12447 9.3005
R8104 VSS.n12575 VSS.n12574 9.3005
R8105 VSS.n12574 VSS.n12573 9.3005
R8106 VSS.n12573 VSS.n12572 9.3005
R8107 VSS.n12541 VSS.n12486 9.3005
R8108 VSS.n12541 VSS.n12540 9.3005
R8109 VSS.n12540 VSS.n12539 9.3005
R8110 VSS.n12530 VSS.n12492 9.3005
R8111 VSS.n12492 VSS.n12491 9.3005
R8112 VSS.n12598 VSS.n12597 9.3005
R8113 VSS.n12599 VSS.n12598 9.3005
R8114 VSS.n12600 VSS.n12599 9.3005
R8115 VSS.n12605 VSS.n12604 9.3005
R8116 VSS.n12604 VSS.n6488 9.3005
R8117 VSS.n12506 VSS.n12503 9.3005
R8118 VSS.n13228 VSS.n13227 9.3005
R8119 VSS.n13266 VSS.n13265 9.3005
R8120 VSS.n12957 VSS.n12956 9.3005
R8121 VSS.n13294 VSS.n13293 9.3005
R8122 VSS.n13273 VSS.n13272 9.3005
R8123 VSS.n13274 VSS.n13273 9.3005
R8124 VSS.n13275 VSS.n13274 9.3005
R8125 VSS.n13241 VSS.n13240 9.3005
R8126 VSS.n13241 VSS.n12991 9.3005
R8127 VSS.n12991 VSS.n12990 9.3005
R8128 VSS.n13221 VSS.n13220 9.3005
R8129 VSS.n13222 VSS.n13221 9.3005
R8130 VSS.n13281 VSS.n13280 9.3005
R8131 VSS.n13280 VSS.n12955 9.3005
R8132 VSS.n12955 VSS.n12954 9.3005
R8133 VSS.n13323 VSS.n13322 9.3005
R8134 VSS.n13322 VSS.n13321 9.3005
R8135 VSS.n13017 VSS.n13015 9.3005
R8136 VSS.n13365 VSS.n13364 9.3005
R8137 VSS.n12881 VSS.n12880 9.3005
R8138 VSS.n13415 VSS.n12906 9.3005
R8139 VSS.n12914 VSS.n12912 9.3005
R8140 VSS.n13380 VSS.n13379 9.3005
R8141 VSS.n13452 VSS.n13451 9.3005
R8142 VSS.n13452 VSS.n12886 9.3005
R8143 VSS.n12886 VSS.n12885 9.3005
R8144 VSS.n13434 VSS.n12894 9.3005
R8145 VSS.n13436 VSS.n13435 9.3005
R8146 VSS.n13428 VSS.n13427 9.3005
R8147 VSS.n13429 VSS.n13428 9.3005
R8148 VSS.n13430 VSS.n13429 9.3005
R8149 VSS.n13418 VSS.n13416 9.3005
R8150 VSS.n13396 VSS.n12907 9.3005
R8151 VSS.n12908 VSS.n12907 9.3005
R8152 VSS.n13410 VSS.n12908 9.3005
R8153 VSS.n13355 VSS.n13354 9.3005
R8154 VSS.n13355 VSS.n12929 9.3005
R8155 VSS.n13359 VSS.n12929 9.3005
R8156 VSS.n13366 VSS.n12926 9.3005
R8157 VSS.n13375 VSS.n12920 9.3005
R8158 VSS.n12920 VSS.n12910 9.3005
R8159 VSS.n12910 VSS.n12909 9.3005
R8160 VSS.n13378 VSS.n12919 9.3005
R8161 VSS.n13393 VSS.n13392 9.3005
R8162 VSS.n13461 VSS.n13460 9.3005
R8163 VSS.n13460 VSS.n13459 9.3005
R8164 VSS.n13308 VSS.n12946 9.3005
R8165 VSS.n13316 VSS.n13315 9.3005
R8166 VSS.n13315 VSS.n13314 9.3005
R8167 VSS.n12939 VSS.n12938 9.3005
R8168 VSS.n13307 VSS.n12938 9.3005
R8169 VSS.n13307 VSS.n13306 9.3005
R8170 VSS.n13345 VSS.n12937 9.3005
R8171 VSS.n13347 VSS.n13346 9.3005
R8172 VSS.n13079 VSS.n13075 9.3005
R8173 VSS.n13057 VSS.n13056 9.3005
R8174 VSS.n13037 VSS.n13036 9.3005
R8175 VSS.n13040 VSS.n13039 9.3005
R8176 VSS.n13167 VSS.n13166 9.3005
R8177 VSS.n13166 VSS.n13165 9.3005
R8178 VSS.n13165 VSS.n13164 9.3005
R8179 VSS.n13133 VSS.n13078 9.3005
R8180 VSS.n13133 VSS.n13132 9.3005
R8181 VSS.n13132 VSS.n13131 9.3005
R8182 VSS.n13122 VSS.n13084 9.3005
R8183 VSS.n13084 VSS.n13083 9.3005
R8184 VSS.n13190 VSS.n13189 9.3005
R8185 VSS.n13191 VSS.n13190 9.3005
R8186 VSS.n13192 VSS.n13191 9.3005
R8187 VSS.n13197 VSS.n13196 9.3005
R8188 VSS.n13196 VSS.n6489 9.3005
R8189 VSS.n13098 VSS.n13095 9.3005
R8190 VSS.n13820 VSS.n13819 9.3005
R8191 VSS.n13858 VSS.n13857 9.3005
R8192 VSS.n13549 VSS.n13548 9.3005
R8193 VSS.n13886 VSS.n13885 9.3005
R8194 VSS.n13865 VSS.n13864 9.3005
R8195 VSS.n13866 VSS.n13865 9.3005
R8196 VSS.n13867 VSS.n13866 9.3005
R8197 VSS.n13833 VSS.n13832 9.3005
R8198 VSS.n13833 VSS.n13583 9.3005
R8199 VSS.n13583 VSS.n13582 9.3005
R8200 VSS.n13813 VSS.n13812 9.3005
R8201 VSS.n13814 VSS.n13813 9.3005
R8202 VSS.n13873 VSS.n13872 9.3005
R8203 VSS.n13872 VSS.n13547 9.3005
R8204 VSS.n13547 VSS.n13546 9.3005
R8205 VSS.n13915 VSS.n13914 9.3005
R8206 VSS.n13914 VSS.n13913 9.3005
R8207 VSS.n13609 VSS.n13607 9.3005
R8208 VSS.n13957 VSS.n13956 9.3005
R8209 VSS.n13473 VSS.n13472 9.3005
R8210 VSS.n14007 VSS.n13498 9.3005
R8211 VSS.n13506 VSS.n13504 9.3005
R8212 VSS.n13972 VSS.n13971 9.3005
R8213 VSS.n14044 VSS.n14043 9.3005
R8214 VSS.n14044 VSS.n13478 9.3005
R8215 VSS.n13478 VSS.n13477 9.3005
R8216 VSS.n14026 VSS.n13486 9.3005
R8217 VSS.n14028 VSS.n14027 9.3005
R8218 VSS.n14020 VSS.n14019 9.3005
R8219 VSS.n14021 VSS.n14020 9.3005
R8220 VSS.n14022 VSS.n14021 9.3005
R8221 VSS.n14010 VSS.n14008 9.3005
R8222 VSS.n13988 VSS.n13499 9.3005
R8223 VSS.n13500 VSS.n13499 9.3005
R8224 VSS.n14002 VSS.n13500 9.3005
R8225 VSS.n13947 VSS.n13946 9.3005
R8226 VSS.n13947 VSS.n13521 9.3005
R8227 VSS.n13951 VSS.n13521 9.3005
R8228 VSS.n13958 VSS.n13518 9.3005
R8229 VSS.n13967 VSS.n13512 9.3005
R8230 VSS.n13512 VSS.n13502 9.3005
R8231 VSS.n13502 VSS.n13501 9.3005
R8232 VSS.n13970 VSS.n13511 9.3005
R8233 VSS.n13985 VSS.n13984 9.3005
R8234 VSS.n14053 VSS.n14052 9.3005
R8235 VSS.n14052 VSS.n14051 9.3005
R8236 VSS.n13900 VSS.n13538 9.3005
R8237 VSS.n13908 VSS.n13907 9.3005
R8238 VSS.n13907 VSS.n13906 9.3005
R8239 VSS.n13531 VSS.n13530 9.3005
R8240 VSS.n13899 VSS.n13530 9.3005
R8241 VSS.n13899 VSS.n13898 9.3005
R8242 VSS.n13937 VSS.n13529 9.3005
R8243 VSS.n13939 VSS.n13938 9.3005
R8244 VSS.n13671 VSS.n13667 9.3005
R8245 VSS.n13649 VSS.n13648 9.3005
R8246 VSS.n13629 VSS.n13628 9.3005
R8247 VSS.n13632 VSS.n13631 9.3005
R8248 VSS.n13759 VSS.n13758 9.3005
R8249 VSS.n13758 VSS.n13757 9.3005
R8250 VSS.n13757 VSS.n13756 9.3005
R8251 VSS.n13725 VSS.n13670 9.3005
R8252 VSS.n13725 VSS.n13724 9.3005
R8253 VSS.n13724 VSS.n13723 9.3005
R8254 VSS.n13714 VSS.n13676 9.3005
R8255 VSS.n13676 VSS.n13675 9.3005
R8256 VSS.n13782 VSS.n13781 9.3005
R8257 VSS.n13783 VSS.n13782 9.3005
R8258 VSS.n13784 VSS.n13783 9.3005
R8259 VSS.n13789 VSS.n13788 9.3005
R8260 VSS.n13788 VSS.n6490 9.3005
R8261 VSS.n13690 VSS.n13687 9.3005
R8262 VSS.n14412 VSS.n14411 9.3005
R8263 VSS.n14450 VSS.n14449 9.3005
R8264 VSS.n14141 VSS.n14140 9.3005
R8265 VSS.n14478 VSS.n14477 9.3005
R8266 VSS.n14457 VSS.n14456 9.3005
R8267 VSS.n14458 VSS.n14457 9.3005
R8268 VSS.n14459 VSS.n14458 9.3005
R8269 VSS.n14425 VSS.n14424 9.3005
R8270 VSS.n14425 VSS.n14175 9.3005
R8271 VSS.n14175 VSS.n14174 9.3005
R8272 VSS.n14405 VSS.n14404 9.3005
R8273 VSS.n14406 VSS.n14405 9.3005
R8274 VSS.n14465 VSS.n14464 9.3005
R8275 VSS.n14464 VSS.n14139 9.3005
R8276 VSS.n14139 VSS.n14138 9.3005
R8277 VSS.n14507 VSS.n14506 9.3005
R8278 VSS.n14506 VSS.n14505 9.3005
R8279 VSS.n14201 VSS.n14199 9.3005
R8280 VSS.n14549 VSS.n14548 9.3005
R8281 VSS.n14065 VSS.n14064 9.3005
R8282 VSS.n14599 VSS.n14090 9.3005
R8283 VSS.n14098 VSS.n14096 9.3005
R8284 VSS.n14564 VSS.n14563 9.3005
R8285 VSS.n14636 VSS.n14635 9.3005
R8286 VSS.n14636 VSS.n14070 9.3005
R8287 VSS.n14070 VSS.n14069 9.3005
R8288 VSS.n14618 VSS.n14078 9.3005
R8289 VSS.n14620 VSS.n14619 9.3005
R8290 VSS.n14612 VSS.n14611 9.3005
R8291 VSS.n14613 VSS.n14612 9.3005
R8292 VSS.n14614 VSS.n14613 9.3005
R8293 VSS.n14602 VSS.n14600 9.3005
R8294 VSS.n14580 VSS.n14091 9.3005
R8295 VSS.n14092 VSS.n14091 9.3005
R8296 VSS.n14594 VSS.n14092 9.3005
R8297 VSS.n14539 VSS.n14538 9.3005
R8298 VSS.n14539 VSS.n14113 9.3005
R8299 VSS.n14543 VSS.n14113 9.3005
R8300 VSS.n14550 VSS.n14110 9.3005
R8301 VSS.n14559 VSS.n14104 9.3005
R8302 VSS.n14104 VSS.n14094 9.3005
R8303 VSS.n14094 VSS.n14093 9.3005
R8304 VSS.n14562 VSS.n14103 9.3005
R8305 VSS.n14577 VSS.n14576 9.3005
R8306 VSS.n14645 VSS.n14644 9.3005
R8307 VSS.n14644 VSS.n14643 9.3005
R8308 VSS.n14492 VSS.n14130 9.3005
R8309 VSS.n14500 VSS.n14499 9.3005
R8310 VSS.n14499 VSS.n14498 9.3005
R8311 VSS.n14123 VSS.n14122 9.3005
R8312 VSS.n14491 VSS.n14122 9.3005
R8313 VSS.n14491 VSS.n14490 9.3005
R8314 VSS.n14529 VSS.n14121 9.3005
R8315 VSS.n14531 VSS.n14530 9.3005
R8316 VSS.n14263 VSS.n14259 9.3005
R8317 VSS.n14241 VSS.n14240 9.3005
R8318 VSS.n14221 VSS.n14220 9.3005
R8319 VSS.n14224 VSS.n14223 9.3005
R8320 VSS.n14351 VSS.n14350 9.3005
R8321 VSS.n14350 VSS.n14349 9.3005
R8322 VSS.n14349 VSS.n14348 9.3005
R8323 VSS.n14317 VSS.n14262 9.3005
R8324 VSS.n14317 VSS.n14316 9.3005
R8325 VSS.n14316 VSS.n14315 9.3005
R8326 VSS.n14306 VSS.n14268 9.3005
R8327 VSS.n14268 VSS.n14267 9.3005
R8328 VSS.n14374 VSS.n14373 9.3005
R8329 VSS.n14375 VSS.n14374 9.3005
R8330 VSS.n14376 VSS.n14375 9.3005
R8331 VSS.n14381 VSS.n14380 9.3005
R8332 VSS.n14380 VSS.n6491 9.3005
R8333 VSS.n14282 VSS.n14279 9.3005
R8334 VSS.n15004 VSS.n15003 9.3005
R8335 VSS.n15042 VSS.n15041 9.3005
R8336 VSS.n14733 VSS.n14732 9.3005
R8337 VSS.n15070 VSS.n15069 9.3005
R8338 VSS.n15049 VSS.n15048 9.3005
R8339 VSS.n15050 VSS.n15049 9.3005
R8340 VSS.n15051 VSS.n15050 9.3005
R8341 VSS.n15017 VSS.n15016 9.3005
R8342 VSS.n15017 VSS.n14767 9.3005
R8343 VSS.n14767 VSS.n14766 9.3005
R8344 VSS.n14997 VSS.n14996 9.3005
R8345 VSS.n14998 VSS.n14997 9.3005
R8346 VSS.n15057 VSS.n15056 9.3005
R8347 VSS.n15056 VSS.n14731 9.3005
R8348 VSS.n14731 VSS.n14730 9.3005
R8349 VSS.n15099 VSS.n15098 9.3005
R8350 VSS.n15098 VSS.n15097 9.3005
R8351 VSS.n14793 VSS.n14791 9.3005
R8352 VSS.n15141 VSS.n15140 9.3005
R8353 VSS.n14657 VSS.n14656 9.3005
R8354 VSS.n15191 VSS.n14682 9.3005
R8355 VSS.n14690 VSS.n14688 9.3005
R8356 VSS.n15156 VSS.n15155 9.3005
R8357 VSS.n15228 VSS.n15227 9.3005
R8358 VSS.n15228 VSS.n14662 9.3005
R8359 VSS.n14662 VSS.n14661 9.3005
R8360 VSS.n15210 VSS.n14670 9.3005
R8361 VSS.n15212 VSS.n15211 9.3005
R8362 VSS.n15204 VSS.n15203 9.3005
R8363 VSS.n15205 VSS.n15204 9.3005
R8364 VSS.n15206 VSS.n15205 9.3005
R8365 VSS.n15194 VSS.n15192 9.3005
R8366 VSS.n15172 VSS.n14683 9.3005
R8367 VSS.n14684 VSS.n14683 9.3005
R8368 VSS.n15186 VSS.n14684 9.3005
R8369 VSS.n15131 VSS.n15130 9.3005
R8370 VSS.n15131 VSS.n14705 9.3005
R8371 VSS.n15135 VSS.n14705 9.3005
R8372 VSS.n15142 VSS.n14702 9.3005
R8373 VSS.n15151 VSS.n14696 9.3005
R8374 VSS.n14696 VSS.n14686 9.3005
R8375 VSS.n14686 VSS.n14685 9.3005
R8376 VSS.n15154 VSS.n14695 9.3005
R8377 VSS.n15169 VSS.n15168 9.3005
R8378 VSS.n15237 VSS.n15236 9.3005
R8379 VSS.n15236 VSS.n15235 9.3005
R8380 VSS.n15084 VSS.n14722 9.3005
R8381 VSS.n15092 VSS.n15091 9.3005
R8382 VSS.n15091 VSS.n15090 9.3005
R8383 VSS.n14715 VSS.n14714 9.3005
R8384 VSS.n15083 VSS.n14714 9.3005
R8385 VSS.n15083 VSS.n15082 9.3005
R8386 VSS.n15121 VSS.n14713 9.3005
R8387 VSS.n15123 VSS.n15122 9.3005
R8388 VSS.n14855 VSS.n14851 9.3005
R8389 VSS.n14833 VSS.n14832 9.3005
R8390 VSS.n14813 VSS.n14812 9.3005
R8391 VSS.n14816 VSS.n14815 9.3005
R8392 VSS.n14943 VSS.n14942 9.3005
R8393 VSS.n14942 VSS.n14941 9.3005
R8394 VSS.n14941 VSS.n14940 9.3005
R8395 VSS.n14909 VSS.n14854 9.3005
R8396 VSS.n14909 VSS.n14908 9.3005
R8397 VSS.n14908 VSS.n14907 9.3005
R8398 VSS.n14898 VSS.n14860 9.3005
R8399 VSS.n14860 VSS.n14859 9.3005
R8400 VSS.n14966 VSS.n14965 9.3005
R8401 VSS.n14967 VSS.n14966 9.3005
R8402 VSS.n14968 VSS.n14967 9.3005
R8403 VSS.n14973 VSS.n14972 9.3005
R8404 VSS.n14972 VSS.n6492 9.3005
R8405 VSS.n14874 VSS.n14871 9.3005
R8406 VSS.n15596 VSS.n15595 9.3005
R8407 VSS.n15634 VSS.n15633 9.3005
R8408 VSS.n15325 VSS.n15324 9.3005
R8409 VSS.n15662 VSS.n15661 9.3005
R8410 VSS.n15641 VSS.n15640 9.3005
R8411 VSS.n15642 VSS.n15641 9.3005
R8412 VSS.n15643 VSS.n15642 9.3005
R8413 VSS.n15609 VSS.n15608 9.3005
R8414 VSS.n15609 VSS.n15359 9.3005
R8415 VSS.n15359 VSS.n15358 9.3005
R8416 VSS.n15589 VSS.n15588 9.3005
R8417 VSS.n15590 VSS.n15589 9.3005
R8418 VSS.n15649 VSS.n15648 9.3005
R8419 VSS.n15648 VSS.n15323 9.3005
R8420 VSS.n15323 VSS.n15322 9.3005
R8421 VSS.n15691 VSS.n15690 9.3005
R8422 VSS.n15690 VSS.n15689 9.3005
R8423 VSS.n15385 VSS.n15383 9.3005
R8424 VSS.n15733 VSS.n15732 9.3005
R8425 VSS.n15249 VSS.n15248 9.3005
R8426 VSS.n15783 VSS.n15274 9.3005
R8427 VSS.n15282 VSS.n15280 9.3005
R8428 VSS.n15748 VSS.n15747 9.3005
R8429 VSS.n15820 VSS.n15819 9.3005
R8430 VSS.n15820 VSS.n15254 9.3005
R8431 VSS.n15254 VSS.n15253 9.3005
R8432 VSS.n15802 VSS.n15262 9.3005
R8433 VSS.n15804 VSS.n15803 9.3005
R8434 VSS.n15796 VSS.n15795 9.3005
R8435 VSS.n15797 VSS.n15796 9.3005
R8436 VSS.n15798 VSS.n15797 9.3005
R8437 VSS.n15786 VSS.n15784 9.3005
R8438 VSS.n15764 VSS.n15275 9.3005
R8439 VSS.n15276 VSS.n15275 9.3005
R8440 VSS.n15778 VSS.n15276 9.3005
R8441 VSS.n15723 VSS.n15722 9.3005
R8442 VSS.n15723 VSS.n15297 9.3005
R8443 VSS.n15727 VSS.n15297 9.3005
R8444 VSS.n15734 VSS.n15294 9.3005
R8445 VSS.n15743 VSS.n15288 9.3005
R8446 VSS.n15288 VSS.n15278 9.3005
R8447 VSS.n15278 VSS.n15277 9.3005
R8448 VSS.n15746 VSS.n15287 9.3005
R8449 VSS.n15761 VSS.n15760 9.3005
R8450 VSS.n15829 VSS.n15828 9.3005
R8451 VSS.n15828 VSS.n15827 9.3005
R8452 VSS.n15676 VSS.n15314 9.3005
R8453 VSS.n15684 VSS.n15683 9.3005
R8454 VSS.n15683 VSS.n15682 9.3005
R8455 VSS.n15307 VSS.n15306 9.3005
R8456 VSS.n15675 VSS.n15306 9.3005
R8457 VSS.n15675 VSS.n15674 9.3005
R8458 VSS.n15713 VSS.n15305 9.3005
R8459 VSS.n15715 VSS.n15714 9.3005
R8460 VSS.n15447 VSS.n15443 9.3005
R8461 VSS.n15425 VSS.n15424 9.3005
R8462 VSS.n15405 VSS.n15404 9.3005
R8463 VSS.n15408 VSS.n15407 9.3005
R8464 VSS.n15535 VSS.n15534 9.3005
R8465 VSS.n15534 VSS.n15533 9.3005
R8466 VSS.n15533 VSS.n15532 9.3005
R8467 VSS.n15501 VSS.n15446 9.3005
R8468 VSS.n15501 VSS.n15500 9.3005
R8469 VSS.n15500 VSS.n15499 9.3005
R8470 VSS.n15490 VSS.n15452 9.3005
R8471 VSS.n15452 VSS.n15451 9.3005
R8472 VSS.n15558 VSS.n15557 9.3005
R8473 VSS.n15559 VSS.n15558 9.3005
R8474 VSS.n15560 VSS.n15559 9.3005
R8475 VSS.n15565 VSS.n15564 9.3005
R8476 VSS.n15564 VSS.n6493 9.3005
R8477 VSS.n15466 VSS.n15463 9.3005
R8478 VSS.n6759 VSS.n6758 9.3005
R8479 VSS.n6780 VSS.n6779 9.3005
R8480 VSS.n6720 VSS.n6719 9.3005
R8481 VSS.n6801 VSS.n6800 9.3005
R8482 VSS.n6786 VSS.n6785 9.3005
R8483 VSS.n6787 VSS.n6786 9.3005
R8484 VSS.n6788 VSS.n6787 9.3005
R8485 VSS.n6767 VSS.n6733 9.3005
R8486 VSS.n6767 VSS.n6766 9.3005
R8487 VSS.n6766 VSS.n6765 9.3005
R8488 VSS.n6752 VSS.n6736 9.3005
R8489 VSS.n6736 VSS.n6735 9.3005
R8490 VSS.n6792 VSS.n6723 9.3005
R8491 VSS.n6792 VSS.n6718 9.3005
R8492 VSS.n6718 VSS.n6717 9.3005
R8493 VSS.n15924 VSS.n15923 9.3005
R8494 VSS.n15923 VSS.n15922 9.3005
R8495 VSS.n15967 VSS.n15966 9.3005
R8496 VSS.n15888 VSS.n15887 9.3005
R8497 VSS.n15843 VSS.n15842 9.3005
R8498 VSS.n15869 VSS.n15868 9.3005
R8499 VSS.n6864 VSS.n6862 9.3005
R8500 VSS.n6882 VSS.n6881 9.3005
R8501 VSS.n15850 VSS.n6908 9.3005
R8502 VSS.n15850 VSS.n15849 9.3005
R8503 VSS.n15849 VSS.n15848 9.3005
R8504 VSS.n6928 VSS.n6899 9.3005
R8505 VSS.n6909 VSS.n6907 9.3005
R8506 VSS.n6898 VSS.n6894 9.3005
R8507 VSS.n6927 VSS.n6894 9.3005
R8508 VSS.n6927 VSS.n6913 9.3005
R8509 VSS.n15867 VSS.n6892 9.3005
R8510 VSS.n6921 VSS.n6920 9.3005
R8511 VSS.n6921 VSS.n6860 9.3005
R8512 VSS.n6860 VSS.n6859 9.3005
R8513 VSS.n15895 VSS.n15894 9.3005
R8514 VSS.n15896 VSS.n15895 9.3005
R8515 VSS.n15897 VSS.n15896 9.3005
R8516 VSS.n15889 VSS.n6855 9.3005
R8517 VSS.n6877 VSS.n6857 9.3005
R8518 VSS.n6858 VSS.n6857 9.3005
R8519 VSS.n15882 VSS.n6858 9.3005
R8520 VSS.n6880 VSS.n6869 9.3005
R8521 VSS.n6916 VSS.n6915 9.3005
R8522 VSS.n6942 VSS.n6934 9.3005
R8523 VSS.n6934 VSS.n6933 9.3005
R8524 VSS.n6823 VSS.n6822 9.3005
R8525 VSS.n15917 VSS.n15916 9.3005
R8526 VSS.n15916 VSS.n15915 9.3005
R8527 VSS.n15910 VSS.n15909 9.3005
R8528 VSS.n15910 VSS.n6812 9.3005
R8529 VSS.n6812 VSS.n6811 9.3005
R8530 VSS.n15904 VSS.n15903 9.3005
R8531 VSS.n15902 VSS.n6838 9.3005
R8532 VSS.n6555 VSS.n6551 9.3005
R8533 VSS.n6533 VSS.n6532 9.3005
R8534 VSS.n6513 VSS.n6512 9.3005
R8535 VSS.n6516 VSS.n6515 9.3005
R8536 VSS.n6643 VSS.n6642 9.3005
R8537 VSS.n6642 VSS.n6641 9.3005
R8538 VSS.n6641 VSS.n6640 9.3005
R8539 VSS.n6609 VSS.n6554 9.3005
R8540 VSS.n6609 VSS.n6608 9.3005
R8541 VSS.n6608 VSS.n6607 9.3005
R8542 VSS.n6598 VSS.n6560 9.3005
R8543 VSS.n6560 VSS.n6559 9.3005
R8544 VSS.n6666 VSS.n6665 9.3005
R8545 VSS.n6667 VSS.n6666 9.3005
R8546 VSS.n6668 VSS.n6667 9.3005
R8547 VSS.n6673 VSS.n6672 9.3005
R8548 VSS.n6672 VSS.n6494 9.3005
R8549 VSS.n6574 VSS.n6571 9.3005
R8550 VSS.n7308 VSS.n7307 9.3005
R8551 VSS.n7346 VSS.n7345 9.3005
R8552 VSS.n7036 VSS.n7035 9.3005
R8553 VSS.n7374 VSS.n7373 9.3005
R8554 VSS.n7353 VSS.n7352 9.3005
R8555 VSS.n7354 VSS.n7353 9.3005
R8556 VSS.n7355 VSS.n7354 9.3005
R8557 VSS.n7321 VSS.n7320 9.3005
R8558 VSS.n7321 VSS.n7070 9.3005
R8559 VSS.n7070 VSS.n7069 9.3005
R8560 VSS.n7301 VSS.n7300 9.3005
R8561 VSS.n7302 VSS.n7301 9.3005
R8562 VSS.n7361 VSS.n7360 9.3005
R8563 VSS.n7360 VSS.n7034 9.3005
R8564 VSS.n7034 VSS.n7033 9.3005
R8565 VSS.n7403 VSS.n7402 9.3005
R8566 VSS.n7402 VSS.n7401 9.3005
R8567 VSS.n7096 VSS.n7094 9.3005
R8568 VSS.n7445 VSS.n7444 9.3005
R8569 VSS.n6960 VSS.n6959 9.3005
R8570 VSS.n7495 VSS.n6985 9.3005
R8571 VSS.n6993 VSS.n6991 9.3005
R8572 VSS.n7460 VSS.n7459 9.3005
R8573 VSS.n7532 VSS.n7531 9.3005
R8574 VSS.n7532 VSS.n6965 9.3005
R8575 VSS.n6965 VSS.n6964 9.3005
R8576 VSS.n7514 VSS.n6973 9.3005
R8577 VSS.n7516 VSS.n7515 9.3005
R8578 VSS.n7508 VSS.n7507 9.3005
R8579 VSS.n7509 VSS.n7508 9.3005
R8580 VSS.n7510 VSS.n7509 9.3005
R8581 VSS.n7498 VSS.n7496 9.3005
R8582 VSS.n7476 VSS.n6986 9.3005
R8583 VSS.n6987 VSS.n6986 9.3005
R8584 VSS.n7490 VSS.n6987 9.3005
R8585 VSS.n7435 VSS.n7434 9.3005
R8586 VSS.n7435 VSS.n7008 9.3005
R8587 VSS.n7439 VSS.n7008 9.3005
R8588 VSS.n7446 VSS.n7005 9.3005
R8589 VSS.n7455 VSS.n6999 9.3005
R8590 VSS.n6999 VSS.n6989 9.3005
R8591 VSS.n6989 VSS.n6988 9.3005
R8592 VSS.n7458 VSS.n6998 9.3005
R8593 VSS.n7473 VSS.n7472 9.3005
R8594 VSS.n7541 VSS.n7540 9.3005
R8595 VSS.n7540 VSS.n7539 9.3005
R8596 VSS.n7388 VSS.n7025 9.3005
R8597 VSS.n7396 VSS.n7395 9.3005
R8598 VSS.n7395 VSS.n7394 9.3005
R8599 VSS.n7018 VSS.n7017 9.3005
R8600 VSS.n7387 VSS.n7017 9.3005
R8601 VSS.n7387 VSS.n7386 9.3005
R8602 VSS.n7425 VSS.n7016 9.3005
R8603 VSS.n7427 VSS.n7426 9.3005
R8604 VSS.n7203 VSS.n7202 9.3005
R8605 VSS.n7241 VSS.n7240 9.3005
R8606 VSS.n7111 VSS.n7110 9.3005
R8607 VSS.n7270 VSS.n7269 9.3005
R8608 VSS.n7248 VSS.n7247 9.3005
R8609 VSS.n7249 VSS.n7248 9.3005
R8610 VSS.n7250 VSS.n7249 9.3005
R8611 VSS.n7216 VSS.n7215 9.3005
R8612 VSS.n7216 VSS.n7147 9.3005
R8613 VSS.n7147 VSS.n7146 9.3005
R8614 VSS.n7196 VSS.n7195 9.3005
R8615 VSS.n7197 VSS.n7196 9.3005
R8616 VSS.n7257 VSS.n7256 9.3005
R8617 VSS.n7256 VSS.n7109 9.3005
R8618 VSS.n7109 VSS.n7108 9.3005
R8619 VSS.n7277 VSS.n7276 9.3005
R8620 VSS.n7276 VSS.n7275 9.3005
R8621 VSS.n7171 VSS.n7169 9.3005
R8622 VSS.n18620 VSS.n18619 9.3005
R8623 VSS.n18658 VSS.n18657 9.3005
R8624 VSS.n134 VSS.n133 9.3005
R8625 VSS.n18686 VSS.n18685 9.3005
R8626 VSS.n18665 VSS.n18664 9.3005
R8627 VSS.n18666 VSS.n18665 9.3005
R8628 VSS.n18667 VSS.n18666 9.3005
R8629 VSS.n18633 VSS.n18632 9.3005
R8630 VSS.n18633 VSS.n168 9.3005
R8631 VSS.n168 VSS.n167 9.3005
R8632 VSS.n18613 VSS.n18612 9.3005
R8633 VSS.n18614 VSS.n18613 9.3005
R8634 VSS.n18673 VSS.n18672 9.3005
R8635 VSS.n18672 VSS.n132 9.3005
R8636 VSS.n132 VSS.n131 9.3005
R8637 VSS.n18715 VSS.n18714 9.3005
R8638 VSS.n18714 VSS.n18713 9.3005
R8639 VSS.n206 VSS.n205 9.3005
R8640 VSS.n18757 VSS.n18756 9.3005
R8641 VSS.n58 VSS.n57 9.3005
R8642 VSS.n18807 VSS.n83 9.3005
R8643 VSS.n91 VSS.n89 9.3005
R8644 VSS.n18772 VSS.n18771 9.3005
R8645 VSS.n18844 VSS.n18843 9.3005
R8646 VSS.n18844 VSS.n63 9.3005
R8647 VSS.n63 VSS.n62 9.3005
R8648 VSS.n18826 VSS.n71 9.3005
R8649 VSS.n18828 VSS.n18827 9.3005
R8650 VSS.n18820 VSS.n18819 9.3005
R8651 VSS.n18821 VSS.n18820 9.3005
R8652 VSS.n18822 VSS.n18821 9.3005
R8653 VSS.n18810 VSS.n18808 9.3005
R8654 VSS.n18788 VSS.n84 9.3005
R8655 VSS.n85 VSS.n84 9.3005
R8656 VSS.n18802 VSS.n85 9.3005
R8657 VSS.n18747 VSS.n18746 9.3005
R8658 VSS.n18747 VSS.n106 9.3005
R8659 VSS.n18751 VSS.n106 9.3005
R8660 VSS.n18758 VSS.n103 9.3005
R8661 VSS.n18767 VSS.n97 9.3005
R8662 VSS.n97 VSS.n87 9.3005
R8663 VSS.n87 VSS.n86 9.3005
R8664 VSS.n18770 VSS.n96 9.3005
R8665 VSS.n18785 VSS.n18784 9.3005
R8666 VSS.n18853 VSS.n18852 9.3005
R8667 VSS.n18852 VSS.n18851 9.3005
R8668 VSS.n18700 VSS.n123 9.3005
R8669 VSS.n18708 VSS.n18707 9.3005
R8670 VSS.n18707 VSS.n18706 9.3005
R8671 VSS.n116 VSS.n115 9.3005
R8672 VSS.n18699 VSS.n115 9.3005
R8673 VSS.n18699 VSS.n18698 9.3005
R8674 VSS.n18737 VSS.n114 9.3005
R8675 VSS.n18739 VSS.n18738 9.3005
R8676 VSS.n366 VSS.n365 9.3005
R8677 VSS.n393 VSS.n392 9.3005
R8678 VSS.n406 VSS.n405 9.3005
R8679 VSS.n404 VSS.n325 9.3005
R8680 VSS.n387 VSS.n386 9.3005
R8681 VSS.n386 VSS.n385 9.3005
R8682 VSS.n385 VSS.n384 9.3005
R8683 VSS.n371 VSS.n370 9.3005
R8684 VSS.n372 VSS.n371 9.3005
R8685 VSS.n373 VSS.n372 9.3005
R8686 VSS.n344 VSS.n343 9.3005
R8687 VSS.n360 VSS.n344 9.3005
R8688 VSS.n396 VSS.n395 9.3005
R8689 VSS.n396 VSS.n329 9.3005
R8690 VSS.n400 VSS.n329 9.3005
R8691 VSS.n18589 VSS.n18588 9.3005
R8692 VSS.n18588 VSS.n18587 9.3005
R8693 VSS.n453 VSS.n452 9.3005
R8694 VSS.n18285 VSS.n18284 9.3005
R8695 VSS.n18286 VSS.n18285 9.3005
R8696 VSS.n18287 VSS.n18286 9.3005
R8697 VSS.n18266 VSS.n18232 9.3005
R8698 VSS.n18266 VSS.n18265 9.3005
R8699 VSS.n18265 VSS.n18264 9.3005
R8700 VSS.n18251 VSS.n18235 9.3005
R8701 VSS.n18235 VSS.n18234 9.3005
R8702 VSS.n18291 VSS.n18222 9.3005
R8703 VSS.n18291 VSS.n18217 9.3005
R8704 VSS.n18217 VSS.n18216 9.3005
R8705 VSS.n18541 VSS.n18540 9.3005
R8706 VSS.n18540 VSS.n18539 9.3005
R8707 VSS.n18584 VSS.n18583 9.3005
R8708 VSS.n18423 VSS.n18421 9.3005
R8709 VSS.n18453 VSS.n18421 9.3005
R8710 VSS.n18453 VSS.n18439 9.3005
R8711 VSS.n18448 VSS.n18447 9.3005
R8712 VSS.n18449 VSS.n18448 9.3005
R8713 VSS.n18450 VSS.n18449 9.3005
R8714 VSS.n18407 VSS.n18386 9.3005
R8715 VSS.n18386 VSS.n18360 9.3005
R8716 VSS.n18495 VSS.n18360 9.3005
R8717 VSS.n18343 VSS.n18340 9.3005
R8718 VSS.n18372 VSS.n18343 9.3005
R8719 VSS.n18372 VSS.n18371 9.3005
R8720 VSS.n18379 VSS.n18378 9.3005
R8721 VSS.n18379 VSS.n18359 9.3005
R8722 VSS.n18383 VSS.n18359 9.3005
R8723 VSS.n18462 VSS.n18461 9.3005
R8724 VSS.n18461 VSS.n18460 9.3005
R8725 VSS.n18534 VSS.n18533 9.3005
R8726 VSS.n18533 VSS.n18532 9.3005
R8727 VSS.n18527 VSS.n18526 9.3005
R8728 VSS.n18527 VSS.n18311 9.3005
R8729 VSS.n18311 VSS.n18310 9.3005
R8730 VSS.n582 VSS.n581 9.3005
R8731 VSS.n603 VSS.n602 9.3005
R8732 VSS.n540 VSS.n539 9.3005
R8733 VSS.n624 VSS.n623 9.3005
R8734 VSS.n609 VSS.n608 9.3005
R8735 VSS.n610 VSS.n609 9.3005
R8736 VSS.n611 VSS.n610 9.3005
R8737 VSS.n590 VSS.n553 9.3005
R8738 VSS.n590 VSS.n589 9.3005
R8739 VSS.n589 VSS.n588 9.3005
R8740 VSS.n575 VSS.n556 9.3005
R8741 VSS.n556 VSS.n555 9.3005
R8742 VSS.n615 VSS.n543 9.3005
R8743 VSS.n615 VSS.n538 9.3005
R8744 VSS.n538 VSS.n537 9.3005
R8745 VSS.n838 VSS.n837 9.3005
R8746 VSS.n837 VSS.n836 9.3005
R8747 VSS.n560 VSS.n559 9.3005
R8748 VSS.n18866 VSS.n18865 9.3005
R8749 VSS.n764 VSS.n730 9.3005
R8750 VSS.n783 VSS.n782 9.3005
R8751 VSS.n781 VSS.n715 9.3005
R8752 VSS.n748 VSS.n747 9.3005
R8753 VSS.n705 VSS.n704 9.3005
R8754 VSS.n818 VSS.n817 9.3005
R8755 VSS.n831 VSS.n830 9.3005
R8756 VSS.n830 VSS.n829 9.3005
R8757 VSS.n646 VSS.n645 9.3005
R8758 VSS.n816 VSS.n661 9.3005
R8759 VSS.n824 VSS.n823 9.3005
R8760 VSS.n824 VSS.n635 9.3005
R8761 VSS.n635 VSS.n634 9.3005
R8762 VSS.n809 VSS.n808 9.3005
R8763 VSS.n810 VSS.n809 9.3005
R8764 VSS.n811 VSS.n810 9.3005
R8765 VSS.n803 VSS.n678 9.3005
R8766 VSS.n802 VSS.n801 9.3005
R8767 VSS.n700 VSS.n680 9.3005
R8768 VSS.n681 VSS.n680 9.3005
R8769 VSS.n796 VSS.n681 9.3005
R8770 VSS.n703 VSS.n692 9.3005
R8771 VSS.n687 VSS.n685 9.3005
R8772 VSS.n753 VSS.n752 9.3005
R8773 VSS.n753 VSS.n683 9.3005
R8774 VSS.n683 VSS.n682 9.3005
R8775 VSS.n721 VSS.n717 9.3005
R8776 VSS.n758 VSS.n717 9.3005
R8777 VSS.n759 VSS.n758 9.3005
R8778 VSS.n763 VSS.n722 9.3005
R8779 VSS.n742 VSS.n48 9.3005
R8780 VSS.n48 VSS.n47 9.3005
R8781 VSS.n47 VSS.n46 9.3005
R8782 VSS.n18874 VSS.n18873 9.3005
R8783 VSS.n18873 VSS.n18872 9.3005
R8784 VSS.n925 VSS.n924 9.3005
R8785 VSS.n946 VSS.n945 9.3005
R8786 VSS.n887 VSS.n886 9.3005
R8787 VSS.n968 VSS.n967 9.3005
R8788 VSS.n952 VSS.n951 9.3005
R8789 VSS.n953 VSS.n952 9.3005
R8790 VSS.n954 VSS.n953 9.3005
R8791 VSS.n933 VSS.n901 9.3005
R8792 VSS.n933 VSS.n932 9.3005
R8793 VSS.n932 VSS.n931 9.3005
R8794 VSS.n920 VSS.n904 9.3005
R8795 VSS.n904 VSS.n903 9.3005
R8796 VSS.n959 VSS.n890 9.3005
R8797 VSS.n959 VSS.n885 9.3005
R8798 VSS.n885 VSS.n884 9.3005
R8799 VSS.n975 VSS.n974 9.3005
R8800 VSS.n974 VSS.n973 9.3005
R8801 VSS.n1018 VSS.n1017 9.3005
R8802 VSS.n1133 VSS.n1132 9.3005
R8803 VSS.n1134 VSS.n1133 9.3005
R8804 VSS.n1135 VSS.n1134 9.3005
R8805 VSS.n1114 VSS.n1082 9.3005
R8806 VSS.n1114 VSS.n1113 9.3005
R8807 VSS.n1113 VSS.n1112 9.3005
R8808 VSS.n1101 VSS.n1085 9.3005
R8809 VSS.n1085 VSS.n1084 9.3005
R8810 VSS.n1140 VSS.n1071 9.3005
R8811 VSS.n1140 VSS.n1066 9.3005
R8812 VSS.n1066 VSS.n1065 9.3005
R8813 VSS.n18001 VSS.n18000 9.3005
R8814 VSS.n18000 VSS.n17999 9.3005
R8815 VSS.n18044 VSS.n18043 9.3005
R8816 VSS.n17565 VSS.n17564 9.3005
R8817 VSS.n17564 VSS.n17563 9.3005
R8818 VSS.n17563 VSS.n17562 9.3005
R8819 VSS.n17531 VSS.n17476 9.3005
R8820 VSS.n17531 VSS.n17530 9.3005
R8821 VSS.n17530 VSS.n17529 9.3005
R8822 VSS.n17520 VSS.n17482 9.3005
R8823 VSS.n17482 VSS.n17481 9.3005
R8824 VSS.n17588 VSS.n17587 9.3005
R8825 VSS.n17589 VSS.n17588 9.3005
R8826 VSS.n17590 VSS.n17589 9.3005
R8827 VSS.n17595 VSS.n17594 9.3005
R8828 VSS.n17594 VSS.n1155 9.3005
R8829 VSS.n17496 VSS.n17493 9.3005
R8830 VSS.n1268 VSS.n1267 9.3005
R8831 VSS.n1269 VSS.n1268 9.3005
R8832 VSS.n1270 VSS.n1269 9.3005
R8833 VSS.n1249 VSS.n1215 9.3005
R8834 VSS.n1249 VSS.n1248 9.3005
R8835 VSS.n1248 VSS.n1247 9.3005
R8836 VSS.n1234 VSS.n1218 9.3005
R8837 VSS.n1218 VSS.n1217 9.3005
R8838 VSS.n1274 VSS.n1205 9.3005
R8839 VSS.n1274 VSS.n1200 9.3005
R8840 VSS.n1200 VSS.n1199 9.3005
R8841 VSS.n17952 VSS.n17951 9.3005
R8842 VSS.n17951 VSS.n17950 9.3005
R8843 VSS.n17995 VSS.n17994 9.3005
R8844 VSS.n17916 VSS.n17915 9.3005
R8845 VSS.n17871 VSS.n17870 9.3005
R8846 VSS.n17897 VSS.n17896 9.3005
R8847 VSS.n1346 VSS.n1344 9.3005
R8848 VSS.n1364 VSS.n1363 9.3005
R8849 VSS.n17878 VSS.n1390 9.3005
R8850 VSS.n17878 VSS.n17877 9.3005
R8851 VSS.n17877 VSS.n17876 9.3005
R8852 VSS.n1410 VSS.n1381 9.3005
R8853 VSS.n1391 VSS.n1389 9.3005
R8854 VSS.n1380 VSS.n1376 9.3005
R8855 VSS.n1409 VSS.n1376 9.3005
R8856 VSS.n1409 VSS.n1395 9.3005
R8857 VSS.n17895 VSS.n1374 9.3005
R8858 VSS.n1403 VSS.n1402 9.3005
R8859 VSS.n1403 VSS.n1342 9.3005
R8860 VSS.n1342 VSS.n1341 9.3005
R8861 VSS.n17923 VSS.n17922 9.3005
R8862 VSS.n17924 VSS.n17923 9.3005
R8863 VSS.n17925 VSS.n17924 9.3005
R8864 VSS.n17917 VSS.n1337 9.3005
R8865 VSS.n1359 VSS.n1339 9.3005
R8866 VSS.n1340 VSS.n1339 9.3005
R8867 VSS.n17910 VSS.n1340 9.3005
R8868 VSS.n1362 VSS.n1351 9.3005
R8869 VSS.n1398 VSS.n1397 9.3005
R8870 VSS.n1424 VSS.n1416 9.3005
R8871 VSS.n1416 VSS.n1415 9.3005
R8872 VSS.n1305 VSS.n1304 9.3005
R8873 VSS.n17945 VSS.n17944 9.3005
R8874 VSS.n17944 VSS.n17943 9.3005
R8875 VSS.n17938 VSS.n17937 9.3005
R8876 VSS.n17938 VSS.n1294 9.3005
R8877 VSS.n1294 VSS.n1293 9.3005
R8878 VSS.n17932 VSS.n17931 9.3005
R8879 VSS.n17930 VSS.n1320 9.3005
R8880 VSS.n17055 VSS.n17054 9.15497
R8881 VSS.n17054 VSS.n17053 9.15497
R8882 VSS.n17647 VSS.n17646 9.15497
R8883 VSS.n17646 VSS.n17645 9.15497
R8884 VSS.n18132 VSS.n251 9.15497
R8885 VSS.n251 VSS.n250 9.15497
R8886 VSS.n9697 VSS.n9696 9.15497
R8887 VSS.n9696 VSS.n9695 9.15497
R8888 VSS.n9605 VSS.n9509 9.15497
R8889 VSS.n9509 VSS.n9508 9.15497
R8890 VSS.n16640 VSS.n16639 9.15497
R8891 VSS.n16639 VSS.n16638 9.15497
R8892 VSS.n16535 VSS.n16534 9.15497
R8893 VSS.n16534 VSS.n16533 9.15497
R8894 VSS.n16047 VSS.n16046 9.15497
R8895 VSS.n16046 VSS.n16045 9.15497
R8896 VSS.n1700 VSS.n1699 9.15497
R8897 VSS.n1699 VSS.n1698 9.15497
R8898 VSS.n1993 VSS.n1992 9.15497
R8899 VSS.n2036 VSS.n1993 9.15497
R8900 VSS.n1897 VSS.n1801 9.15497
R8901 VSS.n1801 VSS.n1800 9.15497
R8902 VSS.n3188 VSS.n3187 9.15497
R8903 VSS.n3187 VSS.n3186 9.15497
R8904 VSS.n3096 VSS.n3000 9.15497
R8905 VSS.n3000 VSS.n2999 9.15497
R8906 VSS.n3780 VSS.n3779 9.15497
R8907 VSS.n3779 VSS.n3778 9.15497
R8908 VSS.n3688 VSS.n3592 9.15497
R8909 VSS.n3592 VSS.n3591 9.15497
R8910 VSS.n4372 VSS.n4371 9.15497
R8911 VSS.n4371 VSS.n4370 9.15497
R8912 VSS.n4280 VSS.n4184 9.15497
R8913 VSS.n4184 VSS.n4183 9.15497
R8914 VSS.n4964 VSS.n4963 9.15497
R8915 VSS.n4963 VSS.n4962 9.15497
R8916 VSS.n4872 VSS.n4776 9.15497
R8917 VSS.n4776 VSS.n4775 9.15497
R8918 VSS.n2589 VSS.n2588 9.15497
R8919 VSS.n2632 VSS.n2589 9.15497
R8920 VSS.n2493 VSS.n2397 9.15497
R8921 VSS.n2397 VSS.n2396 9.15497
R8922 VSS.n5550 VSS.n5549 9.15497
R8923 VSS.n5593 VSS.n5550 9.15497
R8924 VSS.n5454 VSS.n5358 9.15497
R8925 VSS.n5358 VSS.n5357 9.15497
R8926 VSS.n6123 VSS.n6122 9.15497
R8927 VSS.n6166 VSS.n6123 9.15497
R8928 VSS.n6027 VSS.n5931 9.15497
R8929 VSS.n5931 VSS.n5930 9.15497
R8930 VSS.n7921 VSS.n7920 9.15497
R8931 VSS.n7920 VSS.n7919 9.15497
R8932 VSS.n7829 VSS.n7733 9.15497
R8933 VSS.n7733 VSS.n7732 9.15497
R8934 VSS.n8513 VSS.n8512 9.15497
R8935 VSS.n8512 VSS.n8511 9.15497
R8936 VSS.n8421 VSS.n8325 9.15497
R8937 VSS.n8325 VSS.n8324 9.15497
R8938 VSS.n9105 VSS.n9104 9.15497
R8939 VSS.n9104 VSS.n9103 9.15497
R8940 VSS.n9013 VSS.n8917 9.15497
R8941 VSS.n8917 VSS.n8916 9.15497
R8942 VSS.n10289 VSS.n10288 9.15497
R8943 VSS.n10288 VSS.n10287 9.15497
R8944 VSS.n10197 VSS.n10101 9.15497
R8945 VSS.n10101 VSS.n10100 9.15497
R8946 VSS.n10881 VSS.n10880 9.15497
R8947 VSS.n10880 VSS.n10879 9.15497
R8948 VSS.n10789 VSS.n10693 9.15497
R8949 VSS.n10693 VSS.n10692 9.15497
R8950 VSS.n11473 VSS.n11472 9.15497
R8951 VSS.n11472 VSS.n11471 9.15497
R8952 VSS.n11381 VSS.n11285 9.15497
R8953 VSS.n11285 VSS.n11284 9.15497
R8954 VSS.n12065 VSS.n12064 9.15497
R8955 VSS.n12064 VSS.n12063 9.15497
R8956 VSS.n11973 VSS.n11877 9.15497
R8957 VSS.n11877 VSS.n11876 9.15497
R8958 VSS.n12657 VSS.n12656 9.15497
R8959 VSS.n12656 VSS.n12655 9.15497
R8960 VSS.n12565 VSS.n12469 9.15497
R8961 VSS.n12469 VSS.n12468 9.15497
R8962 VSS.n13249 VSS.n13248 9.15497
R8963 VSS.n13248 VSS.n13247 9.15497
R8964 VSS.n13157 VSS.n13061 9.15497
R8965 VSS.n13061 VSS.n13060 9.15497
R8966 VSS.n13841 VSS.n13840 9.15497
R8967 VSS.n13840 VSS.n13839 9.15497
R8968 VSS.n13749 VSS.n13653 9.15497
R8969 VSS.n13653 VSS.n13652 9.15497
R8970 VSS.n14433 VSS.n14432 9.15497
R8971 VSS.n14432 VSS.n14431 9.15497
R8972 VSS.n14341 VSS.n14245 9.15497
R8973 VSS.n14245 VSS.n14244 9.15497
R8974 VSS.n15025 VSS.n15024 9.15497
R8975 VSS.n15024 VSS.n15023 9.15497
R8976 VSS.n14933 VSS.n14837 9.15497
R8977 VSS.n14837 VSS.n14836 9.15497
R8978 VSS.n15617 VSS.n15616 9.15497
R8979 VSS.n15616 VSS.n15615 9.15497
R8980 VSS.n15525 VSS.n15429 9.15497
R8981 VSS.n15429 VSS.n15428 9.15497
R8982 VSS.n6729 VSS.n6728 9.15497
R8983 VSS.n6772 VSS.n6729 9.15497
R8984 VSS.n6633 VSS.n6537 9.15497
R8985 VSS.n6537 VSS.n6536 9.15497
R8986 VSS.n7329 VSS.n7328 9.15497
R8987 VSS.n7328 VSS.n7327 9.15497
R8988 VSS.n7224 VSS.n7223 9.15497
R8989 VSS.n7223 VSS.n7222 9.15497
R8990 VSS.n18641 VSS.n18640 9.15497
R8991 VSS.n18640 VSS.n18639 9.15497
R8992 VSS.n379 VSS.n337 9.15497
R8993 VSS.n337 VSS.n336 9.15497
R8994 VSS.n18228 VSS.n18227 9.15497
R8995 VSS.n18271 VSS.n18228 9.15497
R8996 VSS.n549 VSS.n548 9.15497
R8997 VSS.n595 VSS.n549 9.15497
R8998 VSS.n897 VSS.n896 9.15497
R8999 VSS.n938 VSS.n897 9.15497
R9000 VSS.n1078 VSS.n1077 9.15497
R9001 VSS.n1119 VSS.n1078 9.15497
R9002 VSS.n17555 VSS.n17459 9.15497
R9003 VSS.n17459 VSS.n17458 9.15497
R9004 VSS.n1211 VSS.n1210 9.15497
R9005 VSS.n1254 VSS.n1211 9.15497
R9006 VSS.n17994 VSS.n1157 8.44336
R9007 VSS.n17951 VSS.n1198 8.44336
R9008 VSS.n17499 VSS.n17493 8.44336
R9009 VSS.n17594 VSS.n17593 8.44336
R9010 VSS.n18043 VSS.n1022 8.44336
R9011 VSS.n18000 VSS.n1064 8.44336
R9012 VSS.n1017 VSS.n455 8.44336
R9013 VSS.n974 VSS.n883 8.44336
R9014 VSS.n17004 VSS.n16999 8.44336
R9015 VSS.n17128 VSS.n16937 8.44336
R9016 VSS.n17418 VSS.n17413 8.44336
R9017 VSS.n17720 VSS.n17351 8.44336
R9018 VSS.n18583 VSS.n210 8.44336
R9019 VSS.n18540 VSS.n18215 8.44336
R9020 VSS.n18076 VSS.n285 8.44336
R9021 VSS.n18171 VSS.n18170 8.44336
R9022 VSS.n9549 VSS.n9543 8.44336
R9023 VSS.n9644 VSS.n9643 8.44336
R9024 VSS.n9468 VSS.n9463 8.44336
R9025 VSS.n9770 VSS.n9401 8.44336
R9026 VSS.n16485 VSS.n16480 8.44336
R9027 VSS.n16587 VSS.n16418 8.44336
R9028 VSS.n16410 VSS.n16405 8.44336
R9029 VSS.n16713 VSS.n16343 8.44336
R9030 VSS.n1650 VSS.n1645 8.44336
R9031 VSS.n15994 VSS.n1583 8.44336
R9032 VSS.n1756 VSS.n1755 8.44336
R9033 VSS.n16120 VSS.n1515 8.44336
R9034 VSS.n1841 VSS.n1835 8.44336
R9035 VSS.n1936 VSS.n1935 8.44336
R9036 VSS.n2348 VSS.n1760 8.44336
R9037 VSS.n2305 VSS.n1980 8.44336
R9038 VSS.n3040 VSS.n3034 8.44336
R9039 VSS.n3135 VSS.n3134 8.44336
R9040 VSS.n2959 VSS.n2954 8.44336
R9041 VSS.n3261 VSS.n2892 8.44336
R9042 VSS.n3632 VSS.n3626 8.44336
R9043 VSS.n3727 VSS.n3726 8.44336
R9044 VSS.n3551 VSS.n3546 8.44336
R9045 VSS.n3853 VSS.n3484 8.44336
R9046 VSS.n4224 VSS.n4218 8.44336
R9047 VSS.n4319 VSS.n4318 8.44336
R9048 VSS.n4143 VSS.n4138 8.44336
R9049 VSS.n4445 VSS.n4076 8.44336
R9050 VSS.n4816 VSS.n4810 8.44336
R9051 VSS.n4911 VSS.n4910 8.44336
R9052 VSS.n4735 VSS.n4730 8.44336
R9053 VSS.n5037 VSS.n4668 8.44336
R9054 VSS.n2437 VSS.n2431 8.44336
R9055 VSS.n2532 VSS.n2531 8.44336
R9056 VSS.n5313 VSS.n2356 8.44336
R9057 VSS.n5270 VSS.n2576 8.44336
R9058 VSS.n5398 VSS.n5392 8.44336
R9059 VSS.n5493 VSS.n5492 8.44336
R9060 VSS.n5886 VSS.n5317 8.44336
R9061 VSS.n5843 VSS.n5537 8.44336
R9062 VSS.n5971 VSS.n5965 8.44336
R9063 VSS.n6066 VSS.n6065 8.44336
R9064 VSS.n6478 VSS.n5890 8.44336
R9065 VSS.n6435 VSS.n6110 8.44336
R9066 VSS.n7773 VSS.n7767 8.44336
R9067 VSS.n7868 VSS.n7867 8.44336
R9068 VSS.n7692 VSS.n7687 8.44336
R9069 VSS.n7994 VSS.n7625 8.44336
R9070 VSS.n8365 VSS.n8359 8.44336
R9071 VSS.n8460 VSS.n8459 8.44336
R9072 VSS.n8284 VSS.n8279 8.44336
R9073 VSS.n8586 VSS.n8217 8.44336
R9074 VSS.n8957 VSS.n8951 8.44336
R9075 VSS.n9052 VSS.n9051 8.44336
R9076 VSS.n8876 VSS.n8871 8.44336
R9077 VSS.n9178 VSS.n8809 8.44336
R9078 VSS.n10141 VSS.n10135 8.44336
R9079 VSS.n10236 VSS.n10235 8.44336
R9080 VSS.n10060 VSS.n10055 8.44336
R9081 VSS.n10362 VSS.n9993 8.44336
R9082 VSS.n10733 VSS.n10727 8.44336
R9083 VSS.n10828 VSS.n10827 8.44336
R9084 VSS.n10652 VSS.n10647 8.44336
R9085 VSS.n10954 VSS.n10585 8.44336
R9086 VSS.n11325 VSS.n11319 8.44336
R9087 VSS.n11420 VSS.n11419 8.44336
R9088 VSS.n11244 VSS.n11239 8.44336
R9089 VSS.n11546 VSS.n11177 8.44336
R9090 VSS.n11917 VSS.n11911 8.44336
R9091 VSS.n12012 VSS.n12011 8.44336
R9092 VSS.n11836 VSS.n11831 8.44336
R9093 VSS.n12138 VSS.n11769 8.44336
R9094 VSS.n12509 VSS.n12503 8.44336
R9095 VSS.n12604 VSS.n12603 8.44336
R9096 VSS.n12428 VSS.n12423 8.44336
R9097 VSS.n12730 VSS.n12361 8.44336
R9098 VSS.n13101 VSS.n13095 8.44336
R9099 VSS.n13196 VSS.n13195 8.44336
R9100 VSS.n13020 VSS.n13015 8.44336
R9101 VSS.n13322 VSS.n12953 8.44336
R9102 VSS.n13693 VSS.n13687 8.44336
R9103 VSS.n13788 VSS.n13787 8.44336
R9104 VSS.n13612 VSS.n13607 8.44336
R9105 VSS.n13914 VSS.n13545 8.44336
R9106 VSS.n14285 VSS.n14279 8.44336
R9107 VSS.n14380 VSS.n14379 8.44336
R9108 VSS.n14204 VSS.n14199 8.44336
R9109 VSS.n14506 VSS.n14137 8.44336
R9110 VSS.n14877 VSS.n14871 8.44336
R9111 VSS.n14972 VSS.n14971 8.44336
R9112 VSS.n14796 VSS.n14791 8.44336
R9113 VSS.n15098 VSS.n14729 8.44336
R9114 VSS.n15469 VSS.n15463 8.44336
R9115 VSS.n15564 VSS.n15563 8.44336
R9116 VSS.n15388 VSS.n15383 8.44336
R9117 VSS.n15690 VSS.n15321 8.44336
R9118 VSS.n6577 VSS.n6571 8.44336
R9119 VSS.n6672 VSS.n6671 8.44336
R9120 VSS.n15966 VSS.n6496 8.44336
R9121 VSS.n15923 VSS.n6716 8.44336
R9122 VSS.n7174 VSS.n7169 8.44336
R9123 VSS.n7276 VSS.n7107 8.44336
R9124 VSS.n7099 VSS.n7094 8.44336
R9125 VSS.n7402 VSS.n7032 8.44336
R9126 VSS.n452 VSS.n289 8.44336
R9127 VSS.n18588 VSS.n198 8.44336
R9128 VSS.n205 VSS.n204 8.44336
R9129 VSS.n18714 VSS.n130 8.44336
R9130 VSS.n559 VSS.n558 8.44336
R9131 VSS.n837 VSS.n536 8.44336
R9132 VSS.n17117 VSS.n17111 7.69581
R9133 VSS.n17260 VSS.n16866 7.69581
R9134 VSS.n17709 VSS.n17703 7.69581
R9135 VSS.n17852 VSS.n17280 7.69581
R9136 VSS.n18529 VSS.n18309 7.69581
R9137 VSS.n18456 VSS.n18437 7.69581
R9138 VSS.n9759 VSS.n9753 7.69581
R9139 VSS.n9903 VSS.n9331 7.69581
R9140 VSS.n16702 VSS.n16696 7.69581
R9141 VSS.n16846 VSS.n16273 7.69581
R9142 VSS.n16109 VSS.n16103 7.69581
R9143 VSS.n16253 VSS.n1445 7.69581
R9144 VSS.n2294 VSS.n2074 7.69581
R9145 VSS.n2227 VSS.n2176 7.69581
R9146 VSS.n3250 VSS.n3244 7.69581
R9147 VSS.n3394 VSS.n2822 7.69581
R9148 VSS.n3842 VSS.n3836 7.69581
R9149 VSS.n3986 VSS.n3414 7.69581
R9150 VSS.n4434 VSS.n4428 7.69581
R9151 VSS.n4578 VSS.n4006 7.69581
R9152 VSS.n5026 VSS.n5020 7.69581
R9153 VSS.n5170 VSS.n4598 7.69581
R9154 VSS.n5259 VSS.n2670 7.69581
R9155 VSS.n5192 VSS.n2772 7.69581
R9156 VSS.n5832 VSS.n5631 7.69581
R9157 VSS.n5746 VSS.n7 7.69581
R9158 VSS.n6424 VSS.n6204 7.69581
R9159 VSS.n6357 VSS.n6306 7.69581
R9160 VSS.n7983 VSS.n7977 7.69581
R9161 VSS.n8127 VSS.n7555 7.69581
R9162 VSS.n8575 VSS.n8569 7.69581
R9163 VSS.n8719 VSS.n8147 7.69581
R9164 VSS.n9167 VSS.n9161 7.69581
R9165 VSS.n9311 VSS.n8739 7.69581
R9166 VSS.n10351 VSS.n10345 7.69581
R9167 VSS.n10495 VSS.n9923 7.69581
R9168 VSS.n10943 VSS.n10937 7.69581
R9169 VSS.n11087 VSS.n10515 7.69581
R9170 VSS.n11535 VSS.n11529 7.69581
R9171 VSS.n11679 VSS.n11107 7.69581
R9172 VSS.n12127 VSS.n12121 7.69581
R9173 VSS.n12271 VSS.n11699 7.69581
R9174 VSS.n12719 VSS.n12713 7.69581
R9175 VSS.n12863 VSS.n12291 7.69581
R9176 VSS.n13311 VSS.n13305 7.69581
R9177 VSS.n13455 VSS.n12883 7.69581
R9178 VSS.n13903 VSS.n13897 7.69581
R9179 VSS.n14047 VSS.n13475 7.69581
R9180 VSS.n14495 VSS.n14489 7.69581
R9181 VSS.n14639 VSS.n14067 7.69581
R9182 VSS.n15087 VSS.n15081 7.69581
R9183 VSS.n15231 VSS.n14659 7.69581
R9184 VSS.n15679 VSS.n15673 7.69581
R9185 VSS.n15823 VSS.n15251 7.69581
R9186 VSS.n15912 VSS.n6810 7.69581
R9187 VSS.n15845 VSS.n6912 7.69581
R9188 VSS.n7391 VSS.n7385 7.69581
R9189 VSS.n7535 VSS.n6962 7.69581
R9190 VSS.n18703 VSS.n18697 7.69581
R9191 VSS.n18847 VSS.n60 7.69581
R9192 VSS.n826 VSS.n633 7.69581
R9193 VSS.n18869 VSS.n45 7.69581
R9194 VSS.n17940 VSS.n1292 7.69581
R9195 VSS.n17873 VSS.n1394 7.69581
R9196 VSS.n17911 VSS.n1323 7.61296
R9197 VSS.n1407 VSS.n1406 7.61296
R9198 VSS.n17590 VSS.t409 7.26922
R9199 VSS.n17167 VSS.n17166 6.39585
R9200 VSS.n17217 VSS.n16881 6.39585
R9201 VSS.n17759 VSS.n17758 6.39585
R9202 VSS.n17809 VSS.n17295 6.39585
R9203 VSS.n9809 VSS.n9808 6.39585
R9204 VSS.n9859 VSS.n9345 6.39585
R9205 VSS.n16752 VSS.n16751 6.39585
R9206 VSS.n16802 VSS.n16287 6.39585
R9207 VSS.n16159 VSS.n16158 6.39585
R9208 VSS.n16209 VSS.n1459 6.39585
R9209 VSS.n2265 VSS.n2105 6.39585
R9210 VSS.n2189 VSS.n2188 6.39585
R9211 VSS.n3300 VSS.n3299 6.39585
R9212 VSS.n3350 VSS.n2836 6.39585
R9213 VSS.n3892 VSS.n3891 6.39585
R9214 VSS.n3942 VSS.n3428 6.39585
R9215 VSS.n4484 VSS.n4483 6.39585
R9216 VSS.n4534 VSS.n4020 6.39585
R9217 VSS.n5076 VSS.n5075 6.39585
R9218 VSS.n5126 VSS.n4612 6.39585
R9219 VSS.n5230 VSS.n2701 6.39585
R9220 VSS.n2785 VSS.n2784 6.39585
R9221 VSS.n5803 VSS.n5662 6.39585
R9222 VSS.n5759 VSS.n5758 6.39585
R9223 VSS.n6395 VSS.n6235 6.39585
R9224 VSS.n6319 VSS.n6318 6.39585
R9225 VSS.n8033 VSS.n8032 6.39585
R9226 VSS.n8083 VSS.n7569 6.39585
R9227 VSS.n8625 VSS.n8624 6.39585
R9228 VSS.n8675 VSS.n8161 6.39585
R9229 VSS.n9217 VSS.n9216 6.39585
R9230 VSS.n9267 VSS.n8753 6.39585
R9231 VSS.n10401 VSS.n10400 6.39585
R9232 VSS.n10451 VSS.n9937 6.39585
R9233 VSS.n10993 VSS.n10992 6.39585
R9234 VSS.n11043 VSS.n10529 6.39585
R9235 VSS.n11585 VSS.n11584 6.39585
R9236 VSS.n11635 VSS.n11121 6.39585
R9237 VSS.n12177 VSS.n12176 6.39585
R9238 VSS.n12227 VSS.n11713 6.39585
R9239 VSS.n12769 VSS.n12768 6.39585
R9240 VSS.n12819 VSS.n12305 6.39585
R9241 VSS.n13361 VSS.n13360 6.39585
R9242 VSS.n13411 VSS.n12897 6.39585
R9243 VSS.n13953 VSS.n13952 6.39585
R9244 VSS.n14003 VSS.n13489 6.39585
R9245 VSS.n14545 VSS.n14544 6.39585
R9246 VSS.n14595 VSS.n14081 6.39585
R9247 VSS.n15137 VSS.n15136 6.39585
R9248 VSS.n15187 VSS.n14673 6.39585
R9249 VSS.n15729 VSS.n15728 6.39585
R9250 VSS.n15779 VSS.n15265 6.39585
R9251 VSS.n15883 VSS.n6841 6.39585
R9252 VSS.n6925 VSS.n6924 6.39585
R9253 VSS.n7441 VSS.n7440 6.39585
R9254 VSS.n7491 VSS.n6976 6.39585
R9255 VSS.n18753 VSS.n18752 6.39585
R9256 VSS.n18803 VSS.n74 6.39585
R9257 VSS.n18382 VSS.n18361 6.39585
R9258 VSS.n18494 VSS.n18384 6.39585
R9259 VSS.n797 VSS.n664 6.39585
R9260 VSS.n755 VSS.n745 6.39585
R9261 VSS.n10202 VSS.t635 6.22398
R9262 VSS.n18137 VSS.t466 6.21519
R9263 VSS.n16563 VSS.t528 6.21519
R9264 VSS.n1728 VSS.t323 6.21519
R9265 VSS.n1902 VSS.t206 6.21519
R9266 VSS.n3101 VSS.t281 6.21519
R9267 VSS.n3693 VSS.t264 6.21519
R9268 VSS.n4285 VSS.t320 6.21519
R9269 VSS.n4877 VSS.t191 6.21519
R9270 VSS.n2498 VSS.t148 6.21519
R9271 VSS.n5459 VSS.t383 6.21519
R9272 VSS.n6032 VSS.t55 6.21519
R9273 VSS.n7834 VSS.t427 6.21519
R9274 VSS.n8426 VSS.t200 6.21519
R9275 VSS.n9018 VSS.t108 6.21519
R9276 VSS.n10794 VSS.t303 6.21519
R9277 VSS.n11386 VSS.t534 6.21519
R9278 VSS.n11978 VSS.t602 6.21519
R9279 VSS.n12570 VSS.t623 6.21519
R9280 VSS.n13162 VSS.t193 6.21519
R9281 VSS.n13754 VSS.t367 6.21519
R9282 VSS.n14346 VSS.t300 6.21519
R9283 VSS.n14938 VSS.t403 6.21519
R9284 VSS.n15530 VSS.t470 6.21519
R9285 VSS.n6638 VSS.t435 6.21519
R9286 VSS.n7252 VSS.t502 6.21519
R9287 VSS.t13 VSS.n399 6.21519
R9288 VSS.n956 VSS.t234 6.21519
R9289 VSS.n1137 VSS.t255 6.21519
R9290 VSS.n9610 VSS.t249 6.20642
R9291 VSS.n1244 VSS.n1218 5.62907
R9292 VSS.n1272 VSS.n1200 5.62907
R9293 VSS.n17523 VSS.n17482 5.62907
R9294 VSS.n17589 VSS.n17427 5.62907
R9295 VSS.n1109 VSS.n1085 5.62907
R9296 VSS.n1138 VSS.n1066 5.62907
R9297 VSS.n928 VSS.n904 5.62907
R9298 VSS.n957 VSS.n885 5.62907
R9299 VSS.n17027 VSS.n16988 5.62907
R9300 VSS.n17083 VSS.n16939 5.62907
R9301 VSS.n17619 VSS.n17402 5.62907
R9302 VSS.n17675 VSS.n17353 5.62907
R9303 VSS.n18261 VSS.n18235 5.62907
R9304 VSS.n18289 VSS.n18217 5.62907
R9305 VSS.n18100 VSS.n274 5.62907
R9306 VSS.n18166 VSS.n219 5.62907
R9307 VSS.n9573 VSS.n9532 5.62907
R9308 VSS.n9639 VSS.n9477 5.62907
R9309 VSS.n9669 VSS.n9452 5.62907
R9310 VSS.n9725 VSS.n9403 5.62907
R9311 VSS.n16507 VSS.n16469 5.62907
R9312 VSS.n16564 VSS.n16420 5.62907
R9313 VSS.n16612 VSS.n16394 5.62907
R9314 VSS.n16668 VSS.n16345 5.62907
R9315 VSS.n1672 VSS.n1634 5.62907
R9316 VSS.n1729 VSS.n1585 5.62907
R9317 VSS.n16019 VSS.n1566 5.62907
R9318 VSS.n16075 VSS.n1517 5.62907
R9319 VSS.n1865 VSS.n1824 5.62907
R9320 VSS.n1931 VSS.n1769 5.62907
R9321 VSS.n2026 VSS.n2000 5.62907
R9322 VSS.n2054 VSS.n1982 5.62907
R9323 VSS.n3064 VSS.n3023 5.62907
R9324 VSS.n3130 VSS.n2968 5.62907
R9325 VSS.n3160 VSS.n2943 5.62907
R9326 VSS.n3216 VSS.n2894 5.62907
R9327 VSS.n3656 VSS.n3615 5.62907
R9328 VSS.n3722 VSS.n3560 5.62907
R9329 VSS.n3752 VSS.n3535 5.62907
R9330 VSS.n3808 VSS.n3486 5.62907
R9331 VSS.n4248 VSS.n4207 5.62907
R9332 VSS.n4314 VSS.n4152 5.62907
R9333 VSS.n4344 VSS.n4127 5.62907
R9334 VSS.n4400 VSS.n4078 5.62907
R9335 VSS.n4840 VSS.n4799 5.62907
R9336 VSS.n4906 VSS.n4744 5.62907
R9337 VSS.n4936 VSS.n4719 5.62907
R9338 VSS.n4992 VSS.n4670 5.62907
R9339 VSS.n2461 VSS.n2420 5.62907
R9340 VSS.n2527 VSS.n2365 5.62907
R9341 VSS.n2622 VSS.n2596 5.62907
R9342 VSS.n2650 VSS.n2578 5.62907
R9343 VSS.n5422 VSS.n5381 5.62907
R9344 VSS.n5488 VSS.n5326 5.62907
R9345 VSS.n5583 VSS.n5557 5.62907
R9346 VSS.n5611 VSS.n5539 5.62907
R9347 VSS.n5995 VSS.n5954 5.62907
R9348 VSS.n6061 VSS.n5899 5.62907
R9349 VSS.n6156 VSS.n6130 5.62907
R9350 VSS.n6184 VSS.n6112 5.62907
R9351 VSS.n7797 VSS.n7756 5.62907
R9352 VSS.n7863 VSS.n7701 5.62907
R9353 VSS.n7893 VSS.n7676 5.62907
R9354 VSS.n7949 VSS.n7627 5.62907
R9355 VSS.n8389 VSS.n8348 5.62907
R9356 VSS.n8455 VSS.n8293 5.62907
R9357 VSS.n8485 VSS.n8268 5.62907
R9358 VSS.n8541 VSS.n8219 5.62907
R9359 VSS.n8981 VSS.n8940 5.62907
R9360 VSS.n9047 VSS.n8885 5.62907
R9361 VSS.n9077 VSS.n8860 5.62907
R9362 VSS.n9133 VSS.n8811 5.62907
R9363 VSS.n10165 VSS.n10124 5.62907
R9364 VSS.n10231 VSS.n10069 5.62907
R9365 VSS.n10261 VSS.n10044 5.62907
R9366 VSS.n10317 VSS.n9995 5.62907
R9367 VSS.n10757 VSS.n10716 5.62907
R9368 VSS.n10823 VSS.n10661 5.62907
R9369 VSS.n10853 VSS.n10636 5.62907
R9370 VSS.n10909 VSS.n10587 5.62907
R9371 VSS.n11349 VSS.n11308 5.62907
R9372 VSS.n11415 VSS.n11253 5.62907
R9373 VSS.n11445 VSS.n11228 5.62907
R9374 VSS.n11501 VSS.n11179 5.62907
R9375 VSS.n11941 VSS.n11900 5.62907
R9376 VSS.n12007 VSS.n11845 5.62907
R9377 VSS.n12037 VSS.n11820 5.62907
R9378 VSS.n12093 VSS.n11771 5.62907
R9379 VSS.n12533 VSS.n12492 5.62907
R9380 VSS.n12599 VSS.n12437 5.62907
R9381 VSS.n12629 VSS.n12412 5.62907
R9382 VSS.n12685 VSS.n12363 5.62907
R9383 VSS.n13125 VSS.n13084 5.62907
R9384 VSS.n13191 VSS.n13029 5.62907
R9385 VSS.n13221 VSS.n13004 5.62907
R9386 VSS.n13277 VSS.n12955 5.62907
R9387 VSS.n13717 VSS.n13676 5.62907
R9388 VSS.n13783 VSS.n13621 5.62907
R9389 VSS.n13813 VSS.n13596 5.62907
R9390 VSS.n13869 VSS.n13547 5.62907
R9391 VSS.n14309 VSS.n14268 5.62907
R9392 VSS.n14375 VSS.n14213 5.62907
R9393 VSS.n14405 VSS.n14188 5.62907
R9394 VSS.n14461 VSS.n14139 5.62907
R9395 VSS.n14901 VSS.n14860 5.62907
R9396 VSS.n14967 VSS.n14805 5.62907
R9397 VSS.n14997 VSS.n14780 5.62907
R9398 VSS.n15053 VSS.n14731 5.62907
R9399 VSS.n15493 VSS.n15452 5.62907
R9400 VSS.n15559 VSS.n15397 5.62907
R9401 VSS.n15589 VSS.n15372 5.62907
R9402 VSS.n15645 VSS.n15323 5.62907
R9403 VSS.n6601 VSS.n6560 5.62907
R9404 VSS.n6667 VSS.n6505 5.62907
R9405 VSS.n6762 VSS.n6736 5.62907
R9406 VSS.n6790 VSS.n6718 5.62907
R9407 VSS.n7196 VSS.n7158 5.62907
R9408 VSS.n7253 VSS.n7109 5.62907
R9409 VSS.n7301 VSS.n7083 5.62907
R9410 VSS.n7357 VSS.n7034 5.62907
R9411 VSS.n362 VSS.n344 5.62907
R9412 VSS.n398 VSS.n329 5.62907
R9413 VSS.n18613 VSS.n181 5.62907
R9414 VSS.n18669 VSS.n132 5.62907
R9415 VSS.n585 VSS.n556 5.62907
R9416 VSS.n613 VSS.n538 5.62907
R9417 VSS.n16867 VSS.n16865 5.33568
R9418 VSS.n17123 VSS.n17106 5.33568
R9419 VSS.n17281 VSS.n17279 5.33568
R9420 VSS.n17715 VSS.n17698 5.33568
R9421 VSS.n9332 VSS.n9330 5.33568
R9422 VSS.n9765 VSS.n9748 5.33568
R9423 VSS.n16274 VSS.n16272 5.33568
R9424 VSS.n16708 VSS.n16691 5.33568
R9425 VSS.n1446 VSS.n1444 5.33568
R9426 VSS.n16115 VSS.n16098 5.33568
R9427 VSS.n2205 VSS.n2204 5.33568
R9428 VSS.n2300 VSS.n2071 5.33568
R9429 VSS.n2823 VSS.n2821 5.33568
R9430 VSS.n3256 VSS.n3239 5.33568
R9431 VSS.n3415 VSS.n3413 5.33568
R9432 VSS.n3848 VSS.n3831 5.33568
R9433 VSS.n4007 VSS.n4005 5.33568
R9434 VSS.n4440 VSS.n4423 5.33568
R9435 VSS.n4599 VSS.n4597 5.33568
R9436 VSS.n5032 VSS.n5015 5.33568
R9437 VSS.n2801 VSS.n2800 5.33568
R9438 VSS.n5265 VSS.n2667 5.33568
R9439 VSS.n8 VSS.n6 5.33568
R9440 VSS.n5838 VSS.n5628 5.33568
R9441 VSS.n6335 VSS.n6334 5.33568
R9442 VSS.n6430 VSS.n6201 5.33568
R9443 VSS.n7556 VSS.n7554 5.33568
R9444 VSS.n7989 VSS.n7972 5.33568
R9445 VSS.n8148 VSS.n8146 5.33568
R9446 VSS.n8581 VSS.n8564 5.33568
R9447 VSS.n8740 VSS.n8738 5.33568
R9448 VSS.n9173 VSS.n9156 5.33568
R9449 VSS.n9924 VSS.n9922 5.33568
R9450 VSS.n10357 VSS.n10340 5.33568
R9451 VSS.n10516 VSS.n10514 5.33568
R9452 VSS.n10949 VSS.n10932 5.33568
R9453 VSS.n11108 VSS.n11106 5.33568
R9454 VSS.n11541 VSS.n11524 5.33568
R9455 VSS.n11700 VSS.n11698 5.33568
R9456 VSS.n12133 VSS.n12116 5.33568
R9457 VSS.n12292 VSS.n12290 5.33568
R9458 VSS.n12725 VSS.n12708 5.33568
R9459 VSS.n12884 VSS.n12882 5.33568
R9460 VSS.n13317 VSS.n13300 5.33568
R9461 VSS.n13476 VSS.n13474 5.33568
R9462 VSS.n13909 VSS.n13892 5.33568
R9463 VSS.n14068 VSS.n14066 5.33568
R9464 VSS.n14501 VSS.n14484 5.33568
R9465 VSS.n14660 VSS.n14658 5.33568
R9466 VSS.n15093 VSS.n15076 5.33568
R9467 VSS.n15252 VSS.n15250 5.33568
R9468 VSS.n15685 VSS.n15668 5.33568
R9469 VSS.n6941 VSS.n6940 5.33568
R9470 VSS.n15918 VSS.n6807 5.33568
R9471 VSS.n6963 VSS.n6961 5.33568
R9472 VSS.n7397 VSS.n7380 5.33568
R9473 VSS.n61 VSS.n59 5.33568
R9474 VSS.n18709 VSS.n18692 5.33568
R9475 VSS.n18438 VSS.n18436 5.33568
R9476 VSS.n18535 VSS.n18306 5.33568
R9477 VSS.n832 VSS.n630 5.33568
R9478 VSS.n18875 VSS.n42 5.33568
R9479 VSS.n1423 VSS.n1422 5.33568
R9480 VSS.n17946 VSS.n1289 5.33568
R9481 VSS.n17529 VSS.n17528 4.84631
R9482 VSS.n17562 VSS.n17559 4.84631
R9483 VSS.n1251 VSS.n1210 4.84621
R9484 VSS.n1257 VSS.n1210 4.84621
R9485 VSS.n1116 VSS.n1077 4.84621
R9486 VSS.n1122 VSS.n1077 4.84621
R9487 VSS.n17055 VSS.n16970 4.84621
R9488 VSS.n17055 VSS.n16971 4.84621
R9489 VSS.n17555 VSS.n17460 4.84621
R9490 VSS.n17556 VSS.n17555 4.84621
R9491 VSS.n17647 VSS.n17384 4.84621
R9492 VSS.n17647 VSS.n17385 4.84621
R9493 VSS.n18268 VSS.n18227 4.84621
R9494 VSS.n18274 VSS.n18227 4.84621
R9495 VSS.n18132 VSS.n252 4.84621
R9496 VSS.n18133 VSS.n18132 4.84621
R9497 VSS.n9697 VSS.n9434 4.84621
R9498 VSS.n9697 VSS.n9435 4.84621
R9499 VSS.n9605 VSS.n9510 4.84621
R9500 VSS.n9606 VSS.n9605 4.84621
R9501 VSS.n16640 VSS.n16376 4.84621
R9502 VSS.n16640 VSS.n16377 4.84621
R9503 VSS.n16535 VSS.n16453 4.84621
R9504 VSS.n16535 VSS.n16454 4.84621
R9505 VSS.n16047 VSS.n1548 4.84621
R9506 VSS.n16047 VSS.n1549 4.84621
R9507 VSS.n1700 VSS.n1618 4.84621
R9508 VSS.n1700 VSS.n1619 4.84621
R9509 VSS.n2033 VSS.n1992 4.84621
R9510 VSS.n2039 VSS.n1992 4.84621
R9511 VSS.n1897 VSS.n1802 4.84621
R9512 VSS.n1898 VSS.n1897 4.84621
R9513 VSS.n3188 VSS.n2925 4.84621
R9514 VSS.n3188 VSS.n2926 4.84621
R9515 VSS.n3096 VSS.n3001 4.84621
R9516 VSS.n3097 VSS.n3096 4.84621
R9517 VSS.n3780 VSS.n3517 4.84621
R9518 VSS.n3780 VSS.n3518 4.84621
R9519 VSS.n3688 VSS.n3593 4.84621
R9520 VSS.n3689 VSS.n3688 4.84621
R9521 VSS.n4372 VSS.n4109 4.84621
R9522 VSS.n4372 VSS.n4110 4.84621
R9523 VSS.n4280 VSS.n4185 4.84621
R9524 VSS.n4281 VSS.n4280 4.84621
R9525 VSS.n4964 VSS.n4701 4.84621
R9526 VSS.n4964 VSS.n4702 4.84621
R9527 VSS.n4872 VSS.n4777 4.84621
R9528 VSS.n4873 VSS.n4872 4.84621
R9529 VSS.n2629 VSS.n2588 4.84621
R9530 VSS.n2635 VSS.n2588 4.84621
R9531 VSS.n2493 VSS.n2398 4.84621
R9532 VSS.n2494 VSS.n2493 4.84621
R9533 VSS.n5590 VSS.n5549 4.84621
R9534 VSS.n5596 VSS.n5549 4.84621
R9535 VSS.n5454 VSS.n5359 4.84621
R9536 VSS.n5455 VSS.n5454 4.84621
R9537 VSS.n6163 VSS.n6122 4.84621
R9538 VSS.n6169 VSS.n6122 4.84621
R9539 VSS.n6027 VSS.n5932 4.84621
R9540 VSS.n6028 VSS.n6027 4.84621
R9541 VSS.n7921 VSS.n7658 4.84621
R9542 VSS.n7921 VSS.n7659 4.84621
R9543 VSS.n7829 VSS.n7734 4.84621
R9544 VSS.n7830 VSS.n7829 4.84621
R9545 VSS.n8513 VSS.n8250 4.84621
R9546 VSS.n8513 VSS.n8251 4.84621
R9547 VSS.n8421 VSS.n8326 4.84621
R9548 VSS.n8422 VSS.n8421 4.84621
R9549 VSS.n9105 VSS.n8842 4.84621
R9550 VSS.n9105 VSS.n8843 4.84621
R9551 VSS.n9013 VSS.n8918 4.84621
R9552 VSS.n9014 VSS.n9013 4.84621
R9553 VSS.n10289 VSS.n10026 4.84621
R9554 VSS.n10289 VSS.n10027 4.84621
R9555 VSS.n10197 VSS.n10102 4.84621
R9556 VSS.n10198 VSS.n10197 4.84621
R9557 VSS.n10881 VSS.n10618 4.84621
R9558 VSS.n10881 VSS.n10619 4.84621
R9559 VSS.n10789 VSS.n10694 4.84621
R9560 VSS.n10790 VSS.n10789 4.84621
R9561 VSS.n11473 VSS.n11210 4.84621
R9562 VSS.n11473 VSS.n11211 4.84621
R9563 VSS.n11381 VSS.n11286 4.84621
R9564 VSS.n11382 VSS.n11381 4.84621
R9565 VSS.n12065 VSS.n11802 4.84621
R9566 VSS.n12065 VSS.n11803 4.84621
R9567 VSS.n11973 VSS.n11878 4.84621
R9568 VSS.n11974 VSS.n11973 4.84621
R9569 VSS.n12657 VSS.n12394 4.84621
R9570 VSS.n12657 VSS.n12395 4.84621
R9571 VSS.n12565 VSS.n12470 4.84621
R9572 VSS.n12566 VSS.n12565 4.84621
R9573 VSS.n13249 VSS.n12986 4.84621
R9574 VSS.n13249 VSS.n12987 4.84621
R9575 VSS.n13157 VSS.n13062 4.84621
R9576 VSS.n13158 VSS.n13157 4.84621
R9577 VSS.n13841 VSS.n13578 4.84621
R9578 VSS.n13841 VSS.n13579 4.84621
R9579 VSS.n13749 VSS.n13654 4.84621
R9580 VSS.n13750 VSS.n13749 4.84621
R9581 VSS.n14433 VSS.n14170 4.84621
R9582 VSS.n14433 VSS.n14171 4.84621
R9583 VSS.n14341 VSS.n14246 4.84621
R9584 VSS.n14342 VSS.n14341 4.84621
R9585 VSS.n15025 VSS.n14762 4.84621
R9586 VSS.n15025 VSS.n14763 4.84621
R9587 VSS.n14933 VSS.n14838 4.84621
R9588 VSS.n14934 VSS.n14933 4.84621
R9589 VSS.n15617 VSS.n15354 4.84621
R9590 VSS.n15617 VSS.n15355 4.84621
R9591 VSS.n15525 VSS.n15430 4.84621
R9592 VSS.n15526 VSS.n15525 4.84621
R9593 VSS.n6769 VSS.n6728 4.84621
R9594 VSS.n6775 VSS.n6728 4.84621
R9595 VSS.n6633 VSS.n6538 4.84621
R9596 VSS.n6634 VSS.n6633 4.84621
R9597 VSS.n7329 VSS.n7065 4.84621
R9598 VSS.n7329 VSS.n7066 4.84621
R9599 VSS.n7224 VSS.n7142 4.84621
R9600 VSS.n7224 VSS.n7143 4.84621
R9601 VSS.n18641 VSS.n163 4.84621
R9602 VSS.n18641 VSS.n164 4.84621
R9603 VSS.n379 VSS.n377 4.84621
R9604 VSS.n380 VSS.n379 4.84621
R9605 VSS.n592 VSS.n548 4.84621
R9606 VSS.n598 VSS.n548 4.84621
R9607 VSS.n935 VSS.n896 4.84621
R9608 VSS.n941 VSS.n896 4.84621
R9609 VSS.n1228 VSS.n1222 4.6505
R9610 VSS.n1095 VSS.n1089 4.6505
R9611 VSS.n17011 VSS.n16990 4.6505
R9612 VSS.n17505 VSS.n17483 4.6505
R9613 VSS.n17603 VSS.n17404 4.6505
R9614 VSS.n18245 VSS.n18239 4.6505
R9615 VSS.n18082 VSS.n275 4.6505
R9616 VSS.n9653 VSS.n9454 4.6505
R9617 VSS.n9555 VSS.n9533 4.6505
R9618 VSS.n16596 VSS.n16396 4.6505
R9619 VSS.n16491 VSS.n16471 4.6505
R9620 VSS.n16003 VSS.n1568 4.6505
R9621 VSS.n1656 VSS.n1636 4.6505
R9622 VSS.n2010 VSS.n2004 4.6505
R9623 VSS.n1847 VSS.n1825 4.6505
R9624 VSS.n3144 VSS.n2945 4.6505
R9625 VSS.n3046 VSS.n3024 4.6505
R9626 VSS.n3736 VSS.n3537 4.6505
R9627 VSS.n3638 VSS.n3616 4.6505
R9628 VSS.n4328 VSS.n4129 4.6505
R9629 VSS.n4230 VSS.n4208 4.6505
R9630 VSS.n4920 VSS.n4721 4.6505
R9631 VSS.n4822 VSS.n4800 4.6505
R9632 VSS.n2606 VSS.n2600 4.6505
R9633 VSS.n2443 VSS.n2421 4.6505
R9634 VSS.n5567 VSS.n5561 4.6505
R9635 VSS.n5404 VSS.n5382 4.6505
R9636 VSS.n6140 VSS.n6134 4.6505
R9637 VSS.n5977 VSS.n5955 4.6505
R9638 VSS.n7877 VSS.n7678 4.6505
R9639 VSS.n7779 VSS.n7757 4.6505
R9640 VSS.n8469 VSS.n8270 4.6505
R9641 VSS.n8371 VSS.n8349 4.6505
R9642 VSS.n9061 VSS.n8862 4.6505
R9643 VSS.n8963 VSS.n8941 4.6505
R9644 VSS.n10245 VSS.n10046 4.6505
R9645 VSS.n10147 VSS.n10125 4.6505
R9646 VSS.n10837 VSS.n10638 4.6505
R9647 VSS.n10739 VSS.n10717 4.6505
R9648 VSS.n11429 VSS.n11230 4.6505
R9649 VSS.n11331 VSS.n11309 4.6505
R9650 VSS.n12021 VSS.n11822 4.6505
R9651 VSS.n11923 VSS.n11901 4.6505
R9652 VSS.n12613 VSS.n12414 4.6505
R9653 VSS.n12515 VSS.n12493 4.6505
R9654 VSS.n13205 VSS.n13006 4.6505
R9655 VSS.n13107 VSS.n13085 4.6505
R9656 VSS.n13797 VSS.n13598 4.6505
R9657 VSS.n13699 VSS.n13677 4.6505
R9658 VSS.n14389 VSS.n14190 4.6505
R9659 VSS.n14291 VSS.n14269 4.6505
R9660 VSS.n14981 VSS.n14782 4.6505
R9661 VSS.n14883 VSS.n14861 4.6505
R9662 VSS.n15573 VSS.n15374 4.6505
R9663 VSS.n15475 VSS.n15453 4.6505
R9664 VSS.n6746 VSS.n6740 4.6505
R9665 VSS.n6583 VSS.n6561 4.6505
R9666 VSS.n7285 VSS.n7085 4.6505
R9667 VSS.n7180 VSS.n7160 4.6505
R9668 VSS.n18597 VSS.n183 4.6505
R9669 VSS.n356 VSS.n355 4.6505
R9670 VSS.n569 VSS.n565 4.6505
R9671 VSS.n914 VSS.n908 4.6505
R9672 VSS.n17163 VSS.n16916 4.61769
R9673 VSS.n17238 VSS.n16880 4.61769
R9674 VSS.n17755 VSS.n17330 4.61769
R9675 VSS.n17830 VSS.n17294 4.61769
R9676 VSS.n18368 VSS.n18362 4.61769
R9677 VSS.n18452 VSS.n18440 4.61769
R9678 VSS.n9805 VSS.n9380 4.61769
R9679 VSS.n9880 VSS.n9344 4.61769
R9680 VSS.n16748 VSS.n16322 4.61769
R9681 VSS.n16823 VSS.n16286 4.61769
R9682 VSS.n16155 VSS.n1494 4.61769
R9683 VSS.n16230 VSS.n1458 4.61769
R9684 VSS.n2282 VSS.n2104 4.61769
R9685 VSS.n2195 VSS.n2175 4.61769
R9686 VSS.n3296 VSS.n2871 4.61769
R9687 VSS.n3371 VSS.n2835 4.61769
R9688 VSS.n3888 VSS.n3463 4.61769
R9689 VSS.n3963 VSS.n3427 4.61769
R9690 VSS.n4480 VSS.n4055 4.61769
R9691 VSS.n4555 VSS.n4019 4.61769
R9692 VSS.n5072 VSS.n4647 4.61769
R9693 VSS.n5147 VSS.n4611 4.61769
R9694 VSS.n5247 VSS.n2700 4.61769
R9695 VSS.n2791 VSS.n2771 4.61769
R9696 VSS.n5820 VSS.n5661 4.61769
R9697 VSS.n5765 VSS.n5745 4.61769
R9698 VSS.n6412 VSS.n6234 4.61769
R9699 VSS.n6325 VSS.n6305 4.61769
R9700 VSS.n8029 VSS.n7604 4.61769
R9701 VSS.n8104 VSS.n7568 4.61769
R9702 VSS.n8621 VSS.n8196 4.61769
R9703 VSS.n8696 VSS.n8160 4.61769
R9704 VSS.n9213 VSS.n8788 4.61769
R9705 VSS.n9288 VSS.n8752 4.61769
R9706 VSS.n10397 VSS.n9972 4.61769
R9707 VSS.n10472 VSS.n9936 4.61769
R9708 VSS.n10989 VSS.n10564 4.61769
R9709 VSS.n11064 VSS.n10528 4.61769
R9710 VSS.n11581 VSS.n11156 4.61769
R9711 VSS.n11656 VSS.n11120 4.61769
R9712 VSS.n12173 VSS.n11748 4.61769
R9713 VSS.n12248 VSS.n11712 4.61769
R9714 VSS.n12765 VSS.n12340 4.61769
R9715 VSS.n12840 VSS.n12304 4.61769
R9716 VSS.n13357 VSS.n12932 4.61769
R9717 VSS.n13432 VSS.n12896 4.61769
R9718 VSS.n13949 VSS.n13524 4.61769
R9719 VSS.n14024 VSS.n13488 4.61769
R9720 VSS.n14541 VSS.n14116 4.61769
R9721 VSS.n14616 VSS.n14080 4.61769
R9722 VSS.n15133 VSS.n14708 4.61769
R9723 VSS.n15208 VSS.n14672 4.61769
R9724 VSS.n15725 VSS.n15300 4.61769
R9725 VSS.n15800 VSS.n15264 4.61769
R9726 VSS.n15900 VSS.n6840 4.61769
R9727 VSS.n6931 VSS.n6911 4.61769
R9728 VSS.n7437 VSS.n7011 4.61769
R9729 VSS.n7512 VSS.n6975 4.61769
R9730 VSS.n18749 VSS.n109 4.61769
R9731 VSS.n18824 VSS.n73 4.61769
R9732 VSS.n814 VSS.n663 4.61769
R9733 VSS.n761 VSS.n744 4.61769
R9734 VSS.n17928 VSS.n1322 4.61769
R9735 VSS.n1413 VSS.n1393 4.61769
R9736 VSS.n1278 VSS.n1277 4.5005
R9737 VSS.n1281 VSS.n1280 4.5005
R9738 VSS.n1264 VSS.n1263 4.5005
R9739 VSS.n1239 VSS.n1238 4.5005
R9740 VSS.n1230 VSS.n1229 4.5005
R9741 VSS.n1231 VSS.n1223 4.5005
R9742 VSS.n1227 VSS.n1224 4.5005
R9743 VSS.n1188 VSS.n1186 4.5005
R9744 VSS.n17962 VSS.n17961 4.5005
R9745 VSS.n17969 VSS.n1178 4.5005
R9746 VSS.n17976 VSS.n17975 4.5005
R9747 VSS.n17977 VSS.n1170 4.5005
R9748 VSS.n1235 VSS.n1167 4.5005
R9749 VSS.n17984 VSS.n17983 4.5005
R9750 VSS.n17968 VSS.n17967 4.5005
R9751 VSS.n1279 VSS.n1203 4.5005
R9752 VSS.n17992 VSS.n17991 4.5005
R9753 VSS.n1276 VSS.n1204 4.5005
R9754 VSS.n1276 VSS.n1275 4.5005
R9755 VSS.n1237 VSS.n1236 4.5005
R9756 VSS.n1236 VSS.n1214 4.5005
R9757 VSS.n1233 VSS.n1232 4.5005
R9758 VSS.n1266 VSS.n1265 4.5005
R9759 VSS.n1266 VSS.n1259 4.5005
R9760 VSS.n17954 VSS.n1196 4.5005
R9761 VSS.n17954 VSS.n17953 4.5005
R9762 VSS.n1144 VSS.n1143 4.5005
R9763 VSS.n1147 VSS.n1146 4.5005
R9764 VSS.n1129 VSS.n1128 4.5005
R9765 VSS.n1104 VSS.n1032 4.5005
R9766 VSS.n1097 VSS.n1096 4.5005
R9767 VSS.n1098 VSS.n1090 4.5005
R9768 VSS.n18041 VSS.n18040 4.5005
R9769 VSS.n1094 VSS.n1091 4.5005
R9770 VSS.n1142 VSS.n1070 4.5005
R9771 VSS.n1142 VSS.n1141 4.5005
R9772 VSS.n1054 VSS.n1052 4.5005
R9773 VSS.n18011 VSS.n18010 4.5005
R9774 VSS.n18018 VSS.n1044 4.5005
R9775 VSS.n18025 VSS.n18024 4.5005
R9776 VSS.n1076 VSS.n1040 4.5005
R9777 VSS.n18026 VSS.n1035 4.5005
R9778 VSS.n1103 VSS.n1102 4.5005
R9779 VSS.n1103 VSS.n1081 4.5005
R9780 VSS.n18033 VSS.n18032 4.5005
R9781 VSS.n1100 VSS.n1099 4.5005
R9782 VSS.n18017 VSS.n18016 4.5005
R9783 VSS.n1131 VSS.n1130 4.5005
R9784 VSS.n1131 VSS.n1124 4.5005
R9785 VSS.n1145 VSS.n1069 4.5005
R9786 VSS.n18003 VSS.n1062 4.5005
R9787 VSS.n18003 VSS.n18002 4.5005
R9788 VSS.n17255 VSS.n17254 4.5005
R9789 VSS.n17196 VSS.n16900 4.5005
R9790 VSS.n17159 VSS.n17158 4.5005
R9791 VSS.n17109 VSS.n17107 4.5005
R9792 VSS.n17138 VSS.n17137 4.5005
R9793 VSS.n17149 VSS.n17148 4.5005
R9794 VSS.n17150 VSS.n17149 4.5005
R9795 VSS.n17183 VSS.n17182 4.5005
R9796 VSS.n17156 VSS.n17155 4.5005
R9797 VSS.n16909 VSS.n16908 4.5005
R9798 VSS.n16918 VSS.n16909 4.5005
R9799 VSS.n17249 VSS.n17248 4.5005
R9800 VSS.n17223 VSS.n16889 4.5005
R9801 VSS.n17223 VSS.n16883 4.5005
R9802 VSS.n17230 VSS.n16885 4.5005
R9803 VSS.n17201 VSS.n17197 4.5005
R9804 VSS.n17201 VSS.n17200 4.5005
R9805 VSS.n17204 VSS.n17195 4.5005
R9806 VSS.n17188 VSS.n17187 4.5005
R9807 VSS.n17187 VSS.n16895 4.5005
R9808 VSS.n17253 VSS.n16873 4.5005
R9809 VSS.n16877 VSS.n16871 4.5005
R9810 VSS.n16871 VSS.n16870 4.5005
R9811 VSS.n17211 VSS.n17210 4.5005
R9812 VSS.n17212 VSS.n17211 4.5005
R9813 VSS.n16886 VSS.n16884 4.5005
R9814 VSS.n17268 VSS.n17267 4.5005
R9815 VSS.n17140 VSS.n17139 4.5005
R9816 VSS.n17141 VSS.n16929 4.5005
R9817 VSS.n16948 VSS.n16943 4.5005
R9818 VSS.n17098 VSS.n17097 4.5005
R9819 VSS.n17075 VSS.n16958 4.5005
R9820 VSS.n16986 VSS.n16984 4.5005
R9821 VSS.n17014 VSS.n17012 4.5005
R9822 VSS.n17013 VSS.n16991 4.5005
R9823 VSS.n17016 VSS.n17015 4.5005
R9824 VSS.n17074 VSS.n17073 4.5005
R9825 VSS.n16960 VSS.n16947 4.5005
R9826 VSS.n17064 VSS.n17063 4.5005
R9827 VSS.n16969 VSS.n16967 4.5005
R9828 VSS.n16981 VSS.n16980 4.5005
R9829 VSS.n17036 VSS.n17035 4.5005
R9830 VSS.n16993 VSS.n16983 4.5005
R9831 VSS.n17065 VSS.n16962 4.5005
R9832 VSS.n17096 VSS.n16942 4.5005
R9833 VSS.n17010 VSS.n17009 4.5005
R9834 VSS.n16950 VSS.n16949 4.5005
R9835 VSS.n17085 VSS.n16950 4.5005
R9836 VSS.n16979 VSS.n16977 4.5005
R9837 VSS.n16977 VSS.n16976 4.5005
R9838 VSS.n17025 VSS.n16992 4.5005
R9839 VSS.n17077 VSS.n17076 4.5005
R9840 VSS.n17077 VSS.n16956 4.5005
R9841 VSS.n17132 VSS.n17131 4.5005
R9842 VSS.n17131 VSS.n17130 4.5005
R9843 VSS.n17584 VSS.n17431 4.5005
R9844 VSS.n17583 VSS.n17582 4.5005
R9845 VSS.n17453 VSS.n17452 4.5005
R9846 VSS.n17535 VSS.n17534 4.5005
R9847 VSS.n17508 VSS.n17506 4.5005
R9848 VSS.n17507 VSS.n17484 4.5005
R9849 VSS.n17504 VSS.n17503 4.5005
R9850 VSS.n17510 VSS.n17509 4.5005
R9851 VSS.n17586 VSS.n17585 4.5005
R9852 VSS.n17586 VSS.n17429 4.5005
R9853 VSS.n17442 VSS.n17441 4.5005
R9854 VSS.n17573 VSS.n17572 4.5005
R9855 VSS.n17465 VSS.n17464 4.5005
R9856 VSS.n17544 VSS.n17543 4.5005
R9857 VSS.n17554 VSS.n17462 4.5005
R9858 VSS.n17542 VSS.n17541 4.5005
R9859 VSS.n17533 VSS.n17472 4.5005
R9860 VSS.n17533 VSS.n17532 4.5005
R9861 VSS.n17487 VSS.n17471 4.5005
R9862 VSS.n17519 VSS.n17485 4.5005
R9863 VSS.n17446 VSS.n17444 4.5005
R9864 VSS.n17451 VSS.n17447 4.5005
R9865 VSS.n17449 VSS.n17447 4.5005
R9866 VSS.n17581 VSS.n17433 4.5005
R9867 VSS.n17598 VSS.n17597 4.5005
R9868 VSS.n17597 VSS.n17596 4.5005
R9869 VSS.n17847 VSS.n17846 4.5005
R9870 VSS.n17788 VSS.n17314 4.5005
R9871 VSS.n17751 VSS.n17750 4.5005
R9872 VSS.n17701 VSS.n17699 4.5005
R9873 VSS.n17730 VSS.n17729 4.5005
R9874 VSS.n17741 VSS.n17740 4.5005
R9875 VSS.n17742 VSS.n17741 4.5005
R9876 VSS.n17775 VSS.n17774 4.5005
R9877 VSS.n17748 VSS.n17747 4.5005
R9878 VSS.n17323 VSS.n17322 4.5005
R9879 VSS.n17332 VSS.n17323 4.5005
R9880 VSS.n17841 VSS.n17840 4.5005
R9881 VSS.n17815 VSS.n17303 4.5005
R9882 VSS.n17815 VSS.n17297 4.5005
R9883 VSS.n17822 VSS.n17299 4.5005
R9884 VSS.n17793 VSS.n17789 4.5005
R9885 VSS.n17793 VSS.n17792 4.5005
R9886 VSS.n17796 VSS.n17787 4.5005
R9887 VSS.n17780 VSS.n17779 4.5005
R9888 VSS.n17779 VSS.n17309 4.5005
R9889 VSS.n17845 VSS.n17287 4.5005
R9890 VSS.n17291 VSS.n17285 4.5005
R9891 VSS.n17285 VSS.n17284 4.5005
R9892 VSS.n17803 VSS.n17802 4.5005
R9893 VSS.n17804 VSS.n17803 4.5005
R9894 VSS.n17300 VSS.n17298 4.5005
R9895 VSS.n17860 VSS.n17859 4.5005
R9896 VSS.n17732 VSS.n17731 4.5005
R9897 VSS.n17733 VSS.n17343 4.5005
R9898 VSS.n17362 VSS.n17357 4.5005
R9899 VSS.n17690 VSS.n17689 4.5005
R9900 VSS.n17667 VSS.n17372 4.5005
R9901 VSS.n17400 VSS.n17398 4.5005
R9902 VSS.n17606 VSS.n17604 4.5005
R9903 VSS.n17605 VSS.n17405 4.5005
R9904 VSS.n17608 VSS.n17607 4.5005
R9905 VSS.n17666 VSS.n17665 4.5005
R9906 VSS.n17374 VSS.n17361 4.5005
R9907 VSS.n17656 VSS.n17655 4.5005
R9908 VSS.n17383 VSS.n17381 4.5005
R9909 VSS.n17395 VSS.n17394 4.5005
R9910 VSS.n17628 VSS.n17627 4.5005
R9911 VSS.n17407 VSS.n17397 4.5005
R9912 VSS.n17657 VSS.n17376 4.5005
R9913 VSS.n17688 VSS.n17356 4.5005
R9914 VSS.n17602 VSS.n17601 4.5005
R9915 VSS.n17364 VSS.n17363 4.5005
R9916 VSS.n17677 VSS.n17364 4.5005
R9917 VSS.n17393 VSS.n17391 4.5005
R9918 VSS.n17391 VSS.n17390 4.5005
R9919 VSS.n17617 VSS.n17406 4.5005
R9920 VSS.n17669 VSS.n17668 4.5005
R9921 VSS.n17669 VSS.n17370 4.5005
R9922 VSS.n17724 VSS.n17723 4.5005
R9923 VSS.n17723 VSS.n17722 4.5005
R9924 VSS.n18295 VSS.n18294 4.5005
R9925 VSS.n18298 VSS.n18297 4.5005
R9926 VSS.n18281 VSS.n18280 4.5005
R9927 VSS.n18256 VSS.n18255 4.5005
R9928 VSS.n18247 VSS.n18246 4.5005
R9929 VSS.n18248 VSS.n18240 4.5005
R9930 VSS.n18581 VSS.n18580 4.5005
R9931 VSS.n18244 VSS.n18241 4.5005
R9932 VSS.n18293 VSS.n18221 4.5005
R9933 VSS.n18293 VSS.n18292 4.5005
R9934 VSS.n18205 VSS.n18203 4.5005
R9935 VSS.n18551 VSS.n18550 4.5005
R9936 VSS.n18558 VSS.n18195 4.5005
R9937 VSS.n18565 VSS.n18564 4.5005
R9938 VSS.n18566 VSS.n18187 4.5005
R9939 VSS.n18252 VSS.n18184 4.5005
R9940 VSS.n18254 VSS.n18253 4.5005
R9941 VSS.n18253 VSS.n18231 4.5005
R9942 VSS.n18573 VSS.n18572 4.5005
R9943 VSS.n18250 VSS.n18249 4.5005
R9944 VSS.n18557 VSS.n18556 4.5005
R9945 VSS.n18283 VSS.n18282 4.5005
R9946 VSS.n18283 VSS.n18276 4.5005
R9947 VSS.n18296 VSS.n18220 4.5005
R9948 VSS.n18543 VSS.n18213 4.5005
R9949 VSS.n18543 VSS.n18542 4.5005
R9950 VSS.n18475 VSS.n18474 4.5005
R9951 VSS.n18397 VSS.n18394 4.5005
R9952 VSS.n18514 VSS.n18513 4.5005
R9953 VSS.n18324 VSS.n18307 4.5005
R9954 VSS.n18332 VSS.n18331 4.5005
R9955 VSS.n18525 VSS.n18524 4.5005
R9956 VSS.n18525 VSS.n18313 4.5005
R9957 VSS.n18377 VSS.n18374 4.5005
R9958 VSS.n18517 VSS.n18338 4.5005
R9959 VSS.n18512 VSS.n18341 4.5005
R9960 VSS.n18512 VSS.n18511 4.5005
R9961 VSS.n18433 VSS.n18431 4.5005
R9962 VSS.n18391 VSS.n18389 4.5005
R9963 VSS.n18441 VSS.n18389 4.5005
R9964 VSS.n18418 VSS.n18416 4.5005
R9965 VSS.n18406 VSS.n18395 4.5005
R9966 VSS.n18406 VSS.n18405 4.5005
R9967 VSS.n18411 VSS.n18388 4.5005
R9968 VSS.n18501 VSS.n18500 4.5005
R9969 VSS.n18500 VSS.n18499 4.5005
R9970 VSS.n18473 VSS.n18425 4.5005
R9971 VSS.n18478 VSS.n18477 4.5005
R9972 VSS.n18479 VSS.n18478 4.5005
R9973 VSS.n18401 VSS.n18400 4.5005
R9974 VSS.n18401 VSS.n18358 4.5005
R9975 VSS.n18444 VSS.n18443 4.5005
R9976 VSS.n18464 VSS.n18463 4.5005
R9977 VSS.n18320 VSS.n18314 4.5005
R9978 VSS.n18333 VSS.n18321 4.5005
R9979 VSS.n18161 VSS.n223 4.5005
R9980 VSS.n18160 VSS.n18159 4.5005
R9981 VSS.n245 VSS.n244 4.5005
R9982 VSS.n18112 VSS.n18111 4.5005
R9983 VSS.n18085 VSS.n18083 4.5005
R9984 VSS.n18084 VSS.n276 4.5005
R9985 VSS.n18087 VSS.n18086 4.5005
R9986 VSS.n234 VSS.n233 4.5005
R9987 VSS.n18150 VSS.n18149 4.5005
R9988 VSS.n257 VSS.n256 4.5005
R9989 VSS.n18121 VSS.n18120 4.5005
R9990 VSS.n18119 VSS.n18118 4.5005
R9991 VSS.n279 VSS.n263 4.5005
R9992 VSS.n238 VSS.n236 4.5005
R9993 VSS.n18158 VSS.n225 4.5005
R9994 VSS.n18081 VSS.n18080 4.5005
R9995 VSS.n18163 VSS.n18162 4.5005
R9996 VSS.n18163 VSS.n221 4.5005
R9997 VSS.n18131 VSS.n254 4.5005
R9998 VSS.n18110 VSS.n264 4.5005
R9999 VSS.n18110 VSS.n18109 4.5005
R10000 VSS.n18096 VSS.n277 4.5005
R10001 VSS.n243 VSS.n239 4.5005
R10002 VSS.n241 VSS.n239 4.5005
R10003 VSS.n18175 VSS.n18174 4.5005
R10004 VSS.n18174 VSS.n18173 4.5005
R10005 VSS.n9412 VSS.n9407 4.5005
R10006 VSS.n9740 VSS.n9739 4.5005
R10007 VSS.n9717 VSS.n9422 4.5005
R10008 VSS.n9450 VSS.n9448 4.5005
R10009 VSS.n9656 VSS.n9654 4.5005
R10010 VSS.n9655 VSS.n9455 4.5005
R10011 VSS.n9658 VSS.n9657 4.5005
R10012 VSS.n9716 VSS.n9715 4.5005
R10013 VSS.n9424 VSS.n9411 4.5005
R10014 VSS.n9706 VSS.n9705 4.5005
R10015 VSS.n9433 VSS.n9431 4.5005
R10016 VSS.n9445 VSS.n9444 4.5005
R10017 VSS.n9678 VSS.n9677 4.5005
R10018 VSS.n9457 VSS.n9447 4.5005
R10019 VSS.n9707 VSS.n9426 4.5005
R10020 VSS.n9738 VSS.n9406 4.5005
R10021 VSS.n9652 VSS.n9651 4.5005
R10022 VSS.n9414 VSS.n9413 4.5005
R10023 VSS.n9727 VSS.n9414 4.5005
R10024 VSS.n9443 VSS.n9441 4.5005
R10025 VSS.n9441 VSS.n9440 4.5005
R10026 VSS.n9667 VSS.n9456 4.5005
R10027 VSS.n9719 VSS.n9718 4.5005
R10028 VSS.n9719 VSS.n9420 4.5005
R10029 VSS.n9774 VSS.n9773 4.5005
R10030 VSS.n9773 VSS.n9772 4.5005
R10031 VSS.n9897 VSS.n9337 4.5005
R10032 VSS.n9838 VSS.n9364 4.5005
R10033 VSS.n9801 VSS.n9800 4.5005
R10034 VSS.n9751 VSS.n9749 4.5005
R10035 VSS.n9780 VSS.n9779 4.5005
R10036 VSS.n9791 VSS.n9790 4.5005
R10037 VSS.n9792 VSS.n9791 4.5005
R10038 VSS.n9825 VSS.n9824 4.5005
R10039 VSS.n9798 VSS.n9797 4.5005
R10040 VSS.n9373 VSS.n9372 4.5005
R10041 VSS.n9382 VSS.n9373 4.5005
R10042 VSS.n9892 VSS.n9891 4.5005
R10043 VSS.n9865 VSS.n9353 4.5005
R10044 VSS.n9865 VSS.n9347 4.5005
R10045 VSS.n9872 VSS.n9349 4.5005
R10046 VSS.n9843 VSS.n9839 4.5005
R10047 VSS.n9843 VSS.n9842 4.5005
R10048 VSS.n9846 VSS.n9837 4.5005
R10049 VSS.n9830 VSS.n9829 4.5005
R10050 VSS.n9829 VSS.n9359 4.5005
R10051 VSS.n9896 VSS.n9895 4.5005
R10052 VSS.n9338 VSS.n9336 4.5005
R10053 VSS.n9336 VSS.n9335 4.5005
R10054 VSS.n9853 VSS.n9852 4.5005
R10055 VSS.n9854 VSS.n9853 4.5005
R10056 VSS.n9350 VSS.n9348 4.5005
R10057 VSS.n9911 VSS.n9910 4.5005
R10058 VSS.n9782 VSS.n9781 4.5005
R10059 VSS.n9783 VSS.n9393 4.5005
R10060 VSS.n9634 VSS.n9481 4.5005
R10061 VSS.n9633 VSS.n9632 4.5005
R10062 VSS.n9558 VSS.n9556 4.5005
R10063 VSS.n9557 VSS.n9534 4.5005
R10064 VSS.n9592 VSS.n9591 4.5005
R10065 VSS.n9537 VSS.n9521 4.5005
R10066 VSS.n9560 VSS.n9559 4.5005
R10067 VSS.n9492 VSS.n9491 4.5005
R10068 VSS.n9623 VSS.n9622 4.5005
R10069 VSS.n9515 VSS.n9514 4.5005
R10070 VSS.n9594 VSS.n9593 4.5005
R10071 VSS.n9496 VSS.n9494 4.5005
R10072 VSS.n9503 VSS.n9502 4.5005
R10073 VSS.n9631 VSS.n9483 4.5005
R10074 VSS.n9585 VSS.n9584 4.5005
R10075 VSS.n9583 VSS.n9522 4.5005
R10076 VSS.n9583 VSS.n9582 4.5005
R10077 VSS.n9569 VSS.n9535 4.5005
R10078 VSS.n9554 VSS.n9553 4.5005
R10079 VSS.n9636 VSS.n9635 4.5005
R10080 VSS.n9636 VSS.n9479 4.5005
R10081 VSS.n9604 VSS.n9512 4.5005
R10082 VSS.n9501 VSS.n9497 4.5005
R10083 VSS.n9499 VSS.n9497 4.5005
R10084 VSS.n9648 VSS.n9647 4.5005
R10085 VSS.n9647 VSS.n9646 4.5005
R10086 VSS.n16354 VSS.n16349 4.5005
R10087 VSS.n16683 VSS.n16682 4.5005
R10088 VSS.n16660 VSS.n16364 4.5005
R10089 VSS.n16392 VSS.n16390 4.5005
R10090 VSS.n16599 VSS.n16597 4.5005
R10091 VSS.n16598 VSS.n16397 4.5005
R10092 VSS.n16601 VSS.n16600 4.5005
R10093 VSS.n16659 VSS.n16658 4.5005
R10094 VSS.n16366 VSS.n16353 4.5005
R10095 VSS.n16649 VSS.n16648 4.5005
R10096 VSS.n16375 VSS.n16373 4.5005
R10097 VSS.n16387 VSS.n16386 4.5005
R10098 VSS.n16621 VSS.n16620 4.5005
R10099 VSS.n16399 VSS.n16389 4.5005
R10100 VSS.n16650 VSS.n16368 4.5005
R10101 VSS.n16681 VSS.n16348 4.5005
R10102 VSS.n16595 VSS.n16594 4.5005
R10103 VSS.n16356 VSS.n16355 4.5005
R10104 VSS.n16670 VSS.n16356 4.5005
R10105 VSS.n16385 VSS.n16383 4.5005
R10106 VSS.n16383 VSS.n16382 4.5005
R10107 VSS.n16610 VSS.n16398 4.5005
R10108 VSS.n16662 VSS.n16661 4.5005
R10109 VSS.n16662 VSS.n16362 4.5005
R10110 VSS.n16717 VSS.n16716 4.5005
R10111 VSS.n16716 VSS.n16715 4.5005
R10112 VSS.n16840 VSS.n16279 4.5005
R10113 VSS.n16781 VSS.n16306 4.5005
R10114 VSS.n16744 VSS.n16743 4.5005
R10115 VSS.n16694 VSS.n16692 4.5005
R10116 VSS.n16723 VSS.n16722 4.5005
R10117 VSS.n16734 VSS.n16733 4.5005
R10118 VSS.n16735 VSS.n16734 4.5005
R10119 VSS.n16768 VSS.n16767 4.5005
R10120 VSS.n16741 VSS.n16740 4.5005
R10121 VSS.n16315 VSS.n16314 4.5005
R10122 VSS.n16324 VSS.n16315 4.5005
R10123 VSS.n16835 VSS.n16834 4.5005
R10124 VSS.n16808 VSS.n16295 4.5005
R10125 VSS.n16808 VSS.n16289 4.5005
R10126 VSS.n16815 VSS.n16291 4.5005
R10127 VSS.n16786 VSS.n16782 4.5005
R10128 VSS.n16786 VSS.n16785 4.5005
R10129 VSS.n16789 VSS.n16780 4.5005
R10130 VSS.n16773 VSS.n16772 4.5005
R10131 VSS.n16772 VSS.n16301 4.5005
R10132 VSS.n16839 VSS.n16838 4.5005
R10133 VSS.n16280 VSS.n16278 4.5005
R10134 VSS.n16278 VSS.n16277 4.5005
R10135 VSS.n16796 VSS.n16795 4.5005
R10136 VSS.n16797 VSS.n16796 4.5005
R10137 VSS.n16292 VSS.n16290 4.5005
R10138 VSS.n16854 VSS.n16853 4.5005
R10139 VSS.n16725 VSS.n16724 4.5005
R10140 VSS.n16726 VSS.n16335 4.5005
R10141 VSS.n16429 VSS.n16424 4.5005
R10142 VSS.n16579 VSS.n16578 4.5005
R10143 VSS.n16555 VSS.n16439 4.5005
R10144 VSS.n16516 VSS.n16515 4.5005
R10145 VSS.n16494 VSS.n16492 4.5005
R10146 VSS.n16493 VSS.n16472 4.5005
R10147 VSS.n16496 VSS.n16495 4.5005
R10148 VSS.n16554 VSS.n16553 4.5005
R10149 VSS.n16441 VSS.n16428 4.5005
R10150 VSS.n16544 VSS.n16543 4.5005
R10151 VSS.n16450 VSS.n16448 4.5005
R10152 VSS.n16464 VSS.n16463 4.5005
R10153 VSS.n16474 VSS.n16466 4.5005
R10154 VSS.n16545 VSS.n16443 4.5005
R10155 VSS.n16577 VSS.n16423 4.5005
R10156 VSS.n16490 VSS.n16489 4.5005
R10157 VSS.n16431 VSS.n16430 4.5005
R10158 VSS.n16566 VSS.n16431 4.5005
R10159 VSS.n16536 VSS.n16449 4.5005
R10160 VSS.n16462 VSS.n16460 4.5005
R10161 VSS.n16460 VSS.n16459 4.5005
R10162 VSS.n16505 VSS.n16473 4.5005
R10163 VSS.n16557 VSS.n16556 4.5005
R10164 VSS.n16557 VSS.n16437 4.5005
R10165 VSS.n16591 VSS.n16590 4.5005
R10166 VSS.n16590 VSS.n16589 4.5005
R10167 VSS.n1526 VSS.n1521 4.5005
R10168 VSS.n16090 VSS.n16089 4.5005
R10169 VSS.n16067 VSS.n1536 4.5005
R10170 VSS.n1564 VSS.n1562 4.5005
R10171 VSS.n16006 VSS.n16004 4.5005
R10172 VSS.n16005 VSS.n1569 4.5005
R10173 VSS.n16008 VSS.n16007 4.5005
R10174 VSS.n16066 VSS.n16065 4.5005
R10175 VSS.n1538 VSS.n1525 4.5005
R10176 VSS.n16056 VSS.n16055 4.5005
R10177 VSS.n1547 VSS.n1545 4.5005
R10178 VSS.n1559 VSS.n1558 4.5005
R10179 VSS.n16028 VSS.n16027 4.5005
R10180 VSS.n1571 VSS.n1561 4.5005
R10181 VSS.n16057 VSS.n1540 4.5005
R10182 VSS.n16088 VSS.n1520 4.5005
R10183 VSS.n16002 VSS.n16001 4.5005
R10184 VSS.n1528 VSS.n1527 4.5005
R10185 VSS.n16077 VSS.n1528 4.5005
R10186 VSS.n1557 VSS.n1555 4.5005
R10187 VSS.n1555 VSS.n1554 4.5005
R10188 VSS.n16017 VSS.n1570 4.5005
R10189 VSS.n16069 VSS.n16068 4.5005
R10190 VSS.n16069 VSS.n1534 4.5005
R10191 VSS.n16124 VSS.n16123 4.5005
R10192 VSS.n16123 VSS.n16122 4.5005
R10193 VSS.n16247 VSS.n1451 4.5005
R10194 VSS.n16188 VSS.n1478 4.5005
R10195 VSS.n16151 VSS.n16150 4.5005
R10196 VSS.n16101 VSS.n16099 4.5005
R10197 VSS.n16130 VSS.n16129 4.5005
R10198 VSS.n16141 VSS.n16140 4.5005
R10199 VSS.n16142 VSS.n16141 4.5005
R10200 VSS.n16175 VSS.n16174 4.5005
R10201 VSS.n16148 VSS.n16147 4.5005
R10202 VSS.n1487 VSS.n1486 4.5005
R10203 VSS.n1496 VSS.n1487 4.5005
R10204 VSS.n16242 VSS.n16241 4.5005
R10205 VSS.n16215 VSS.n1467 4.5005
R10206 VSS.n16215 VSS.n1461 4.5005
R10207 VSS.n16222 VSS.n1463 4.5005
R10208 VSS.n16193 VSS.n16189 4.5005
R10209 VSS.n16193 VSS.n16192 4.5005
R10210 VSS.n16196 VSS.n16187 4.5005
R10211 VSS.n16180 VSS.n16179 4.5005
R10212 VSS.n16179 VSS.n1473 4.5005
R10213 VSS.n16246 VSS.n16245 4.5005
R10214 VSS.n1452 VSS.n1450 4.5005
R10215 VSS.n1450 VSS.n1449 4.5005
R10216 VSS.n16203 VSS.n16202 4.5005
R10217 VSS.n16204 VSS.n16203 4.5005
R10218 VSS.n1464 VSS.n1462 4.5005
R10219 VSS.n16261 VSS.n16260 4.5005
R10220 VSS.n16132 VSS.n16131 4.5005
R10221 VSS.n16133 VSS.n1507 4.5005
R10222 VSS.n1594 VSS.n1589 4.5005
R10223 VSS.n1744 VSS.n1743 4.5005
R10224 VSS.n1720 VSS.n1604 4.5005
R10225 VSS.n1681 VSS.n1680 4.5005
R10226 VSS.n1659 VSS.n1657 4.5005
R10227 VSS.n1658 VSS.n1637 4.5005
R10228 VSS.n1661 VSS.n1660 4.5005
R10229 VSS.n1719 VSS.n1718 4.5005
R10230 VSS.n1606 VSS.n1593 4.5005
R10231 VSS.n1709 VSS.n1708 4.5005
R10232 VSS.n1615 VSS.n1613 4.5005
R10233 VSS.n1629 VSS.n1628 4.5005
R10234 VSS.n1639 VSS.n1631 4.5005
R10235 VSS.n1710 VSS.n1608 4.5005
R10236 VSS.n1742 VSS.n1588 4.5005
R10237 VSS.n1655 VSS.n1654 4.5005
R10238 VSS.n1596 VSS.n1595 4.5005
R10239 VSS.n1731 VSS.n1596 4.5005
R10240 VSS.n1701 VSS.n1614 4.5005
R10241 VSS.n1627 VSS.n1625 4.5005
R10242 VSS.n1625 VSS.n1624 4.5005
R10243 VSS.n1670 VSS.n1638 4.5005
R10244 VSS.n1722 VSS.n1721 4.5005
R10245 VSS.n1722 VSS.n1602 4.5005
R10246 VSS.n15998 VSS.n15997 4.5005
R10247 VSS.n15997 VSS.n15996 4.5005
R10248 VSS.n2060 VSS.n2059 4.5005
R10249 VSS.n2063 VSS.n2062 4.5005
R10250 VSS.n2046 VSS.n2045 4.5005
R10251 VSS.n2021 VSS.n2020 4.5005
R10252 VSS.n2012 VSS.n2011 4.5005
R10253 VSS.n2013 VSS.n2005 4.5005
R10254 VSS.n2009 VSS.n2006 4.5005
R10255 VSS.n1970 VSS.n1968 4.5005
R10256 VSS.n2316 VSS.n2315 4.5005
R10257 VSS.n2323 VSS.n1960 4.5005
R10258 VSS.n2330 VSS.n2329 4.5005
R10259 VSS.n2331 VSS.n1952 4.5005
R10260 VSS.n2017 VSS.n1949 4.5005
R10261 VSS.n2338 VSS.n2337 4.5005
R10262 VSS.n2322 VSS.n2321 4.5005
R10263 VSS.n2061 VSS.n1985 4.5005
R10264 VSS.n2346 VSS.n2345 4.5005
R10265 VSS.n2058 VSS.n1986 4.5005
R10266 VSS.n2058 VSS.n2057 4.5005
R10267 VSS.n2019 VSS.n2018 4.5005
R10268 VSS.n2018 VSS.n1996 4.5005
R10269 VSS.n2015 VSS.n2014 4.5005
R10270 VSS.n2048 VSS.n2047 4.5005
R10271 VSS.n2048 VSS.n2041 4.5005
R10272 VSS.n2308 VSS.n1978 4.5005
R10273 VSS.n2308 VSS.n2307 4.5005
R10274 VSS.n2211 VSS.n2210 4.5005
R10275 VSS.n2181 VSS.n2130 4.5005
R10276 VSS.n2275 VSS.n2274 4.5005
R10277 VSS.n2088 VSS.n2072 4.5005
R10278 VSS.n2096 VSS.n2095 4.5005
R10279 VSS.n2289 VSS.n2080 4.5005
R10280 VSS.n2080 VSS.n2078 4.5005
R10281 VSS.n2143 VSS.n2142 4.5005
R10282 VSS.n2114 VSS.n2113 4.5005
R10283 VSS.n2273 VSS.n2109 4.5005
R10284 VSS.n2109 VSS.n2107 4.5005
R10285 VSS.n2216 VSS.n2200 4.5005
R10286 VSS.n2247 VSS.n2246 4.5005
R10287 VSS.n2248 VSS.n2247 4.5005
R10288 VSS.n2242 VSS.n2161 4.5005
R10289 VSS.n2183 VSS.n2182 4.5005
R10290 VSS.n2183 VSS.n2178 4.5005
R10291 VSS.n2252 VSS.n2154 4.5005
R10292 VSS.n2148 VSS.n2147 4.5005
R10293 VSS.n2147 VSS.n2125 4.5005
R10294 VSS.n2212 VSS.n2208 4.5005
R10295 VSS.n2234 VSS.n2170 4.5005
R10296 VSS.n2234 VSS.n2233 4.5005
R10297 VSS.n2259 VSS.n2258 4.5005
R10298 VSS.n2260 VSS.n2259 4.5005
R10299 VSS.n2245 VSS.n2159 4.5005
R10300 VSS.n2201 VSS.n2199 4.5005
R10301 VSS.n2081 VSS.n2079 4.5005
R10302 VSS.n2097 VSS.n2085 4.5005
R10303 VSS.n1926 VSS.n1773 4.5005
R10304 VSS.n1925 VSS.n1924 4.5005
R10305 VSS.n1795 VSS.n1794 4.5005
R10306 VSS.n1877 VSS.n1876 4.5005
R10307 VSS.n1850 VSS.n1848 4.5005
R10308 VSS.n1849 VSS.n1826 4.5005
R10309 VSS.n1852 VSS.n1851 4.5005
R10310 VSS.n1784 VSS.n1783 4.5005
R10311 VSS.n1915 VSS.n1914 4.5005
R10312 VSS.n1807 VSS.n1806 4.5005
R10313 VSS.n1886 VSS.n1885 4.5005
R10314 VSS.n1884 VSS.n1883 4.5005
R10315 VSS.n1829 VSS.n1813 4.5005
R10316 VSS.n1788 VSS.n1786 4.5005
R10317 VSS.n1923 VSS.n1775 4.5005
R10318 VSS.n1846 VSS.n1845 4.5005
R10319 VSS.n1928 VSS.n1927 4.5005
R10320 VSS.n1928 VSS.n1771 4.5005
R10321 VSS.n1896 VSS.n1804 4.5005
R10322 VSS.n1875 VSS.n1814 4.5005
R10323 VSS.n1875 VSS.n1874 4.5005
R10324 VSS.n1861 VSS.n1827 4.5005
R10325 VSS.n1793 VSS.n1789 4.5005
R10326 VSS.n1791 VSS.n1789 4.5005
R10327 VSS.n1940 VSS.n1939 4.5005
R10328 VSS.n1939 VSS.n1938 4.5005
R10329 VSS.n2903 VSS.n2898 4.5005
R10330 VSS.n3231 VSS.n3230 4.5005
R10331 VSS.n3208 VSS.n2913 4.5005
R10332 VSS.n2941 VSS.n2939 4.5005
R10333 VSS.n3147 VSS.n3145 4.5005
R10334 VSS.n3146 VSS.n2946 4.5005
R10335 VSS.n3149 VSS.n3148 4.5005
R10336 VSS.n3207 VSS.n3206 4.5005
R10337 VSS.n2915 VSS.n2902 4.5005
R10338 VSS.n3197 VSS.n3196 4.5005
R10339 VSS.n2924 VSS.n2922 4.5005
R10340 VSS.n2936 VSS.n2935 4.5005
R10341 VSS.n3169 VSS.n3168 4.5005
R10342 VSS.n2948 VSS.n2938 4.5005
R10343 VSS.n3198 VSS.n2917 4.5005
R10344 VSS.n3229 VSS.n2897 4.5005
R10345 VSS.n3143 VSS.n3142 4.5005
R10346 VSS.n2905 VSS.n2904 4.5005
R10347 VSS.n3218 VSS.n2905 4.5005
R10348 VSS.n2934 VSS.n2932 4.5005
R10349 VSS.n2932 VSS.n2931 4.5005
R10350 VSS.n3158 VSS.n2947 4.5005
R10351 VSS.n3210 VSS.n3209 4.5005
R10352 VSS.n3210 VSS.n2911 4.5005
R10353 VSS.n3265 VSS.n3264 4.5005
R10354 VSS.n3264 VSS.n3263 4.5005
R10355 VSS.n3388 VSS.n2828 4.5005
R10356 VSS.n3329 VSS.n2855 4.5005
R10357 VSS.n3292 VSS.n3291 4.5005
R10358 VSS.n3242 VSS.n3240 4.5005
R10359 VSS.n3271 VSS.n3270 4.5005
R10360 VSS.n3282 VSS.n3281 4.5005
R10361 VSS.n3283 VSS.n3282 4.5005
R10362 VSS.n3316 VSS.n3315 4.5005
R10363 VSS.n3289 VSS.n3288 4.5005
R10364 VSS.n2864 VSS.n2863 4.5005
R10365 VSS.n2873 VSS.n2864 4.5005
R10366 VSS.n3383 VSS.n3382 4.5005
R10367 VSS.n3356 VSS.n2844 4.5005
R10368 VSS.n3356 VSS.n2838 4.5005
R10369 VSS.n3363 VSS.n2840 4.5005
R10370 VSS.n3334 VSS.n3330 4.5005
R10371 VSS.n3334 VSS.n3333 4.5005
R10372 VSS.n3337 VSS.n3328 4.5005
R10373 VSS.n3321 VSS.n3320 4.5005
R10374 VSS.n3320 VSS.n2850 4.5005
R10375 VSS.n3387 VSS.n3386 4.5005
R10376 VSS.n2829 VSS.n2827 4.5005
R10377 VSS.n2827 VSS.n2826 4.5005
R10378 VSS.n3344 VSS.n3343 4.5005
R10379 VSS.n3345 VSS.n3344 4.5005
R10380 VSS.n2841 VSS.n2839 4.5005
R10381 VSS.n3402 VSS.n3401 4.5005
R10382 VSS.n3273 VSS.n3272 4.5005
R10383 VSS.n3274 VSS.n2884 4.5005
R10384 VSS.n3125 VSS.n2972 4.5005
R10385 VSS.n3124 VSS.n3123 4.5005
R10386 VSS.n2994 VSS.n2993 4.5005
R10387 VSS.n3076 VSS.n3075 4.5005
R10388 VSS.n3049 VSS.n3047 4.5005
R10389 VSS.n3048 VSS.n3025 4.5005
R10390 VSS.n3051 VSS.n3050 4.5005
R10391 VSS.n2983 VSS.n2982 4.5005
R10392 VSS.n3114 VSS.n3113 4.5005
R10393 VSS.n3006 VSS.n3005 4.5005
R10394 VSS.n3085 VSS.n3084 4.5005
R10395 VSS.n3083 VSS.n3082 4.5005
R10396 VSS.n3028 VSS.n3012 4.5005
R10397 VSS.n2987 VSS.n2985 4.5005
R10398 VSS.n3122 VSS.n2974 4.5005
R10399 VSS.n3045 VSS.n3044 4.5005
R10400 VSS.n3127 VSS.n3126 4.5005
R10401 VSS.n3127 VSS.n2970 4.5005
R10402 VSS.n3095 VSS.n3003 4.5005
R10403 VSS.n3074 VSS.n3013 4.5005
R10404 VSS.n3074 VSS.n3073 4.5005
R10405 VSS.n3060 VSS.n3026 4.5005
R10406 VSS.n2992 VSS.n2988 4.5005
R10407 VSS.n2990 VSS.n2988 4.5005
R10408 VSS.n3139 VSS.n3138 4.5005
R10409 VSS.n3138 VSS.n3137 4.5005
R10410 VSS.n3495 VSS.n3490 4.5005
R10411 VSS.n3823 VSS.n3822 4.5005
R10412 VSS.n3800 VSS.n3505 4.5005
R10413 VSS.n3533 VSS.n3531 4.5005
R10414 VSS.n3739 VSS.n3737 4.5005
R10415 VSS.n3738 VSS.n3538 4.5005
R10416 VSS.n3741 VSS.n3740 4.5005
R10417 VSS.n3799 VSS.n3798 4.5005
R10418 VSS.n3507 VSS.n3494 4.5005
R10419 VSS.n3789 VSS.n3788 4.5005
R10420 VSS.n3516 VSS.n3514 4.5005
R10421 VSS.n3528 VSS.n3527 4.5005
R10422 VSS.n3761 VSS.n3760 4.5005
R10423 VSS.n3540 VSS.n3530 4.5005
R10424 VSS.n3790 VSS.n3509 4.5005
R10425 VSS.n3821 VSS.n3489 4.5005
R10426 VSS.n3735 VSS.n3734 4.5005
R10427 VSS.n3497 VSS.n3496 4.5005
R10428 VSS.n3810 VSS.n3497 4.5005
R10429 VSS.n3526 VSS.n3524 4.5005
R10430 VSS.n3524 VSS.n3523 4.5005
R10431 VSS.n3750 VSS.n3539 4.5005
R10432 VSS.n3802 VSS.n3801 4.5005
R10433 VSS.n3802 VSS.n3503 4.5005
R10434 VSS.n3857 VSS.n3856 4.5005
R10435 VSS.n3856 VSS.n3855 4.5005
R10436 VSS.n3980 VSS.n3420 4.5005
R10437 VSS.n3921 VSS.n3447 4.5005
R10438 VSS.n3884 VSS.n3883 4.5005
R10439 VSS.n3834 VSS.n3832 4.5005
R10440 VSS.n3863 VSS.n3862 4.5005
R10441 VSS.n3874 VSS.n3873 4.5005
R10442 VSS.n3875 VSS.n3874 4.5005
R10443 VSS.n3908 VSS.n3907 4.5005
R10444 VSS.n3881 VSS.n3880 4.5005
R10445 VSS.n3456 VSS.n3455 4.5005
R10446 VSS.n3465 VSS.n3456 4.5005
R10447 VSS.n3975 VSS.n3974 4.5005
R10448 VSS.n3948 VSS.n3436 4.5005
R10449 VSS.n3948 VSS.n3430 4.5005
R10450 VSS.n3955 VSS.n3432 4.5005
R10451 VSS.n3926 VSS.n3922 4.5005
R10452 VSS.n3926 VSS.n3925 4.5005
R10453 VSS.n3929 VSS.n3920 4.5005
R10454 VSS.n3913 VSS.n3912 4.5005
R10455 VSS.n3912 VSS.n3442 4.5005
R10456 VSS.n3979 VSS.n3978 4.5005
R10457 VSS.n3421 VSS.n3419 4.5005
R10458 VSS.n3419 VSS.n3418 4.5005
R10459 VSS.n3936 VSS.n3935 4.5005
R10460 VSS.n3937 VSS.n3936 4.5005
R10461 VSS.n3433 VSS.n3431 4.5005
R10462 VSS.n3994 VSS.n3993 4.5005
R10463 VSS.n3865 VSS.n3864 4.5005
R10464 VSS.n3866 VSS.n3476 4.5005
R10465 VSS.n3717 VSS.n3564 4.5005
R10466 VSS.n3716 VSS.n3715 4.5005
R10467 VSS.n3586 VSS.n3585 4.5005
R10468 VSS.n3668 VSS.n3667 4.5005
R10469 VSS.n3641 VSS.n3639 4.5005
R10470 VSS.n3640 VSS.n3617 4.5005
R10471 VSS.n3643 VSS.n3642 4.5005
R10472 VSS.n3575 VSS.n3574 4.5005
R10473 VSS.n3706 VSS.n3705 4.5005
R10474 VSS.n3598 VSS.n3597 4.5005
R10475 VSS.n3677 VSS.n3676 4.5005
R10476 VSS.n3675 VSS.n3674 4.5005
R10477 VSS.n3620 VSS.n3604 4.5005
R10478 VSS.n3579 VSS.n3577 4.5005
R10479 VSS.n3714 VSS.n3566 4.5005
R10480 VSS.n3637 VSS.n3636 4.5005
R10481 VSS.n3719 VSS.n3718 4.5005
R10482 VSS.n3719 VSS.n3562 4.5005
R10483 VSS.n3687 VSS.n3595 4.5005
R10484 VSS.n3666 VSS.n3605 4.5005
R10485 VSS.n3666 VSS.n3665 4.5005
R10486 VSS.n3652 VSS.n3618 4.5005
R10487 VSS.n3584 VSS.n3580 4.5005
R10488 VSS.n3582 VSS.n3580 4.5005
R10489 VSS.n3731 VSS.n3730 4.5005
R10490 VSS.n3730 VSS.n3729 4.5005
R10491 VSS.n4087 VSS.n4082 4.5005
R10492 VSS.n4415 VSS.n4414 4.5005
R10493 VSS.n4392 VSS.n4097 4.5005
R10494 VSS.n4125 VSS.n4123 4.5005
R10495 VSS.n4331 VSS.n4329 4.5005
R10496 VSS.n4330 VSS.n4130 4.5005
R10497 VSS.n4333 VSS.n4332 4.5005
R10498 VSS.n4391 VSS.n4390 4.5005
R10499 VSS.n4099 VSS.n4086 4.5005
R10500 VSS.n4381 VSS.n4380 4.5005
R10501 VSS.n4108 VSS.n4106 4.5005
R10502 VSS.n4120 VSS.n4119 4.5005
R10503 VSS.n4353 VSS.n4352 4.5005
R10504 VSS.n4132 VSS.n4122 4.5005
R10505 VSS.n4382 VSS.n4101 4.5005
R10506 VSS.n4413 VSS.n4081 4.5005
R10507 VSS.n4327 VSS.n4326 4.5005
R10508 VSS.n4089 VSS.n4088 4.5005
R10509 VSS.n4402 VSS.n4089 4.5005
R10510 VSS.n4118 VSS.n4116 4.5005
R10511 VSS.n4116 VSS.n4115 4.5005
R10512 VSS.n4342 VSS.n4131 4.5005
R10513 VSS.n4394 VSS.n4393 4.5005
R10514 VSS.n4394 VSS.n4095 4.5005
R10515 VSS.n4449 VSS.n4448 4.5005
R10516 VSS.n4448 VSS.n4447 4.5005
R10517 VSS.n4572 VSS.n4012 4.5005
R10518 VSS.n4513 VSS.n4039 4.5005
R10519 VSS.n4476 VSS.n4475 4.5005
R10520 VSS.n4426 VSS.n4424 4.5005
R10521 VSS.n4455 VSS.n4454 4.5005
R10522 VSS.n4466 VSS.n4465 4.5005
R10523 VSS.n4467 VSS.n4466 4.5005
R10524 VSS.n4500 VSS.n4499 4.5005
R10525 VSS.n4473 VSS.n4472 4.5005
R10526 VSS.n4048 VSS.n4047 4.5005
R10527 VSS.n4057 VSS.n4048 4.5005
R10528 VSS.n4567 VSS.n4566 4.5005
R10529 VSS.n4540 VSS.n4028 4.5005
R10530 VSS.n4540 VSS.n4022 4.5005
R10531 VSS.n4547 VSS.n4024 4.5005
R10532 VSS.n4518 VSS.n4514 4.5005
R10533 VSS.n4518 VSS.n4517 4.5005
R10534 VSS.n4521 VSS.n4512 4.5005
R10535 VSS.n4505 VSS.n4504 4.5005
R10536 VSS.n4504 VSS.n4034 4.5005
R10537 VSS.n4571 VSS.n4570 4.5005
R10538 VSS.n4013 VSS.n4011 4.5005
R10539 VSS.n4011 VSS.n4010 4.5005
R10540 VSS.n4528 VSS.n4527 4.5005
R10541 VSS.n4529 VSS.n4528 4.5005
R10542 VSS.n4025 VSS.n4023 4.5005
R10543 VSS.n4586 VSS.n4585 4.5005
R10544 VSS.n4457 VSS.n4456 4.5005
R10545 VSS.n4458 VSS.n4068 4.5005
R10546 VSS.n4309 VSS.n4156 4.5005
R10547 VSS.n4308 VSS.n4307 4.5005
R10548 VSS.n4178 VSS.n4177 4.5005
R10549 VSS.n4260 VSS.n4259 4.5005
R10550 VSS.n4233 VSS.n4231 4.5005
R10551 VSS.n4232 VSS.n4209 4.5005
R10552 VSS.n4235 VSS.n4234 4.5005
R10553 VSS.n4167 VSS.n4166 4.5005
R10554 VSS.n4298 VSS.n4297 4.5005
R10555 VSS.n4190 VSS.n4189 4.5005
R10556 VSS.n4269 VSS.n4268 4.5005
R10557 VSS.n4267 VSS.n4266 4.5005
R10558 VSS.n4212 VSS.n4196 4.5005
R10559 VSS.n4171 VSS.n4169 4.5005
R10560 VSS.n4306 VSS.n4158 4.5005
R10561 VSS.n4229 VSS.n4228 4.5005
R10562 VSS.n4311 VSS.n4310 4.5005
R10563 VSS.n4311 VSS.n4154 4.5005
R10564 VSS.n4279 VSS.n4187 4.5005
R10565 VSS.n4258 VSS.n4197 4.5005
R10566 VSS.n4258 VSS.n4257 4.5005
R10567 VSS.n4244 VSS.n4210 4.5005
R10568 VSS.n4176 VSS.n4172 4.5005
R10569 VSS.n4174 VSS.n4172 4.5005
R10570 VSS.n4323 VSS.n4322 4.5005
R10571 VSS.n4322 VSS.n4321 4.5005
R10572 VSS.n4679 VSS.n4674 4.5005
R10573 VSS.n5007 VSS.n5006 4.5005
R10574 VSS.n4984 VSS.n4689 4.5005
R10575 VSS.n4717 VSS.n4715 4.5005
R10576 VSS.n4923 VSS.n4921 4.5005
R10577 VSS.n4922 VSS.n4722 4.5005
R10578 VSS.n4925 VSS.n4924 4.5005
R10579 VSS.n4983 VSS.n4982 4.5005
R10580 VSS.n4691 VSS.n4678 4.5005
R10581 VSS.n4973 VSS.n4972 4.5005
R10582 VSS.n4700 VSS.n4698 4.5005
R10583 VSS.n4712 VSS.n4711 4.5005
R10584 VSS.n4945 VSS.n4944 4.5005
R10585 VSS.n4724 VSS.n4714 4.5005
R10586 VSS.n4974 VSS.n4693 4.5005
R10587 VSS.n5005 VSS.n4673 4.5005
R10588 VSS.n4919 VSS.n4918 4.5005
R10589 VSS.n4681 VSS.n4680 4.5005
R10590 VSS.n4994 VSS.n4681 4.5005
R10591 VSS.n4710 VSS.n4708 4.5005
R10592 VSS.n4708 VSS.n4707 4.5005
R10593 VSS.n4934 VSS.n4723 4.5005
R10594 VSS.n4986 VSS.n4985 4.5005
R10595 VSS.n4986 VSS.n4687 4.5005
R10596 VSS.n5041 VSS.n5040 4.5005
R10597 VSS.n5040 VSS.n5039 4.5005
R10598 VSS.n5164 VSS.n4604 4.5005
R10599 VSS.n5105 VSS.n4631 4.5005
R10600 VSS.n5068 VSS.n5067 4.5005
R10601 VSS.n5018 VSS.n5016 4.5005
R10602 VSS.n5047 VSS.n5046 4.5005
R10603 VSS.n5058 VSS.n5057 4.5005
R10604 VSS.n5059 VSS.n5058 4.5005
R10605 VSS.n5092 VSS.n5091 4.5005
R10606 VSS.n5065 VSS.n5064 4.5005
R10607 VSS.n4640 VSS.n4639 4.5005
R10608 VSS.n4649 VSS.n4640 4.5005
R10609 VSS.n5159 VSS.n5158 4.5005
R10610 VSS.n5132 VSS.n4620 4.5005
R10611 VSS.n5132 VSS.n4614 4.5005
R10612 VSS.n5139 VSS.n4616 4.5005
R10613 VSS.n5110 VSS.n5106 4.5005
R10614 VSS.n5110 VSS.n5109 4.5005
R10615 VSS.n5113 VSS.n5104 4.5005
R10616 VSS.n5097 VSS.n5096 4.5005
R10617 VSS.n5096 VSS.n4626 4.5005
R10618 VSS.n5163 VSS.n5162 4.5005
R10619 VSS.n4605 VSS.n4603 4.5005
R10620 VSS.n4603 VSS.n4602 4.5005
R10621 VSS.n5120 VSS.n5119 4.5005
R10622 VSS.n5121 VSS.n5120 4.5005
R10623 VSS.n4617 VSS.n4615 4.5005
R10624 VSS.n5178 VSS.n5177 4.5005
R10625 VSS.n5049 VSS.n5048 4.5005
R10626 VSS.n5050 VSS.n4660 4.5005
R10627 VSS.n4901 VSS.n4748 4.5005
R10628 VSS.n4900 VSS.n4899 4.5005
R10629 VSS.n4770 VSS.n4769 4.5005
R10630 VSS.n4852 VSS.n4851 4.5005
R10631 VSS.n4825 VSS.n4823 4.5005
R10632 VSS.n4824 VSS.n4801 4.5005
R10633 VSS.n4827 VSS.n4826 4.5005
R10634 VSS.n4759 VSS.n4758 4.5005
R10635 VSS.n4890 VSS.n4889 4.5005
R10636 VSS.n4782 VSS.n4781 4.5005
R10637 VSS.n4861 VSS.n4860 4.5005
R10638 VSS.n4859 VSS.n4858 4.5005
R10639 VSS.n4804 VSS.n4788 4.5005
R10640 VSS.n4763 VSS.n4761 4.5005
R10641 VSS.n4898 VSS.n4750 4.5005
R10642 VSS.n4821 VSS.n4820 4.5005
R10643 VSS.n4903 VSS.n4902 4.5005
R10644 VSS.n4903 VSS.n4746 4.5005
R10645 VSS.n4871 VSS.n4779 4.5005
R10646 VSS.n4850 VSS.n4789 4.5005
R10647 VSS.n4850 VSS.n4849 4.5005
R10648 VSS.n4836 VSS.n4802 4.5005
R10649 VSS.n4768 VSS.n4764 4.5005
R10650 VSS.n4766 VSS.n4764 4.5005
R10651 VSS.n4915 VSS.n4914 4.5005
R10652 VSS.n4914 VSS.n4913 4.5005
R10653 VSS.n2656 VSS.n2655 4.5005
R10654 VSS.n2659 VSS.n2658 4.5005
R10655 VSS.n2642 VSS.n2641 4.5005
R10656 VSS.n2617 VSS.n2616 4.5005
R10657 VSS.n2608 VSS.n2607 4.5005
R10658 VSS.n2609 VSS.n2601 4.5005
R10659 VSS.n2605 VSS.n2602 4.5005
R10660 VSS.n2566 VSS.n2564 4.5005
R10661 VSS.n5281 VSS.n5280 4.5005
R10662 VSS.n5288 VSS.n2556 4.5005
R10663 VSS.n5295 VSS.n5294 4.5005
R10664 VSS.n5296 VSS.n2548 4.5005
R10665 VSS.n2613 VSS.n2545 4.5005
R10666 VSS.n5303 VSS.n5302 4.5005
R10667 VSS.n5287 VSS.n5286 4.5005
R10668 VSS.n2657 VSS.n2581 4.5005
R10669 VSS.n5311 VSS.n5310 4.5005
R10670 VSS.n2654 VSS.n2582 4.5005
R10671 VSS.n2654 VSS.n2653 4.5005
R10672 VSS.n2615 VSS.n2614 4.5005
R10673 VSS.n2614 VSS.n2592 4.5005
R10674 VSS.n2611 VSS.n2610 4.5005
R10675 VSS.n2644 VSS.n2643 4.5005
R10676 VSS.n2644 VSS.n2637 4.5005
R10677 VSS.n5273 VSS.n2574 4.5005
R10678 VSS.n5273 VSS.n5272 4.5005
R10679 VSS.n2807 VSS.n2806 4.5005
R10680 VSS.n2777 VSS.n2726 4.5005
R10681 VSS.n5240 VSS.n5239 4.5005
R10682 VSS.n2684 VSS.n2668 4.5005
R10683 VSS.n2692 VSS.n2691 4.5005
R10684 VSS.n5254 VSS.n2676 4.5005
R10685 VSS.n2676 VSS.n2674 4.5005
R10686 VSS.n2739 VSS.n2738 4.5005
R10687 VSS.n2710 VSS.n2709 4.5005
R10688 VSS.n5238 VSS.n2705 4.5005
R10689 VSS.n2705 VSS.n2703 4.5005
R10690 VSS.n2812 VSS.n2796 4.5005
R10691 VSS.n5212 VSS.n5211 4.5005
R10692 VSS.n5213 VSS.n5212 4.5005
R10693 VSS.n5207 VSS.n2757 4.5005
R10694 VSS.n2779 VSS.n2778 4.5005
R10695 VSS.n2779 VSS.n2774 4.5005
R10696 VSS.n5217 VSS.n2750 4.5005
R10697 VSS.n2744 VSS.n2743 4.5005
R10698 VSS.n2743 VSS.n2721 4.5005
R10699 VSS.n2808 VSS.n2804 4.5005
R10700 VSS.n5199 VSS.n2766 4.5005
R10701 VSS.n5199 VSS.n5198 4.5005
R10702 VSS.n5224 VSS.n5223 4.5005
R10703 VSS.n5225 VSS.n5224 4.5005
R10704 VSS.n5210 VSS.n2755 4.5005
R10705 VSS.n2797 VSS.n2795 4.5005
R10706 VSS.n2677 VSS.n2675 4.5005
R10707 VSS.n2693 VSS.n2681 4.5005
R10708 VSS.n2522 VSS.n2369 4.5005
R10709 VSS.n2521 VSS.n2520 4.5005
R10710 VSS.n2391 VSS.n2390 4.5005
R10711 VSS.n2473 VSS.n2472 4.5005
R10712 VSS.n2446 VSS.n2444 4.5005
R10713 VSS.n2445 VSS.n2422 4.5005
R10714 VSS.n2448 VSS.n2447 4.5005
R10715 VSS.n2380 VSS.n2379 4.5005
R10716 VSS.n2511 VSS.n2510 4.5005
R10717 VSS.n2403 VSS.n2402 4.5005
R10718 VSS.n2482 VSS.n2481 4.5005
R10719 VSS.n2480 VSS.n2479 4.5005
R10720 VSS.n2425 VSS.n2409 4.5005
R10721 VSS.n2384 VSS.n2382 4.5005
R10722 VSS.n2519 VSS.n2371 4.5005
R10723 VSS.n2442 VSS.n2441 4.5005
R10724 VSS.n2524 VSS.n2523 4.5005
R10725 VSS.n2524 VSS.n2367 4.5005
R10726 VSS.n2492 VSS.n2400 4.5005
R10727 VSS.n2471 VSS.n2410 4.5005
R10728 VSS.n2471 VSS.n2470 4.5005
R10729 VSS.n2457 VSS.n2423 4.5005
R10730 VSS.n2389 VSS.n2385 4.5005
R10731 VSS.n2387 VSS.n2385 4.5005
R10732 VSS.n2536 VSS.n2535 4.5005
R10733 VSS.n2535 VSS.n2534 4.5005
R10734 VSS.n5617 VSS.n5616 4.5005
R10735 VSS.n5620 VSS.n5619 4.5005
R10736 VSS.n5603 VSS.n5602 4.5005
R10737 VSS.n5578 VSS.n5577 4.5005
R10738 VSS.n5569 VSS.n5568 4.5005
R10739 VSS.n5570 VSS.n5562 4.5005
R10740 VSS.n5566 VSS.n5563 4.5005
R10741 VSS.n5527 VSS.n5525 4.5005
R10742 VSS.n5854 VSS.n5853 4.5005
R10743 VSS.n5861 VSS.n5517 4.5005
R10744 VSS.n5868 VSS.n5867 4.5005
R10745 VSS.n5869 VSS.n5509 4.5005
R10746 VSS.n5574 VSS.n5506 4.5005
R10747 VSS.n5876 VSS.n5875 4.5005
R10748 VSS.n5860 VSS.n5859 4.5005
R10749 VSS.n5618 VSS.n5542 4.5005
R10750 VSS.n5884 VSS.n5883 4.5005
R10751 VSS.n5615 VSS.n5543 4.5005
R10752 VSS.n5615 VSS.n5614 4.5005
R10753 VSS.n5576 VSS.n5575 4.5005
R10754 VSS.n5575 VSS.n5553 4.5005
R10755 VSS.n5572 VSS.n5571 4.5005
R10756 VSS.n5605 VSS.n5604 4.5005
R10757 VSS.n5605 VSS.n5598 4.5005
R10758 VSS.n5846 VSS.n5535 4.5005
R10759 VSS.n5846 VSS.n5845 4.5005
R10760 VSS.n5739 VSS.n5729 4.5005
R10761 VSS.n5751 VSS.n5687 4.5005
R10762 VSS.n5813 VSS.n5812 4.5005
R10763 VSS.n5645 VSS.n5629 4.5005
R10764 VSS.n5653 VSS.n5652 4.5005
R10765 VSS.n5827 VSS.n5637 4.5005
R10766 VSS.n5637 VSS.n5635 4.5005
R10767 VSS.n5700 VSS.n5699 4.5005
R10768 VSS.n5671 VSS.n5670 4.5005
R10769 VSS.n5811 VSS.n5666 4.5005
R10770 VSS.n5666 VSS.n5664 4.5005
R10771 VSS.n5734 VSS.n5733 4.5005
R10772 VSS.n5785 VSS.n5784 4.5005
R10773 VSS.n5786 VSS.n5785 4.5005
R10774 VSS.n5780 VSS.n5718 4.5005
R10775 VSS.n5753 VSS.n5752 4.5005
R10776 VSS.n5753 VSS.n5748 4.5005
R10777 VSS.n5790 VSS.n5711 4.5005
R10778 VSS.n5705 VSS.n5704 4.5005
R10779 VSS.n5704 VSS.n5682 4.5005
R10780 VSS.n5738 VSS.n5737 4.5005
R10781 VSS.n5772 VSS.n5727 4.5005
R10782 VSS.n5772 VSS.n5771 4.5005
R10783 VSS.n5797 VSS.n5796 4.5005
R10784 VSS.n5798 VSS.n5797 4.5005
R10785 VSS.n5783 VSS.n5716 4.5005
R10786 VSS.n18884 VSS.n18883 4.5005
R10787 VSS.n5638 VSS.n5636 4.5005
R10788 VSS.n5654 VSS.n5642 4.5005
R10789 VSS.n5483 VSS.n5330 4.5005
R10790 VSS.n5482 VSS.n5481 4.5005
R10791 VSS.n5352 VSS.n5351 4.5005
R10792 VSS.n5434 VSS.n5433 4.5005
R10793 VSS.n5407 VSS.n5405 4.5005
R10794 VSS.n5406 VSS.n5383 4.5005
R10795 VSS.n5409 VSS.n5408 4.5005
R10796 VSS.n5341 VSS.n5340 4.5005
R10797 VSS.n5472 VSS.n5471 4.5005
R10798 VSS.n5364 VSS.n5363 4.5005
R10799 VSS.n5443 VSS.n5442 4.5005
R10800 VSS.n5441 VSS.n5440 4.5005
R10801 VSS.n5386 VSS.n5370 4.5005
R10802 VSS.n5345 VSS.n5343 4.5005
R10803 VSS.n5480 VSS.n5332 4.5005
R10804 VSS.n5403 VSS.n5402 4.5005
R10805 VSS.n5485 VSS.n5484 4.5005
R10806 VSS.n5485 VSS.n5328 4.5005
R10807 VSS.n5453 VSS.n5361 4.5005
R10808 VSS.n5432 VSS.n5371 4.5005
R10809 VSS.n5432 VSS.n5431 4.5005
R10810 VSS.n5418 VSS.n5384 4.5005
R10811 VSS.n5350 VSS.n5346 4.5005
R10812 VSS.n5348 VSS.n5346 4.5005
R10813 VSS.n5497 VSS.n5496 4.5005
R10814 VSS.n5496 VSS.n5495 4.5005
R10815 VSS.n6190 VSS.n6189 4.5005
R10816 VSS.n6193 VSS.n6192 4.5005
R10817 VSS.n6176 VSS.n6175 4.5005
R10818 VSS.n6151 VSS.n6150 4.5005
R10819 VSS.n6142 VSS.n6141 4.5005
R10820 VSS.n6143 VSS.n6135 4.5005
R10821 VSS.n6139 VSS.n6136 4.5005
R10822 VSS.n6100 VSS.n6098 4.5005
R10823 VSS.n6446 VSS.n6445 4.5005
R10824 VSS.n6453 VSS.n6090 4.5005
R10825 VSS.n6460 VSS.n6459 4.5005
R10826 VSS.n6461 VSS.n6082 4.5005
R10827 VSS.n6147 VSS.n6079 4.5005
R10828 VSS.n6468 VSS.n6467 4.5005
R10829 VSS.n6452 VSS.n6451 4.5005
R10830 VSS.n6191 VSS.n6115 4.5005
R10831 VSS.n6476 VSS.n6475 4.5005
R10832 VSS.n6188 VSS.n6116 4.5005
R10833 VSS.n6188 VSS.n6187 4.5005
R10834 VSS.n6149 VSS.n6148 4.5005
R10835 VSS.n6148 VSS.n6126 4.5005
R10836 VSS.n6145 VSS.n6144 4.5005
R10837 VSS.n6178 VSS.n6177 4.5005
R10838 VSS.n6178 VSS.n6171 4.5005
R10839 VSS.n6438 VSS.n6108 4.5005
R10840 VSS.n6438 VSS.n6437 4.5005
R10841 VSS.n6341 VSS.n6340 4.5005
R10842 VSS.n6311 VSS.n6260 4.5005
R10843 VSS.n6405 VSS.n6404 4.5005
R10844 VSS.n6218 VSS.n6202 4.5005
R10845 VSS.n6226 VSS.n6225 4.5005
R10846 VSS.n6419 VSS.n6210 4.5005
R10847 VSS.n6210 VSS.n6208 4.5005
R10848 VSS.n6273 VSS.n6272 4.5005
R10849 VSS.n6244 VSS.n6243 4.5005
R10850 VSS.n6403 VSS.n6239 4.5005
R10851 VSS.n6239 VSS.n6237 4.5005
R10852 VSS.n6346 VSS.n6330 4.5005
R10853 VSS.n6377 VSS.n6376 4.5005
R10854 VSS.n6378 VSS.n6377 4.5005
R10855 VSS.n6372 VSS.n6291 4.5005
R10856 VSS.n6313 VSS.n6312 4.5005
R10857 VSS.n6313 VSS.n6308 4.5005
R10858 VSS.n6382 VSS.n6284 4.5005
R10859 VSS.n6278 VSS.n6277 4.5005
R10860 VSS.n6277 VSS.n6255 4.5005
R10861 VSS.n6342 VSS.n6338 4.5005
R10862 VSS.n6364 VSS.n6300 4.5005
R10863 VSS.n6364 VSS.n6363 4.5005
R10864 VSS.n6389 VSS.n6388 4.5005
R10865 VSS.n6390 VSS.n6389 4.5005
R10866 VSS.n6375 VSS.n6289 4.5005
R10867 VSS.n6331 VSS.n6329 4.5005
R10868 VSS.n6211 VSS.n6209 4.5005
R10869 VSS.n6227 VSS.n6215 4.5005
R10870 VSS.n6056 VSS.n5903 4.5005
R10871 VSS.n6055 VSS.n6054 4.5005
R10872 VSS.n5925 VSS.n5924 4.5005
R10873 VSS.n6007 VSS.n6006 4.5005
R10874 VSS.n5980 VSS.n5978 4.5005
R10875 VSS.n5979 VSS.n5956 4.5005
R10876 VSS.n5982 VSS.n5981 4.5005
R10877 VSS.n5914 VSS.n5913 4.5005
R10878 VSS.n6045 VSS.n6044 4.5005
R10879 VSS.n5937 VSS.n5936 4.5005
R10880 VSS.n6016 VSS.n6015 4.5005
R10881 VSS.n6014 VSS.n6013 4.5005
R10882 VSS.n5959 VSS.n5943 4.5005
R10883 VSS.n5918 VSS.n5916 4.5005
R10884 VSS.n6053 VSS.n5905 4.5005
R10885 VSS.n5976 VSS.n5975 4.5005
R10886 VSS.n6058 VSS.n6057 4.5005
R10887 VSS.n6058 VSS.n5901 4.5005
R10888 VSS.n6026 VSS.n5934 4.5005
R10889 VSS.n6005 VSS.n5944 4.5005
R10890 VSS.n6005 VSS.n6004 4.5005
R10891 VSS.n5991 VSS.n5957 4.5005
R10892 VSS.n5923 VSS.n5919 4.5005
R10893 VSS.n5921 VSS.n5919 4.5005
R10894 VSS.n6070 VSS.n6069 4.5005
R10895 VSS.n6069 VSS.n6068 4.5005
R10896 VSS.n7636 VSS.n7631 4.5005
R10897 VSS.n7964 VSS.n7963 4.5005
R10898 VSS.n7941 VSS.n7646 4.5005
R10899 VSS.n7674 VSS.n7672 4.5005
R10900 VSS.n7880 VSS.n7878 4.5005
R10901 VSS.n7879 VSS.n7679 4.5005
R10902 VSS.n7882 VSS.n7881 4.5005
R10903 VSS.n7940 VSS.n7939 4.5005
R10904 VSS.n7648 VSS.n7635 4.5005
R10905 VSS.n7930 VSS.n7929 4.5005
R10906 VSS.n7657 VSS.n7655 4.5005
R10907 VSS.n7669 VSS.n7668 4.5005
R10908 VSS.n7902 VSS.n7901 4.5005
R10909 VSS.n7681 VSS.n7671 4.5005
R10910 VSS.n7931 VSS.n7650 4.5005
R10911 VSS.n7962 VSS.n7630 4.5005
R10912 VSS.n7876 VSS.n7875 4.5005
R10913 VSS.n7638 VSS.n7637 4.5005
R10914 VSS.n7951 VSS.n7638 4.5005
R10915 VSS.n7667 VSS.n7665 4.5005
R10916 VSS.n7665 VSS.n7664 4.5005
R10917 VSS.n7891 VSS.n7680 4.5005
R10918 VSS.n7943 VSS.n7942 4.5005
R10919 VSS.n7943 VSS.n7644 4.5005
R10920 VSS.n7998 VSS.n7997 4.5005
R10921 VSS.n7997 VSS.n7996 4.5005
R10922 VSS.n8121 VSS.n7561 4.5005
R10923 VSS.n8062 VSS.n7588 4.5005
R10924 VSS.n8025 VSS.n8024 4.5005
R10925 VSS.n7975 VSS.n7973 4.5005
R10926 VSS.n8004 VSS.n8003 4.5005
R10927 VSS.n8015 VSS.n8014 4.5005
R10928 VSS.n8016 VSS.n8015 4.5005
R10929 VSS.n8049 VSS.n8048 4.5005
R10930 VSS.n8022 VSS.n8021 4.5005
R10931 VSS.n7597 VSS.n7596 4.5005
R10932 VSS.n7606 VSS.n7597 4.5005
R10933 VSS.n8116 VSS.n8115 4.5005
R10934 VSS.n8089 VSS.n7577 4.5005
R10935 VSS.n8089 VSS.n7571 4.5005
R10936 VSS.n8096 VSS.n7573 4.5005
R10937 VSS.n8067 VSS.n8063 4.5005
R10938 VSS.n8067 VSS.n8066 4.5005
R10939 VSS.n8070 VSS.n8061 4.5005
R10940 VSS.n8054 VSS.n8053 4.5005
R10941 VSS.n8053 VSS.n7583 4.5005
R10942 VSS.n8120 VSS.n8119 4.5005
R10943 VSS.n7562 VSS.n7560 4.5005
R10944 VSS.n7560 VSS.n7559 4.5005
R10945 VSS.n8077 VSS.n8076 4.5005
R10946 VSS.n8078 VSS.n8077 4.5005
R10947 VSS.n7574 VSS.n7572 4.5005
R10948 VSS.n8135 VSS.n8134 4.5005
R10949 VSS.n8006 VSS.n8005 4.5005
R10950 VSS.n8007 VSS.n7617 4.5005
R10951 VSS.n7858 VSS.n7705 4.5005
R10952 VSS.n7857 VSS.n7856 4.5005
R10953 VSS.n7727 VSS.n7726 4.5005
R10954 VSS.n7809 VSS.n7808 4.5005
R10955 VSS.n7782 VSS.n7780 4.5005
R10956 VSS.n7781 VSS.n7758 4.5005
R10957 VSS.n7784 VSS.n7783 4.5005
R10958 VSS.n7716 VSS.n7715 4.5005
R10959 VSS.n7847 VSS.n7846 4.5005
R10960 VSS.n7739 VSS.n7738 4.5005
R10961 VSS.n7818 VSS.n7817 4.5005
R10962 VSS.n7816 VSS.n7815 4.5005
R10963 VSS.n7761 VSS.n7745 4.5005
R10964 VSS.n7720 VSS.n7718 4.5005
R10965 VSS.n7855 VSS.n7707 4.5005
R10966 VSS.n7778 VSS.n7777 4.5005
R10967 VSS.n7860 VSS.n7859 4.5005
R10968 VSS.n7860 VSS.n7703 4.5005
R10969 VSS.n7828 VSS.n7736 4.5005
R10970 VSS.n7807 VSS.n7746 4.5005
R10971 VSS.n7807 VSS.n7806 4.5005
R10972 VSS.n7793 VSS.n7759 4.5005
R10973 VSS.n7725 VSS.n7721 4.5005
R10974 VSS.n7723 VSS.n7721 4.5005
R10975 VSS.n7872 VSS.n7871 4.5005
R10976 VSS.n7871 VSS.n7870 4.5005
R10977 VSS.n8228 VSS.n8223 4.5005
R10978 VSS.n8556 VSS.n8555 4.5005
R10979 VSS.n8533 VSS.n8238 4.5005
R10980 VSS.n8266 VSS.n8264 4.5005
R10981 VSS.n8472 VSS.n8470 4.5005
R10982 VSS.n8471 VSS.n8271 4.5005
R10983 VSS.n8474 VSS.n8473 4.5005
R10984 VSS.n8532 VSS.n8531 4.5005
R10985 VSS.n8240 VSS.n8227 4.5005
R10986 VSS.n8522 VSS.n8521 4.5005
R10987 VSS.n8249 VSS.n8247 4.5005
R10988 VSS.n8261 VSS.n8260 4.5005
R10989 VSS.n8494 VSS.n8493 4.5005
R10990 VSS.n8273 VSS.n8263 4.5005
R10991 VSS.n8523 VSS.n8242 4.5005
R10992 VSS.n8554 VSS.n8222 4.5005
R10993 VSS.n8468 VSS.n8467 4.5005
R10994 VSS.n8230 VSS.n8229 4.5005
R10995 VSS.n8543 VSS.n8230 4.5005
R10996 VSS.n8259 VSS.n8257 4.5005
R10997 VSS.n8257 VSS.n8256 4.5005
R10998 VSS.n8483 VSS.n8272 4.5005
R10999 VSS.n8535 VSS.n8534 4.5005
R11000 VSS.n8535 VSS.n8236 4.5005
R11001 VSS.n8590 VSS.n8589 4.5005
R11002 VSS.n8589 VSS.n8588 4.5005
R11003 VSS.n8713 VSS.n8153 4.5005
R11004 VSS.n8654 VSS.n8180 4.5005
R11005 VSS.n8617 VSS.n8616 4.5005
R11006 VSS.n8567 VSS.n8565 4.5005
R11007 VSS.n8596 VSS.n8595 4.5005
R11008 VSS.n8607 VSS.n8606 4.5005
R11009 VSS.n8608 VSS.n8607 4.5005
R11010 VSS.n8641 VSS.n8640 4.5005
R11011 VSS.n8614 VSS.n8613 4.5005
R11012 VSS.n8189 VSS.n8188 4.5005
R11013 VSS.n8198 VSS.n8189 4.5005
R11014 VSS.n8708 VSS.n8707 4.5005
R11015 VSS.n8681 VSS.n8169 4.5005
R11016 VSS.n8681 VSS.n8163 4.5005
R11017 VSS.n8688 VSS.n8165 4.5005
R11018 VSS.n8659 VSS.n8655 4.5005
R11019 VSS.n8659 VSS.n8658 4.5005
R11020 VSS.n8662 VSS.n8653 4.5005
R11021 VSS.n8646 VSS.n8645 4.5005
R11022 VSS.n8645 VSS.n8175 4.5005
R11023 VSS.n8712 VSS.n8711 4.5005
R11024 VSS.n8154 VSS.n8152 4.5005
R11025 VSS.n8152 VSS.n8151 4.5005
R11026 VSS.n8669 VSS.n8668 4.5005
R11027 VSS.n8670 VSS.n8669 4.5005
R11028 VSS.n8166 VSS.n8164 4.5005
R11029 VSS.n8727 VSS.n8726 4.5005
R11030 VSS.n8598 VSS.n8597 4.5005
R11031 VSS.n8599 VSS.n8209 4.5005
R11032 VSS.n8450 VSS.n8297 4.5005
R11033 VSS.n8449 VSS.n8448 4.5005
R11034 VSS.n8319 VSS.n8318 4.5005
R11035 VSS.n8401 VSS.n8400 4.5005
R11036 VSS.n8374 VSS.n8372 4.5005
R11037 VSS.n8373 VSS.n8350 4.5005
R11038 VSS.n8376 VSS.n8375 4.5005
R11039 VSS.n8308 VSS.n8307 4.5005
R11040 VSS.n8439 VSS.n8438 4.5005
R11041 VSS.n8331 VSS.n8330 4.5005
R11042 VSS.n8410 VSS.n8409 4.5005
R11043 VSS.n8408 VSS.n8407 4.5005
R11044 VSS.n8353 VSS.n8337 4.5005
R11045 VSS.n8312 VSS.n8310 4.5005
R11046 VSS.n8447 VSS.n8299 4.5005
R11047 VSS.n8370 VSS.n8369 4.5005
R11048 VSS.n8452 VSS.n8451 4.5005
R11049 VSS.n8452 VSS.n8295 4.5005
R11050 VSS.n8420 VSS.n8328 4.5005
R11051 VSS.n8399 VSS.n8338 4.5005
R11052 VSS.n8399 VSS.n8398 4.5005
R11053 VSS.n8385 VSS.n8351 4.5005
R11054 VSS.n8317 VSS.n8313 4.5005
R11055 VSS.n8315 VSS.n8313 4.5005
R11056 VSS.n8464 VSS.n8463 4.5005
R11057 VSS.n8463 VSS.n8462 4.5005
R11058 VSS.n8820 VSS.n8815 4.5005
R11059 VSS.n9148 VSS.n9147 4.5005
R11060 VSS.n9125 VSS.n8830 4.5005
R11061 VSS.n8858 VSS.n8856 4.5005
R11062 VSS.n9064 VSS.n9062 4.5005
R11063 VSS.n9063 VSS.n8863 4.5005
R11064 VSS.n9066 VSS.n9065 4.5005
R11065 VSS.n9124 VSS.n9123 4.5005
R11066 VSS.n8832 VSS.n8819 4.5005
R11067 VSS.n9114 VSS.n9113 4.5005
R11068 VSS.n8841 VSS.n8839 4.5005
R11069 VSS.n8853 VSS.n8852 4.5005
R11070 VSS.n9086 VSS.n9085 4.5005
R11071 VSS.n8865 VSS.n8855 4.5005
R11072 VSS.n9115 VSS.n8834 4.5005
R11073 VSS.n9146 VSS.n8814 4.5005
R11074 VSS.n9060 VSS.n9059 4.5005
R11075 VSS.n8822 VSS.n8821 4.5005
R11076 VSS.n9135 VSS.n8822 4.5005
R11077 VSS.n8851 VSS.n8849 4.5005
R11078 VSS.n8849 VSS.n8848 4.5005
R11079 VSS.n9075 VSS.n8864 4.5005
R11080 VSS.n9127 VSS.n9126 4.5005
R11081 VSS.n9127 VSS.n8828 4.5005
R11082 VSS.n9182 VSS.n9181 4.5005
R11083 VSS.n9181 VSS.n9180 4.5005
R11084 VSS.n9305 VSS.n8745 4.5005
R11085 VSS.n9246 VSS.n8772 4.5005
R11086 VSS.n9209 VSS.n9208 4.5005
R11087 VSS.n9159 VSS.n9157 4.5005
R11088 VSS.n9188 VSS.n9187 4.5005
R11089 VSS.n9199 VSS.n9198 4.5005
R11090 VSS.n9200 VSS.n9199 4.5005
R11091 VSS.n9233 VSS.n9232 4.5005
R11092 VSS.n9206 VSS.n9205 4.5005
R11093 VSS.n8781 VSS.n8780 4.5005
R11094 VSS.n8790 VSS.n8781 4.5005
R11095 VSS.n9300 VSS.n9299 4.5005
R11096 VSS.n9273 VSS.n8761 4.5005
R11097 VSS.n9273 VSS.n8755 4.5005
R11098 VSS.n9280 VSS.n8757 4.5005
R11099 VSS.n9251 VSS.n9247 4.5005
R11100 VSS.n9251 VSS.n9250 4.5005
R11101 VSS.n9254 VSS.n9245 4.5005
R11102 VSS.n9238 VSS.n9237 4.5005
R11103 VSS.n9237 VSS.n8767 4.5005
R11104 VSS.n9304 VSS.n9303 4.5005
R11105 VSS.n8746 VSS.n8744 4.5005
R11106 VSS.n8744 VSS.n8743 4.5005
R11107 VSS.n9261 VSS.n9260 4.5005
R11108 VSS.n9262 VSS.n9261 4.5005
R11109 VSS.n8758 VSS.n8756 4.5005
R11110 VSS.n9319 VSS.n9318 4.5005
R11111 VSS.n9190 VSS.n9189 4.5005
R11112 VSS.n9191 VSS.n8801 4.5005
R11113 VSS.n9042 VSS.n8889 4.5005
R11114 VSS.n9041 VSS.n9040 4.5005
R11115 VSS.n8911 VSS.n8910 4.5005
R11116 VSS.n8993 VSS.n8992 4.5005
R11117 VSS.n8966 VSS.n8964 4.5005
R11118 VSS.n8965 VSS.n8942 4.5005
R11119 VSS.n8968 VSS.n8967 4.5005
R11120 VSS.n8900 VSS.n8899 4.5005
R11121 VSS.n9031 VSS.n9030 4.5005
R11122 VSS.n8923 VSS.n8922 4.5005
R11123 VSS.n9002 VSS.n9001 4.5005
R11124 VSS.n9000 VSS.n8999 4.5005
R11125 VSS.n8945 VSS.n8929 4.5005
R11126 VSS.n8904 VSS.n8902 4.5005
R11127 VSS.n9039 VSS.n8891 4.5005
R11128 VSS.n8962 VSS.n8961 4.5005
R11129 VSS.n9044 VSS.n9043 4.5005
R11130 VSS.n9044 VSS.n8887 4.5005
R11131 VSS.n9012 VSS.n8920 4.5005
R11132 VSS.n8991 VSS.n8930 4.5005
R11133 VSS.n8991 VSS.n8990 4.5005
R11134 VSS.n8977 VSS.n8943 4.5005
R11135 VSS.n8909 VSS.n8905 4.5005
R11136 VSS.n8907 VSS.n8905 4.5005
R11137 VSS.n9056 VSS.n9055 4.5005
R11138 VSS.n9055 VSS.n9054 4.5005
R11139 VSS.n10004 VSS.n9999 4.5005
R11140 VSS.n10332 VSS.n10331 4.5005
R11141 VSS.n10309 VSS.n10014 4.5005
R11142 VSS.n10042 VSS.n10040 4.5005
R11143 VSS.n10248 VSS.n10246 4.5005
R11144 VSS.n10247 VSS.n10047 4.5005
R11145 VSS.n10250 VSS.n10249 4.5005
R11146 VSS.n10308 VSS.n10307 4.5005
R11147 VSS.n10016 VSS.n10003 4.5005
R11148 VSS.n10298 VSS.n10297 4.5005
R11149 VSS.n10025 VSS.n10023 4.5005
R11150 VSS.n10037 VSS.n10036 4.5005
R11151 VSS.n10270 VSS.n10269 4.5005
R11152 VSS.n10049 VSS.n10039 4.5005
R11153 VSS.n10299 VSS.n10018 4.5005
R11154 VSS.n10330 VSS.n9998 4.5005
R11155 VSS.n10244 VSS.n10243 4.5005
R11156 VSS.n10006 VSS.n10005 4.5005
R11157 VSS.n10319 VSS.n10006 4.5005
R11158 VSS.n10035 VSS.n10033 4.5005
R11159 VSS.n10033 VSS.n10032 4.5005
R11160 VSS.n10259 VSS.n10048 4.5005
R11161 VSS.n10311 VSS.n10310 4.5005
R11162 VSS.n10311 VSS.n10012 4.5005
R11163 VSS.n10366 VSS.n10365 4.5005
R11164 VSS.n10365 VSS.n10364 4.5005
R11165 VSS.n10489 VSS.n9929 4.5005
R11166 VSS.n10430 VSS.n9956 4.5005
R11167 VSS.n10393 VSS.n10392 4.5005
R11168 VSS.n10343 VSS.n10341 4.5005
R11169 VSS.n10372 VSS.n10371 4.5005
R11170 VSS.n10383 VSS.n10382 4.5005
R11171 VSS.n10384 VSS.n10383 4.5005
R11172 VSS.n10417 VSS.n10416 4.5005
R11173 VSS.n10390 VSS.n10389 4.5005
R11174 VSS.n9965 VSS.n9964 4.5005
R11175 VSS.n9974 VSS.n9965 4.5005
R11176 VSS.n10484 VSS.n10483 4.5005
R11177 VSS.n10457 VSS.n9945 4.5005
R11178 VSS.n10457 VSS.n9939 4.5005
R11179 VSS.n10464 VSS.n9941 4.5005
R11180 VSS.n10435 VSS.n10431 4.5005
R11181 VSS.n10435 VSS.n10434 4.5005
R11182 VSS.n10438 VSS.n10429 4.5005
R11183 VSS.n10422 VSS.n10421 4.5005
R11184 VSS.n10421 VSS.n9951 4.5005
R11185 VSS.n10488 VSS.n10487 4.5005
R11186 VSS.n9930 VSS.n9928 4.5005
R11187 VSS.n9928 VSS.n9927 4.5005
R11188 VSS.n10445 VSS.n10444 4.5005
R11189 VSS.n10446 VSS.n10445 4.5005
R11190 VSS.n9942 VSS.n9940 4.5005
R11191 VSS.n10503 VSS.n10502 4.5005
R11192 VSS.n10374 VSS.n10373 4.5005
R11193 VSS.n10375 VSS.n9985 4.5005
R11194 VSS.n10226 VSS.n10073 4.5005
R11195 VSS.n10225 VSS.n10224 4.5005
R11196 VSS.n10095 VSS.n10094 4.5005
R11197 VSS.n10177 VSS.n10176 4.5005
R11198 VSS.n10150 VSS.n10148 4.5005
R11199 VSS.n10149 VSS.n10126 4.5005
R11200 VSS.n10152 VSS.n10151 4.5005
R11201 VSS.n10084 VSS.n10083 4.5005
R11202 VSS.n10215 VSS.n10214 4.5005
R11203 VSS.n10107 VSS.n10106 4.5005
R11204 VSS.n10186 VSS.n10185 4.5005
R11205 VSS.n10184 VSS.n10183 4.5005
R11206 VSS.n10129 VSS.n10113 4.5005
R11207 VSS.n10088 VSS.n10086 4.5005
R11208 VSS.n10223 VSS.n10075 4.5005
R11209 VSS.n10146 VSS.n10145 4.5005
R11210 VSS.n10228 VSS.n10227 4.5005
R11211 VSS.n10228 VSS.n10071 4.5005
R11212 VSS.n10196 VSS.n10104 4.5005
R11213 VSS.n10175 VSS.n10114 4.5005
R11214 VSS.n10175 VSS.n10174 4.5005
R11215 VSS.n10161 VSS.n10127 4.5005
R11216 VSS.n10093 VSS.n10089 4.5005
R11217 VSS.n10091 VSS.n10089 4.5005
R11218 VSS.n10240 VSS.n10239 4.5005
R11219 VSS.n10239 VSS.n10238 4.5005
R11220 VSS.n10596 VSS.n10591 4.5005
R11221 VSS.n10924 VSS.n10923 4.5005
R11222 VSS.n10901 VSS.n10606 4.5005
R11223 VSS.n10634 VSS.n10632 4.5005
R11224 VSS.n10840 VSS.n10838 4.5005
R11225 VSS.n10839 VSS.n10639 4.5005
R11226 VSS.n10842 VSS.n10841 4.5005
R11227 VSS.n10900 VSS.n10899 4.5005
R11228 VSS.n10608 VSS.n10595 4.5005
R11229 VSS.n10890 VSS.n10889 4.5005
R11230 VSS.n10617 VSS.n10615 4.5005
R11231 VSS.n10629 VSS.n10628 4.5005
R11232 VSS.n10862 VSS.n10861 4.5005
R11233 VSS.n10641 VSS.n10631 4.5005
R11234 VSS.n10891 VSS.n10610 4.5005
R11235 VSS.n10922 VSS.n10590 4.5005
R11236 VSS.n10836 VSS.n10835 4.5005
R11237 VSS.n10598 VSS.n10597 4.5005
R11238 VSS.n10911 VSS.n10598 4.5005
R11239 VSS.n10627 VSS.n10625 4.5005
R11240 VSS.n10625 VSS.n10624 4.5005
R11241 VSS.n10851 VSS.n10640 4.5005
R11242 VSS.n10903 VSS.n10902 4.5005
R11243 VSS.n10903 VSS.n10604 4.5005
R11244 VSS.n10958 VSS.n10957 4.5005
R11245 VSS.n10957 VSS.n10956 4.5005
R11246 VSS.n11081 VSS.n10521 4.5005
R11247 VSS.n11022 VSS.n10548 4.5005
R11248 VSS.n10985 VSS.n10984 4.5005
R11249 VSS.n10935 VSS.n10933 4.5005
R11250 VSS.n10964 VSS.n10963 4.5005
R11251 VSS.n10975 VSS.n10974 4.5005
R11252 VSS.n10976 VSS.n10975 4.5005
R11253 VSS.n11009 VSS.n11008 4.5005
R11254 VSS.n10982 VSS.n10981 4.5005
R11255 VSS.n10557 VSS.n10556 4.5005
R11256 VSS.n10566 VSS.n10557 4.5005
R11257 VSS.n11076 VSS.n11075 4.5005
R11258 VSS.n11049 VSS.n10537 4.5005
R11259 VSS.n11049 VSS.n10531 4.5005
R11260 VSS.n11056 VSS.n10533 4.5005
R11261 VSS.n11027 VSS.n11023 4.5005
R11262 VSS.n11027 VSS.n11026 4.5005
R11263 VSS.n11030 VSS.n11021 4.5005
R11264 VSS.n11014 VSS.n11013 4.5005
R11265 VSS.n11013 VSS.n10543 4.5005
R11266 VSS.n11080 VSS.n11079 4.5005
R11267 VSS.n10522 VSS.n10520 4.5005
R11268 VSS.n10520 VSS.n10519 4.5005
R11269 VSS.n11037 VSS.n11036 4.5005
R11270 VSS.n11038 VSS.n11037 4.5005
R11271 VSS.n10534 VSS.n10532 4.5005
R11272 VSS.n11095 VSS.n11094 4.5005
R11273 VSS.n10966 VSS.n10965 4.5005
R11274 VSS.n10967 VSS.n10577 4.5005
R11275 VSS.n10818 VSS.n10665 4.5005
R11276 VSS.n10817 VSS.n10816 4.5005
R11277 VSS.n10687 VSS.n10686 4.5005
R11278 VSS.n10769 VSS.n10768 4.5005
R11279 VSS.n10742 VSS.n10740 4.5005
R11280 VSS.n10741 VSS.n10718 4.5005
R11281 VSS.n10744 VSS.n10743 4.5005
R11282 VSS.n10676 VSS.n10675 4.5005
R11283 VSS.n10807 VSS.n10806 4.5005
R11284 VSS.n10699 VSS.n10698 4.5005
R11285 VSS.n10778 VSS.n10777 4.5005
R11286 VSS.n10776 VSS.n10775 4.5005
R11287 VSS.n10721 VSS.n10705 4.5005
R11288 VSS.n10680 VSS.n10678 4.5005
R11289 VSS.n10815 VSS.n10667 4.5005
R11290 VSS.n10738 VSS.n10737 4.5005
R11291 VSS.n10820 VSS.n10819 4.5005
R11292 VSS.n10820 VSS.n10663 4.5005
R11293 VSS.n10788 VSS.n10696 4.5005
R11294 VSS.n10767 VSS.n10706 4.5005
R11295 VSS.n10767 VSS.n10766 4.5005
R11296 VSS.n10753 VSS.n10719 4.5005
R11297 VSS.n10685 VSS.n10681 4.5005
R11298 VSS.n10683 VSS.n10681 4.5005
R11299 VSS.n10832 VSS.n10831 4.5005
R11300 VSS.n10831 VSS.n10830 4.5005
R11301 VSS.n11188 VSS.n11183 4.5005
R11302 VSS.n11516 VSS.n11515 4.5005
R11303 VSS.n11493 VSS.n11198 4.5005
R11304 VSS.n11226 VSS.n11224 4.5005
R11305 VSS.n11432 VSS.n11430 4.5005
R11306 VSS.n11431 VSS.n11231 4.5005
R11307 VSS.n11434 VSS.n11433 4.5005
R11308 VSS.n11492 VSS.n11491 4.5005
R11309 VSS.n11200 VSS.n11187 4.5005
R11310 VSS.n11482 VSS.n11481 4.5005
R11311 VSS.n11209 VSS.n11207 4.5005
R11312 VSS.n11221 VSS.n11220 4.5005
R11313 VSS.n11454 VSS.n11453 4.5005
R11314 VSS.n11233 VSS.n11223 4.5005
R11315 VSS.n11483 VSS.n11202 4.5005
R11316 VSS.n11514 VSS.n11182 4.5005
R11317 VSS.n11428 VSS.n11427 4.5005
R11318 VSS.n11190 VSS.n11189 4.5005
R11319 VSS.n11503 VSS.n11190 4.5005
R11320 VSS.n11219 VSS.n11217 4.5005
R11321 VSS.n11217 VSS.n11216 4.5005
R11322 VSS.n11443 VSS.n11232 4.5005
R11323 VSS.n11495 VSS.n11494 4.5005
R11324 VSS.n11495 VSS.n11196 4.5005
R11325 VSS.n11550 VSS.n11549 4.5005
R11326 VSS.n11549 VSS.n11548 4.5005
R11327 VSS.n11673 VSS.n11113 4.5005
R11328 VSS.n11614 VSS.n11140 4.5005
R11329 VSS.n11577 VSS.n11576 4.5005
R11330 VSS.n11527 VSS.n11525 4.5005
R11331 VSS.n11556 VSS.n11555 4.5005
R11332 VSS.n11567 VSS.n11566 4.5005
R11333 VSS.n11568 VSS.n11567 4.5005
R11334 VSS.n11601 VSS.n11600 4.5005
R11335 VSS.n11574 VSS.n11573 4.5005
R11336 VSS.n11149 VSS.n11148 4.5005
R11337 VSS.n11158 VSS.n11149 4.5005
R11338 VSS.n11668 VSS.n11667 4.5005
R11339 VSS.n11641 VSS.n11129 4.5005
R11340 VSS.n11641 VSS.n11123 4.5005
R11341 VSS.n11648 VSS.n11125 4.5005
R11342 VSS.n11619 VSS.n11615 4.5005
R11343 VSS.n11619 VSS.n11618 4.5005
R11344 VSS.n11622 VSS.n11613 4.5005
R11345 VSS.n11606 VSS.n11605 4.5005
R11346 VSS.n11605 VSS.n11135 4.5005
R11347 VSS.n11672 VSS.n11671 4.5005
R11348 VSS.n11114 VSS.n11112 4.5005
R11349 VSS.n11112 VSS.n11111 4.5005
R11350 VSS.n11629 VSS.n11628 4.5005
R11351 VSS.n11630 VSS.n11629 4.5005
R11352 VSS.n11126 VSS.n11124 4.5005
R11353 VSS.n11687 VSS.n11686 4.5005
R11354 VSS.n11558 VSS.n11557 4.5005
R11355 VSS.n11559 VSS.n11169 4.5005
R11356 VSS.n11410 VSS.n11257 4.5005
R11357 VSS.n11409 VSS.n11408 4.5005
R11358 VSS.n11279 VSS.n11278 4.5005
R11359 VSS.n11361 VSS.n11360 4.5005
R11360 VSS.n11334 VSS.n11332 4.5005
R11361 VSS.n11333 VSS.n11310 4.5005
R11362 VSS.n11336 VSS.n11335 4.5005
R11363 VSS.n11268 VSS.n11267 4.5005
R11364 VSS.n11399 VSS.n11398 4.5005
R11365 VSS.n11291 VSS.n11290 4.5005
R11366 VSS.n11370 VSS.n11369 4.5005
R11367 VSS.n11368 VSS.n11367 4.5005
R11368 VSS.n11313 VSS.n11297 4.5005
R11369 VSS.n11272 VSS.n11270 4.5005
R11370 VSS.n11407 VSS.n11259 4.5005
R11371 VSS.n11330 VSS.n11329 4.5005
R11372 VSS.n11412 VSS.n11411 4.5005
R11373 VSS.n11412 VSS.n11255 4.5005
R11374 VSS.n11380 VSS.n11288 4.5005
R11375 VSS.n11359 VSS.n11298 4.5005
R11376 VSS.n11359 VSS.n11358 4.5005
R11377 VSS.n11345 VSS.n11311 4.5005
R11378 VSS.n11277 VSS.n11273 4.5005
R11379 VSS.n11275 VSS.n11273 4.5005
R11380 VSS.n11424 VSS.n11423 4.5005
R11381 VSS.n11423 VSS.n11422 4.5005
R11382 VSS.n11780 VSS.n11775 4.5005
R11383 VSS.n12108 VSS.n12107 4.5005
R11384 VSS.n12085 VSS.n11790 4.5005
R11385 VSS.n11818 VSS.n11816 4.5005
R11386 VSS.n12024 VSS.n12022 4.5005
R11387 VSS.n12023 VSS.n11823 4.5005
R11388 VSS.n12026 VSS.n12025 4.5005
R11389 VSS.n12084 VSS.n12083 4.5005
R11390 VSS.n11792 VSS.n11779 4.5005
R11391 VSS.n12074 VSS.n12073 4.5005
R11392 VSS.n11801 VSS.n11799 4.5005
R11393 VSS.n11813 VSS.n11812 4.5005
R11394 VSS.n12046 VSS.n12045 4.5005
R11395 VSS.n11825 VSS.n11815 4.5005
R11396 VSS.n12075 VSS.n11794 4.5005
R11397 VSS.n12106 VSS.n11774 4.5005
R11398 VSS.n12020 VSS.n12019 4.5005
R11399 VSS.n11782 VSS.n11781 4.5005
R11400 VSS.n12095 VSS.n11782 4.5005
R11401 VSS.n11811 VSS.n11809 4.5005
R11402 VSS.n11809 VSS.n11808 4.5005
R11403 VSS.n12035 VSS.n11824 4.5005
R11404 VSS.n12087 VSS.n12086 4.5005
R11405 VSS.n12087 VSS.n11788 4.5005
R11406 VSS.n12142 VSS.n12141 4.5005
R11407 VSS.n12141 VSS.n12140 4.5005
R11408 VSS.n12265 VSS.n11705 4.5005
R11409 VSS.n12206 VSS.n11732 4.5005
R11410 VSS.n12169 VSS.n12168 4.5005
R11411 VSS.n12119 VSS.n12117 4.5005
R11412 VSS.n12148 VSS.n12147 4.5005
R11413 VSS.n12159 VSS.n12158 4.5005
R11414 VSS.n12160 VSS.n12159 4.5005
R11415 VSS.n12193 VSS.n12192 4.5005
R11416 VSS.n12166 VSS.n12165 4.5005
R11417 VSS.n11741 VSS.n11740 4.5005
R11418 VSS.n11750 VSS.n11741 4.5005
R11419 VSS.n12260 VSS.n12259 4.5005
R11420 VSS.n12233 VSS.n11721 4.5005
R11421 VSS.n12233 VSS.n11715 4.5005
R11422 VSS.n12240 VSS.n11717 4.5005
R11423 VSS.n12211 VSS.n12207 4.5005
R11424 VSS.n12211 VSS.n12210 4.5005
R11425 VSS.n12214 VSS.n12205 4.5005
R11426 VSS.n12198 VSS.n12197 4.5005
R11427 VSS.n12197 VSS.n11727 4.5005
R11428 VSS.n12264 VSS.n12263 4.5005
R11429 VSS.n11706 VSS.n11704 4.5005
R11430 VSS.n11704 VSS.n11703 4.5005
R11431 VSS.n12221 VSS.n12220 4.5005
R11432 VSS.n12222 VSS.n12221 4.5005
R11433 VSS.n11718 VSS.n11716 4.5005
R11434 VSS.n12279 VSS.n12278 4.5005
R11435 VSS.n12150 VSS.n12149 4.5005
R11436 VSS.n12151 VSS.n11761 4.5005
R11437 VSS.n12002 VSS.n11849 4.5005
R11438 VSS.n12001 VSS.n12000 4.5005
R11439 VSS.n11871 VSS.n11870 4.5005
R11440 VSS.n11953 VSS.n11952 4.5005
R11441 VSS.n11926 VSS.n11924 4.5005
R11442 VSS.n11925 VSS.n11902 4.5005
R11443 VSS.n11928 VSS.n11927 4.5005
R11444 VSS.n11860 VSS.n11859 4.5005
R11445 VSS.n11991 VSS.n11990 4.5005
R11446 VSS.n11883 VSS.n11882 4.5005
R11447 VSS.n11962 VSS.n11961 4.5005
R11448 VSS.n11960 VSS.n11959 4.5005
R11449 VSS.n11905 VSS.n11889 4.5005
R11450 VSS.n11864 VSS.n11862 4.5005
R11451 VSS.n11999 VSS.n11851 4.5005
R11452 VSS.n11922 VSS.n11921 4.5005
R11453 VSS.n12004 VSS.n12003 4.5005
R11454 VSS.n12004 VSS.n11847 4.5005
R11455 VSS.n11972 VSS.n11880 4.5005
R11456 VSS.n11951 VSS.n11890 4.5005
R11457 VSS.n11951 VSS.n11950 4.5005
R11458 VSS.n11937 VSS.n11903 4.5005
R11459 VSS.n11869 VSS.n11865 4.5005
R11460 VSS.n11867 VSS.n11865 4.5005
R11461 VSS.n12016 VSS.n12015 4.5005
R11462 VSS.n12015 VSS.n12014 4.5005
R11463 VSS.n12372 VSS.n12367 4.5005
R11464 VSS.n12700 VSS.n12699 4.5005
R11465 VSS.n12677 VSS.n12382 4.5005
R11466 VSS.n12410 VSS.n12408 4.5005
R11467 VSS.n12616 VSS.n12614 4.5005
R11468 VSS.n12615 VSS.n12415 4.5005
R11469 VSS.n12618 VSS.n12617 4.5005
R11470 VSS.n12676 VSS.n12675 4.5005
R11471 VSS.n12384 VSS.n12371 4.5005
R11472 VSS.n12666 VSS.n12665 4.5005
R11473 VSS.n12393 VSS.n12391 4.5005
R11474 VSS.n12405 VSS.n12404 4.5005
R11475 VSS.n12638 VSS.n12637 4.5005
R11476 VSS.n12417 VSS.n12407 4.5005
R11477 VSS.n12667 VSS.n12386 4.5005
R11478 VSS.n12698 VSS.n12366 4.5005
R11479 VSS.n12612 VSS.n12611 4.5005
R11480 VSS.n12374 VSS.n12373 4.5005
R11481 VSS.n12687 VSS.n12374 4.5005
R11482 VSS.n12403 VSS.n12401 4.5005
R11483 VSS.n12401 VSS.n12400 4.5005
R11484 VSS.n12627 VSS.n12416 4.5005
R11485 VSS.n12679 VSS.n12678 4.5005
R11486 VSS.n12679 VSS.n12380 4.5005
R11487 VSS.n12734 VSS.n12733 4.5005
R11488 VSS.n12733 VSS.n12732 4.5005
R11489 VSS.n12857 VSS.n12297 4.5005
R11490 VSS.n12798 VSS.n12324 4.5005
R11491 VSS.n12761 VSS.n12760 4.5005
R11492 VSS.n12711 VSS.n12709 4.5005
R11493 VSS.n12740 VSS.n12739 4.5005
R11494 VSS.n12751 VSS.n12750 4.5005
R11495 VSS.n12752 VSS.n12751 4.5005
R11496 VSS.n12785 VSS.n12784 4.5005
R11497 VSS.n12758 VSS.n12757 4.5005
R11498 VSS.n12333 VSS.n12332 4.5005
R11499 VSS.n12342 VSS.n12333 4.5005
R11500 VSS.n12852 VSS.n12851 4.5005
R11501 VSS.n12825 VSS.n12313 4.5005
R11502 VSS.n12825 VSS.n12307 4.5005
R11503 VSS.n12832 VSS.n12309 4.5005
R11504 VSS.n12803 VSS.n12799 4.5005
R11505 VSS.n12803 VSS.n12802 4.5005
R11506 VSS.n12806 VSS.n12797 4.5005
R11507 VSS.n12790 VSS.n12789 4.5005
R11508 VSS.n12789 VSS.n12319 4.5005
R11509 VSS.n12856 VSS.n12855 4.5005
R11510 VSS.n12298 VSS.n12296 4.5005
R11511 VSS.n12296 VSS.n12295 4.5005
R11512 VSS.n12813 VSS.n12812 4.5005
R11513 VSS.n12814 VSS.n12813 4.5005
R11514 VSS.n12310 VSS.n12308 4.5005
R11515 VSS.n12871 VSS.n12870 4.5005
R11516 VSS.n12742 VSS.n12741 4.5005
R11517 VSS.n12743 VSS.n12353 4.5005
R11518 VSS.n12594 VSS.n12441 4.5005
R11519 VSS.n12593 VSS.n12592 4.5005
R11520 VSS.n12463 VSS.n12462 4.5005
R11521 VSS.n12545 VSS.n12544 4.5005
R11522 VSS.n12518 VSS.n12516 4.5005
R11523 VSS.n12517 VSS.n12494 4.5005
R11524 VSS.n12520 VSS.n12519 4.5005
R11525 VSS.n12452 VSS.n12451 4.5005
R11526 VSS.n12583 VSS.n12582 4.5005
R11527 VSS.n12475 VSS.n12474 4.5005
R11528 VSS.n12554 VSS.n12553 4.5005
R11529 VSS.n12552 VSS.n12551 4.5005
R11530 VSS.n12497 VSS.n12481 4.5005
R11531 VSS.n12456 VSS.n12454 4.5005
R11532 VSS.n12591 VSS.n12443 4.5005
R11533 VSS.n12514 VSS.n12513 4.5005
R11534 VSS.n12596 VSS.n12595 4.5005
R11535 VSS.n12596 VSS.n12439 4.5005
R11536 VSS.n12564 VSS.n12472 4.5005
R11537 VSS.n12543 VSS.n12482 4.5005
R11538 VSS.n12543 VSS.n12542 4.5005
R11539 VSS.n12529 VSS.n12495 4.5005
R11540 VSS.n12461 VSS.n12457 4.5005
R11541 VSS.n12459 VSS.n12457 4.5005
R11542 VSS.n12608 VSS.n12607 4.5005
R11543 VSS.n12607 VSS.n12606 4.5005
R11544 VSS.n12964 VSS.n12959 4.5005
R11545 VSS.n13292 VSS.n13291 4.5005
R11546 VSS.n13269 VSS.n12974 4.5005
R11547 VSS.n13002 VSS.n13000 4.5005
R11548 VSS.n13208 VSS.n13206 4.5005
R11549 VSS.n13207 VSS.n13007 4.5005
R11550 VSS.n13210 VSS.n13209 4.5005
R11551 VSS.n13268 VSS.n13267 4.5005
R11552 VSS.n12976 VSS.n12963 4.5005
R11553 VSS.n13258 VSS.n13257 4.5005
R11554 VSS.n12985 VSS.n12983 4.5005
R11555 VSS.n12997 VSS.n12996 4.5005
R11556 VSS.n13230 VSS.n13229 4.5005
R11557 VSS.n13009 VSS.n12999 4.5005
R11558 VSS.n13259 VSS.n12978 4.5005
R11559 VSS.n13290 VSS.n12958 4.5005
R11560 VSS.n13204 VSS.n13203 4.5005
R11561 VSS.n12966 VSS.n12965 4.5005
R11562 VSS.n13279 VSS.n12966 4.5005
R11563 VSS.n12995 VSS.n12993 4.5005
R11564 VSS.n12993 VSS.n12992 4.5005
R11565 VSS.n13219 VSS.n13008 4.5005
R11566 VSS.n13271 VSS.n13270 4.5005
R11567 VSS.n13271 VSS.n12972 4.5005
R11568 VSS.n13326 VSS.n13325 4.5005
R11569 VSS.n13325 VSS.n13324 4.5005
R11570 VSS.n13449 VSS.n12889 4.5005
R11571 VSS.n13390 VSS.n12916 4.5005
R11572 VSS.n13353 VSS.n13352 4.5005
R11573 VSS.n13303 VSS.n13301 4.5005
R11574 VSS.n13332 VSS.n13331 4.5005
R11575 VSS.n13343 VSS.n13342 4.5005
R11576 VSS.n13344 VSS.n13343 4.5005
R11577 VSS.n13377 VSS.n13376 4.5005
R11578 VSS.n13350 VSS.n13349 4.5005
R11579 VSS.n12925 VSS.n12924 4.5005
R11580 VSS.n12934 VSS.n12925 4.5005
R11581 VSS.n13444 VSS.n13443 4.5005
R11582 VSS.n13417 VSS.n12905 4.5005
R11583 VSS.n13417 VSS.n12899 4.5005
R11584 VSS.n13424 VSS.n12901 4.5005
R11585 VSS.n13395 VSS.n13391 4.5005
R11586 VSS.n13395 VSS.n13394 4.5005
R11587 VSS.n13398 VSS.n13389 4.5005
R11588 VSS.n13382 VSS.n13381 4.5005
R11589 VSS.n13381 VSS.n12911 4.5005
R11590 VSS.n13448 VSS.n13447 4.5005
R11591 VSS.n12890 VSS.n12888 4.5005
R11592 VSS.n12888 VSS.n12887 4.5005
R11593 VSS.n13405 VSS.n13404 4.5005
R11594 VSS.n13406 VSS.n13405 4.5005
R11595 VSS.n12902 VSS.n12900 4.5005
R11596 VSS.n13463 VSS.n13462 4.5005
R11597 VSS.n13334 VSS.n13333 4.5005
R11598 VSS.n13335 VSS.n12945 4.5005
R11599 VSS.n13186 VSS.n13033 4.5005
R11600 VSS.n13185 VSS.n13184 4.5005
R11601 VSS.n13055 VSS.n13054 4.5005
R11602 VSS.n13137 VSS.n13136 4.5005
R11603 VSS.n13110 VSS.n13108 4.5005
R11604 VSS.n13109 VSS.n13086 4.5005
R11605 VSS.n13112 VSS.n13111 4.5005
R11606 VSS.n13044 VSS.n13043 4.5005
R11607 VSS.n13175 VSS.n13174 4.5005
R11608 VSS.n13067 VSS.n13066 4.5005
R11609 VSS.n13146 VSS.n13145 4.5005
R11610 VSS.n13144 VSS.n13143 4.5005
R11611 VSS.n13089 VSS.n13073 4.5005
R11612 VSS.n13048 VSS.n13046 4.5005
R11613 VSS.n13183 VSS.n13035 4.5005
R11614 VSS.n13106 VSS.n13105 4.5005
R11615 VSS.n13188 VSS.n13187 4.5005
R11616 VSS.n13188 VSS.n13031 4.5005
R11617 VSS.n13156 VSS.n13064 4.5005
R11618 VSS.n13135 VSS.n13074 4.5005
R11619 VSS.n13135 VSS.n13134 4.5005
R11620 VSS.n13121 VSS.n13087 4.5005
R11621 VSS.n13053 VSS.n13049 4.5005
R11622 VSS.n13051 VSS.n13049 4.5005
R11623 VSS.n13200 VSS.n13199 4.5005
R11624 VSS.n13199 VSS.n13198 4.5005
R11625 VSS.n13556 VSS.n13551 4.5005
R11626 VSS.n13884 VSS.n13883 4.5005
R11627 VSS.n13861 VSS.n13566 4.5005
R11628 VSS.n13594 VSS.n13592 4.5005
R11629 VSS.n13800 VSS.n13798 4.5005
R11630 VSS.n13799 VSS.n13599 4.5005
R11631 VSS.n13802 VSS.n13801 4.5005
R11632 VSS.n13860 VSS.n13859 4.5005
R11633 VSS.n13568 VSS.n13555 4.5005
R11634 VSS.n13850 VSS.n13849 4.5005
R11635 VSS.n13577 VSS.n13575 4.5005
R11636 VSS.n13589 VSS.n13588 4.5005
R11637 VSS.n13822 VSS.n13821 4.5005
R11638 VSS.n13601 VSS.n13591 4.5005
R11639 VSS.n13851 VSS.n13570 4.5005
R11640 VSS.n13882 VSS.n13550 4.5005
R11641 VSS.n13796 VSS.n13795 4.5005
R11642 VSS.n13558 VSS.n13557 4.5005
R11643 VSS.n13871 VSS.n13558 4.5005
R11644 VSS.n13587 VSS.n13585 4.5005
R11645 VSS.n13585 VSS.n13584 4.5005
R11646 VSS.n13811 VSS.n13600 4.5005
R11647 VSS.n13863 VSS.n13862 4.5005
R11648 VSS.n13863 VSS.n13564 4.5005
R11649 VSS.n13918 VSS.n13917 4.5005
R11650 VSS.n13917 VSS.n13916 4.5005
R11651 VSS.n14041 VSS.n13481 4.5005
R11652 VSS.n13982 VSS.n13508 4.5005
R11653 VSS.n13945 VSS.n13944 4.5005
R11654 VSS.n13895 VSS.n13893 4.5005
R11655 VSS.n13924 VSS.n13923 4.5005
R11656 VSS.n13935 VSS.n13934 4.5005
R11657 VSS.n13936 VSS.n13935 4.5005
R11658 VSS.n13969 VSS.n13968 4.5005
R11659 VSS.n13942 VSS.n13941 4.5005
R11660 VSS.n13517 VSS.n13516 4.5005
R11661 VSS.n13526 VSS.n13517 4.5005
R11662 VSS.n14036 VSS.n14035 4.5005
R11663 VSS.n14009 VSS.n13497 4.5005
R11664 VSS.n14009 VSS.n13491 4.5005
R11665 VSS.n14016 VSS.n13493 4.5005
R11666 VSS.n13987 VSS.n13983 4.5005
R11667 VSS.n13987 VSS.n13986 4.5005
R11668 VSS.n13990 VSS.n13981 4.5005
R11669 VSS.n13974 VSS.n13973 4.5005
R11670 VSS.n13973 VSS.n13503 4.5005
R11671 VSS.n14040 VSS.n14039 4.5005
R11672 VSS.n13482 VSS.n13480 4.5005
R11673 VSS.n13480 VSS.n13479 4.5005
R11674 VSS.n13997 VSS.n13996 4.5005
R11675 VSS.n13998 VSS.n13997 4.5005
R11676 VSS.n13494 VSS.n13492 4.5005
R11677 VSS.n14055 VSS.n14054 4.5005
R11678 VSS.n13926 VSS.n13925 4.5005
R11679 VSS.n13927 VSS.n13537 4.5005
R11680 VSS.n13778 VSS.n13625 4.5005
R11681 VSS.n13777 VSS.n13776 4.5005
R11682 VSS.n13647 VSS.n13646 4.5005
R11683 VSS.n13729 VSS.n13728 4.5005
R11684 VSS.n13702 VSS.n13700 4.5005
R11685 VSS.n13701 VSS.n13678 4.5005
R11686 VSS.n13704 VSS.n13703 4.5005
R11687 VSS.n13636 VSS.n13635 4.5005
R11688 VSS.n13767 VSS.n13766 4.5005
R11689 VSS.n13659 VSS.n13658 4.5005
R11690 VSS.n13738 VSS.n13737 4.5005
R11691 VSS.n13736 VSS.n13735 4.5005
R11692 VSS.n13681 VSS.n13665 4.5005
R11693 VSS.n13640 VSS.n13638 4.5005
R11694 VSS.n13775 VSS.n13627 4.5005
R11695 VSS.n13698 VSS.n13697 4.5005
R11696 VSS.n13780 VSS.n13779 4.5005
R11697 VSS.n13780 VSS.n13623 4.5005
R11698 VSS.n13748 VSS.n13656 4.5005
R11699 VSS.n13727 VSS.n13666 4.5005
R11700 VSS.n13727 VSS.n13726 4.5005
R11701 VSS.n13713 VSS.n13679 4.5005
R11702 VSS.n13645 VSS.n13641 4.5005
R11703 VSS.n13643 VSS.n13641 4.5005
R11704 VSS.n13792 VSS.n13791 4.5005
R11705 VSS.n13791 VSS.n13790 4.5005
R11706 VSS.n14148 VSS.n14143 4.5005
R11707 VSS.n14476 VSS.n14475 4.5005
R11708 VSS.n14453 VSS.n14158 4.5005
R11709 VSS.n14186 VSS.n14184 4.5005
R11710 VSS.n14392 VSS.n14390 4.5005
R11711 VSS.n14391 VSS.n14191 4.5005
R11712 VSS.n14394 VSS.n14393 4.5005
R11713 VSS.n14452 VSS.n14451 4.5005
R11714 VSS.n14160 VSS.n14147 4.5005
R11715 VSS.n14442 VSS.n14441 4.5005
R11716 VSS.n14169 VSS.n14167 4.5005
R11717 VSS.n14181 VSS.n14180 4.5005
R11718 VSS.n14414 VSS.n14413 4.5005
R11719 VSS.n14193 VSS.n14183 4.5005
R11720 VSS.n14443 VSS.n14162 4.5005
R11721 VSS.n14474 VSS.n14142 4.5005
R11722 VSS.n14388 VSS.n14387 4.5005
R11723 VSS.n14150 VSS.n14149 4.5005
R11724 VSS.n14463 VSS.n14150 4.5005
R11725 VSS.n14179 VSS.n14177 4.5005
R11726 VSS.n14177 VSS.n14176 4.5005
R11727 VSS.n14403 VSS.n14192 4.5005
R11728 VSS.n14455 VSS.n14454 4.5005
R11729 VSS.n14455 VSS.n14156 4.5005
R11730 VSS.n14510 VSS.n14509 4.5005
R11731 VSS.n14509 VSS.n14508 4.5005
R11732 VSS.n14633 VSS.n14073 4.5005
R11733 VSS.n14574 VSS.n14100 4.5005
R11734 VSS.n14537 VSS.n14536 4.5005
R11735 VSS.n14487 VSS.n14485 4.5005
R11736 VSS.n14516 VSS.n14515 4.5005
R11737 VSS.n14527 VSS.n14526 4.5005
R11738 VSS.n14528 VSS.n14527 4.5005
R11739 VSS.n14561 VSS.n14560 4.5005
R11740 VSS.n14534 VSS.n14533 4.5005
R11741 VSS.n14109 VSS.n14108 4.5005
R11742 VSS.n14118 VSS.n14109 4.5005
R11743 VSS.n14628 VSS.n14627 4.5005
R11744 VSS.n14601 VSS.n14089 4.5005
R11745 VSS.n14601 VSS.n14083 4.5005
R11746 VSS.n14608 VSS.n14085 4.5005
R11747 VSS.n14579 VSS.n14575 4.5005
R11748 VSS.n14579 VSS.n14578 4.5005
R11749 VSS.n14582 VSS.n14573 4.5005
R11750 VSS.n14566 VSS.n14565 4.5005
R11751 VSS.n14565 VSS.n14095 4.5005
R11752 VSS.n14632 VSS.n14631 4.5005
R11753 VSS.n14074 VSS.n14072 4.5005
R11754 VSS.n14072 VSS.n14071 4.5005
R11755 VSS.n14589 VSS.n14588 4.5005
R11756 VSS.n14590 VSS.n14589 4.5005
R11757 VSS.n14086 VSS.n14084 4.5005
R11758 VSS.n14647 VSS.n14646 4.5005
R11759 VSS.n14518 VSS.n14517 4.5005
R11760 VSS.n14519 VSS.n14129 4.5005
R11761 VSS.n14370 VSS.n14217 4.5005
R11762 VSS.n14369 VSS.n14368 4.5005
R11763 VSS.n14239 VSS.n14238 4.5005
R11764 VSS.n14321 VSS.n14320 4.5005
R11765 VSS.n14294 VSS.n14292 4.5005
R11766 VSS.n14293 VSS.n14270 4.5005
R11767 VSS.n14296 VSS.n14295 4.5005
R11768 VSS.n14228 VSS.n14227 4.5005
R11769 VSS.n14359 VSS.n14358 4.5005
R11770 VSS.n14251 VSS.n14250 4.5005
R11771 VSS.n14330 VSS.n14329 4.5005
R11772 VSS.n14328 VSS.n14327 4.5005
R11773 VSS.n14273 VSS.n14257 4.5005
R11774 VSS.n14232 VSS.n14230 4.5005
R11775 VSS.n14367 VSS.n14219 4.5005
R11776 VSS.n14290 VSS.n14289 4.5005
R11777 VSS.n14372 VSS.n14371 4.5005
R11778 VSS.n14372 VSS.n14215 4.5005
R11779 VSS.n14340 VSS.n14248 4.5005
R11780 VSS.n14319 VSS.n14258 4.5005
R11781 VSS.n14319 VSS.n14318 4.5005
R11782 VSS.n14305 VSS.n14271 4.5005
R11783 VSS.n14237 VSS.n14233 4.5005
R11784 VSS.n14235 VSS.n14233 4.5005
R11785 VSS.n14384 VSS.n14383 4.5005
R11786 VSS.n14383 VSS.n14382 4.5005
R11787 VSS.n14740 VSS.n14735 4.5005
R11788 VSS.n15068 VSS.n15067 4.5005
R11789 VSS.n15045 VSS.n14750 4.5005
R11790 VSS.n14778 VSS.n14776 4.5005
R11791 VSS.n14984 VSS.n14982 4.5005
R11792 VSS.n14983 VSS.n14783 4.5005
R11793 VSS.n14986 VSS.n14985 4.5005
R11794 VSS.n15044 VSS.n15043 4.5005
R11795 VSS.n14752 VSS.n14739 4.5005
R11796 VSS.n15034 VSS.n15033 4.5005
R11797 VSS.n14761 VSS.n14759 4.5005
R11798 VSS.n14773 VSS.n14772 4.5005
R11799 VSS.n15006 VSS.n15005 4.5005
R11800 VSS.n14785 VSS.n14775 4.5005
R11801 VSS.n15035 VSS.n14754 4.5005
R11802 VSS.n15066 VSS.n14734 4.5005
R11803 VSS.n14980 VSS.n14979 4.5005
R11804 VSS.n14742 VSS.n14741 4.5005
R11805 VSS.n15055 VSS.n14742 4.5005
R11806 VSS.n14771 VSS.n14769 4.5005
R11807 VSS.n14769 VSS.n14768 4.5005
R11808 VSS.n14995 VSS.n14784 4.5005
R11809 VSS.n15047 VSS.n15046 4.5005
R11810 VSS.n15047 VSS.n14748 4.5005
R11811 VSS.n15102 VSS.n15101 4.5005
R11812 VSS.n15101 VSS.n15100 4.5005
R11813 VSS.n15225 VSS.n14665 4.5005
R11814 VSS.n15166 VSS.n14692 4.5005
R11815 VSS.n15129 VSS.n15128 4.5005
R11816 VSS.n15079 VSS.n15077 4.5005
R11817 VSS.n15108 VSS.n15107 4.5005
R11818 VSS.n15119 VSS.n15118 4.5005
R11819 VSS.n15120 VSS.n15119 4.5005
R11820 VSS.n15153 VSS.n15152 4.5005
R11821 VSS.n15126 VSS.n15125 4.5005
R11822 VSS.n14701 VSS.n14700 4.5005
R11823 VSS.n14710 VSS.n14701 4.5005
R11824 VSS.n15220 VSS.n15219 4.5005
R11825 VSS.n15193 VSS.n14681 4.5005
R11826 VSS.n15193 VSS.n14675 4.5005
R11827 VSS.n15200 VSS.n14677 4.5005
R11828 VSS.n15171 VSS.n15167 4.5005
R11829 VSS.n15171 VSS.n15170 4.5005
R11830 VSS.n15174 VSS.n15165 4.5005
R11831 VSS.n15158 VSS.n15157 4.5005
R11832 VSS.n15157 VSS.n14687 4.5005
R11833 VSS.n15224 VSS.n15223 4.5005
R11834 VSS.n14666 VSS.n14664 4.5005
R11835 VSS.n14664 VSS.n14663 4.5005
R11836 VSS.n15181 VSS.n15180 4.5005
R11837 VSS.n15182 VSS.n15181 4.5005
R11838 VSS.n14678 VSS.n14676 4.5005
R11839 VSS.n15239 VSS.n15238 4.5005
R11840 VSS.n15110 VSS.n15109 4.5005
R11841 VSS.n15111 VSS.n14721 4.5005
R11842 VSS.n14962 VSS.n14809 4.5005
R11843 VSS.n14961 VSS.n14960 4.5005
R11844 VSS.n14831 VSS.n14830 4.5005
R11845 VSS.n14913 VSS.n14912 4.5005
R11846 VSS.n14886 VSS.n14884 4.5005
R11847 VSS.n14885 VSS.n14862 4.5005
R11848 VSS.n14888 VSS.n14887 4.5005
R11849 VSS.n14820 VSS.n14819 4.5005
R11850 VSS.n14951 VSS.n14950 4.5005
R11851 VSS.n14843 VSS.n14842 4.5005
R11852 VSS.n14922 VSS.n14921 4.5005
R11853 VSS.n14920 VSS.n14919 4.5005
R11854 VSS.n14865 VSS.n14849 4.5005
R11855 VSS.n14824 VSS.n14822 4.5005
R11856 VSS.n14959 VSS.n14811 4.5005
R11857 VSS.n14882 VSS.n14881 4.5005
R11858 VSS.n14964 VSS.n14963 4.5005
R11859 VSS.n14964 VSS.n14807 4.5005
R11860 VSS.n14932 VSS.n14840 4.5005
R11861 VSS.n14911 VSS.n14850 4.5005
R11862 VSS.n14911 VSS.n14910 4.5005
R11863 VSS.n14897 VSS.n14863 4.5005
R11864 VSS.n14829 VSS.n14825 4.5005
R11865 VSS.n14827 VSS.n14825 4.5005
R11866 VSS.n14976 VSS.n14975 4.5005
R11867 VSS.n14975 VSS.n14974 4.5005
R11868 VSS.n15332 VSS.n15327 4.5005
R11869 VSS.n15660 VSS.n15659 4.5005
R11870 VSS.n15637 VSS.n15342 4.5005
R11871 VSS.n15370 VSS.n15368 4.5005
R11872 VSS.n15576 VSS.n15574 4.5005
R11873 VSS.n15575 VSS.n15375 4.5005
R11874 VSS.n15578 VSS.n15577 4.5005
R11875 VSS.n15636 VSS.n15635 4.5005
R11876 VSS.n15344 VSS.n15331 4.5005
R11877 VSS.n15626 VSS.n15625 4.5005
R11878 VSS.n15353 VSS.n15351 4.5005
R11879 VSS.n15365 VSS.n15364 4.5005
R11880 VSS.n15598 VSS.n15597 4.5005
R11881 VSS.n15377 VSS.n15367 4.5005
R11882 VSS.n15627 VSS.n15346 4.5005
R11883 VSS.n15658 VSS.n15326 4.5005
R11884 VSS.n15572 VSS.n15571 4.5005
R11885 VSS.n15334 VSS.n15333 4.5005
R11886 VSS.n15647 VSS.n15334 4.5005
R11887 VSS.n15363 VSS.n15361 4.5005
R11888 VSS.n15361 VSS.n15360 4.5005
R11889 VSS.n15587 VSS.n15376 4.5005
R11890 VSS.n15639 VSS.n15638 4.5005
R11891 VSS.n15639 VSS.n15340 4.5005
R11892 VSS.n15694 VSS.n15693 4.5005
R11893 VSS.n15693 VSS.n15692 4.5005
R11894 VSS.n15817 VSS.n15257 4.5005
R11895 VSS.n15758 VSS.n15284 4.5005
R11896 VSS.n15721 VSS.n15720 4.5005
R11897 VSS.n15671 VSS.n15669 4.5005
R11898 VSS.n15700 VSS.n15699 4.5005
R11899 VSS.n15711 VSS.n15710 4.5005
R11900 VSS.n15712 VSS.n15711 4.5005
R11901 VSS.n15745 VSS.n15744 4.5005
R11902 VSS.n15718 VSS.n15717 4.5005
R11903 VSS.n15293 VSS.n15292 4.5005
R11904 VSS.n15302 VSS.n15293 4.5005
R11905 VSS.n15812 VSS.n15811 4.5005
R11906 VSS.n15785 VSS.n15273 4.5005
R11907 VSS.n15785 VSS.n15267 4.5005
R11908 VSS.n15792 VSS.n15269 4.5005
R11909 VSS.n15763 VSS.n15759 4.5005
R11910 VSS.n15763 VSS.n15762 4.5005
R11911 VSS.n15766 VSS.n15757 4.5005
R11912 VSS.n15750 VSS.n15749 4.5005
R11913 VSS.n15749 VSS.n15279 4.5005
R11914 VSS.n15816 VSS.n15815 4.5005
R11915 VSS.n15258 VSS.n15256 4.5005
R11916 VSS.n15256 VSS.n15255 4.5005
R11917 VSS.n15773 VSS.n15772 4.5005
R11918 VSS.n15774 VSS.n15773 4.5005
R11919 VSS.n15270 VSS.n15268 4.5005
R11920 VSS.n15831 VSS.n15830 4.5005
R11921 VSS.n15702 VSS.n15701 4.5005
R11922 VSS.n15703 VSS.n15313 4.5005
R11923 VSS.n15554 VSS.n15401 4.5005
R11924 VSS.n15553 VSS.n15552 4.5005
R11925 VSS.n15423 VSS.n15422 4.5005
R11926 VSS.n15505 VSS.n15504 4.5005
R11927 VSS.n15478 VSS.n15476 4.5005
R11928 VSS.n15477 VSS.n15454 4.5005
R11929 VSS.n15480 VSS.n15479 4.5005
R11930 VSS.n15412 VSS.n15411 4.5005
R11931 VSS.n15543 VSS.n15542 4.5005
R11932 VSS.n15435 VSS.n15434 4.5005
R11933 VSS.n15514 VSS.n15513 4.5005
R11934 VSS.n15512 VSS.n15511 4.5005
R11935 VSS.n15457 VSS.n15441 4.5005
R11936 VSS.n15416 VSS.n15414 4.5005
R11937 VSS.n15551 VSS.n15403 4.5005
R11938 VSS.n15474 VSS.n15473 4.5005
R11939 VSS.n15556 VSS.n15555 4.5005
R11940 VSS.n15556 VSS.n15399 4.5005
R11941 VSS.n15524 VSS.n15432 4.5005
R11942 VSS.n15503 VSS.n15442 4.5005
R11943 VSS.n15503 VSS.n15502 4.5005
R11944 VSS.n15489 VSS.n15455 4.5005
R11945 VSS.n15421 VSS.n15417 4.5005
R11946 VSS.n15419 VSS.n15417 4.5005
R11947 VSS.n15568 VSS.n15567 4.5005
R11948 VSS.n15567 VSS.n15566 4.5005
R11949 VSS.n6796 VSS.n6795 4.5005
R11950 VSS.n6799 VSS.n6798 4.5005
R11951 VSS.n6782 VSS.n6781 4.5005
R11952 VSS.n6757 VSS.n6756 4.5005
R11953 VSS.n6748 VSS.n6747 4.5005
R11954 VSS.n6749 VSS.n6741 4.5005
R11955 VSS.n6745 VSS.n6742 4.5005
R11956 VSS.n6706 VSS.n6704 4.5005
R11957 VSS.n15934 VSS.n15933 4.5005
R11958 VSS.n15941 VSS.n6696 4.5005
R11959 VSS.n15948 VSS.n15947 4.5005
R11960 VSS.n15949 VSS.n6688 4.5005
R11961 VSS.n6753 VSS.n6685 4.5005
R11962 VSS.n15956 VSS.n15955 4.5005
R11963 VSS.n15940 VSS.n15939 4.5005
R11964 VSS.n6797 VSS.n6721 4.5005
R11965 VSS.n15964 VSS.n15963 4.5005
R11966 VSS.n6794 VSS.n6722 4.5005
R11967 VSS.n6794 VSS.n6793 4.5005
R11968 VSS.n6755 VSS.n6754 4.5005
R11969 VSS.n6754 VSS.n6732 4.5005
R11970 VSS.n6751 VSS.n6750 4.5005
R11971 VSS.n6784 VSS.n6783 4.5005
R11972 VSS.n6784 VSS.n6777 4.5005
R11973 VSS.n15926 VSS.n6714 4.5005
R11974 VSS.n15926 VSS.n15925 4.5005
R11975 VSS.n6947 VSS.n6946 4.5005
R11976 VSS.n6917 VSS.n6866 4.5005
R11977 VSS.n15893 VSS.n15892 4.5005
R11978 VSS.n6824 VSS.n6808 4.5005
R11979 VSS.n6832 VSS.n6831 4.5005
R11980 VSS.n15907 VSS.n6816 4.5005
R11981 VSS.n6816 VSS.n6814 4.5005
R11982 VSS.n6879 VSS.n6878 4.5005
R11983 VSS.n6850 VSS.n6849 4.5005
R11984 VSS.n15891 VSS.n6845 4.5005
R11985 VSS.n6845 VSS.n6843 4.5005
R11986 VSS.n6952 VSS.n6936 4.5005
R11987 VSS.n15865 VSS.n15864 4.5005
R11988 VSS.n15866 VSS.n15865 4.5005
R11989 VSS.n15860 VSS.n6897 4.5005
R11990 VSS.n6919 VSS.n6918 4.5005
R11991 VSS.n6919 VSS.n6914 4.5005
R11992 VSS.n15870 VSS.n6890 4.5005
R11993 VSS.n6884 VSS.n6883 4.5005
R11994 VSS.n6883 VSS.n6861 4.5005
R11995 VSS.n6948 VSS.n6944 4.5005
R11996 VSS.n15852 VSS.n6906 4.5005
R11997 VSS.n15852 VSS.n15851 4.5005
R11998 VSS.n15877 VSS.n15876 4.5005
R11999 VSS.n15878 VSS.n15877 4.5005
R12000 VSS.n15863 VSS.n6895 4.5005
R12001 VSS.n6937 VSS.n6935 4.5005
R12002 VSS.n6817 VSS.n6815 4.5005
R12003 VSS.n6833 VSS.n6821 4.5005
R12004 VSS.n6662 VSS.n6509 4.5005
R12005 VSS.n6661 VSS.n6660 4.5005
R12006 VSS.n6531 VSS.n6530 4.5005
R12007 VSS.n6613 VSS.n6612 4.5005
R12008 VSS.n6586 VSS.n6584 4.5005
R12009 VSS.n6585 VSS.n6562 4.5005
R12010 VSS.n6588 VSS.n6587 4.5005
R12011 VSS.n6520 VSS.n6519 4.5005
R12012 VSS.n6651 VSS.n6650 4.5005
R12013 VSS.n6543 VSS.n6542 4.5005
R12014 VSS.n6622 VSS.n6621 4.5005
R12015 VSS.n6620 VSS.n6619 4.5005
R12016 VSS.n6565 VSS.n6549 4.5005
R12017 VSS.n6524 VSS.n6522 4.5005
R12018 VSS.n6659 VSS.n6511 4.5005
R12019 VSS.n6582 VSS.n6581 4.5005
R12020 VSS.n6664 VSS.n6663 4.5005
R12021 VSS.n6664 VSS.n6507 4.5005
R12022 VSS.n6632 VSS.n6540 4.5005
R12023 VSS.n6611 VSS.n6550 4.5005
R12024 VSS.n6611 VSS.n6610 4.5005
R12025 VSS.n6597 VSS.n6563 4.5005
R12026 VSS.n6529 VSS.n6525 4.5005
R12027 VSS.n6527 VSS.n6525 4.5005
R12028 VSS.n6676 VSS.n6675 4.5005
R12029 VSS.n6675 VSS.n6674 4.5005
R12030 VSS.n7043 VSS.n7038 4.5005
R12031 VSS.n7372 VSS.n7371 4.5005
R12032 VSS.n7349 VSS.n7053 4.5005
R12033 VSS.n7081 VSS.n7079 4.5005
R12034 VSS.n7288 VSS.n7286 4.5005
R12035 VSS.n7287 VSS.n7086 4.5005
R12036 VSS.n7290 VSS.n7289 4.5005
R12037 VSS.n7348 VSS.n7347 4.5005
R12038 VSS.n7055 VSS.n7042 4.5005
R12039 VSS.n7338 VSS.n7337 4.5005
R12040 VSS.n7064 VSS.n7062 4.5005
R12041 VSS.n7076 VSS.n7075 4.5005
R12042 VSS.n7310 VSS.n7309 4.5005
R12043 VSS.n7088 VSS.n7078 4.5005
R12044 VSS.n7339 VSS.n7057 4.5005
R12045 VSS.n7370 VSS.n7037 4.5005
R12046 VSS.n7284 VSS.n7283 4.5005
R12047 VSS.n7045 VSS.n7044 4.5005
R12048 VSS.n7359 VSS.n7045 4.5005
R12049 VSS.n7074 VSS.n7072 4.5005
R12050 VSS.n7072 VSS.n7071 4.5005
R12051 VSS.n7299 VSS.n7087 4.5005
R12052 VSS.n7351 VSS.n7350 4.5005
R12053 VSS.n7351 VSS.n7051 4.5005
R12054 VSS.n7406 VSS.n7405 4.5005
R12055 VSS.n7405 VSS.n7404 4.5005
R12056 VSS.n7529 VSS.n6968 4.5005
R12057 VSS.n7470 VSS.n6995 4.5005
R12058 VSS.n7433 VSS.n7432 4.5005
R12059 VSS.n7383 VSS.n7381 4.5005
R12060 VSS.n7412 VSS.n7411 4.5005
R12061 VSS.n7423 VSS.n7422 4.5005
R12062 VSS.n7424 VSS.n7423 4.5005
R12063 VSS.n7457 VSS.n7456 4.5005
R12064 VSS.n7430 VSS.n7429 4.5005
R12065 VSS.n7004 VSS.n7003 4.5005
R12066 VSS.n7013 VSS.n7004 4.5005
R12067 VSS.n7524 VSS.n7523 4.5005
R12068 VSS.n7497 VSS.n6984 4.5005
R12069 VSS.n7497 VSS.n6978 4.5005
R12070 VSS.n7504 VSS.n6980 4.5005
R12071 VSS.n7475 VSS.n7471 4.5005
R12072 VSS.n7475 VSS.n7474 4.5005
R12073 VSS.n7478 VSS.n7469 4.5005
R12074 VSS.n7462 VSS.n7461 4.5005
R12075 VSS.n7461 VSS.n6990 4.5005
R12076 VSS.n7528 VSS.n7527 4.5005
R12077 VSS.n6969 VSS.n6967 4.5005
R12078 VSS.n6967 VSS.n6966 4.5005
R12079 VSS.n7485 VSS.n7484 4.5005
R12080 VSS.n7486 VSS.n7485 4.5005
R12081 VSS.n6981 VSS.n6979 4.5005
R12082 VSS.n7543 VSS.n7542 4.5005
R12083 VSS.n7414 VSS.n7413 4.5005
R12084 VSS.n7415 VSS.n7024 4.5005
R12085 VSS.n7118 VSS.n7113 4.5005
R12086 VSS.n7268 VSS.n7267 4.5005
R12087 VSS.n7244 VSS.n7128 4.5005
R12088 VSS.n7205 VSS.n7204 4.5005
R12089 VSS.n7183 VSS.n7181 4.5005
R12090 VSS.n7182 VSS.n7161 4.5005
R12091 VSS.n7185 VSS.n7184 4.5005
R12092 VSS.n7243 VSS.n7242 4.5005
R12093 VSS.n7130 VSS.n7117 4.5005
R12094 VSS.n7233 VSS.n7232 4.5005
R12095 VSS.n7139 VSS.n7137 4.5005
R12096 VSS.n7153 VSS.n7152 4.5005
R12097 VSS.n7163 VSS.n7155 4.5005
R12098 VSS.n7234 VSS.n7132 4.5005
R12099 VSS.n7266 VSS.n7112 4.5005
R12100 VSS.n7179 VSS.n7178 4.5005
R12101 VSS.n7120 VSS.n7119 4.5005
R12102 VSS.n7255 VSS.n7120 4.5005
R12103 VSS.n7225 VSS.n7138 4.5005
R12104 VSS.n7151 VSS.n7149 4.5005
R12105 VSS.n7149 VSS.n7148 4.5005
R12106 VSS.n7194 VSS.n7162 4.5005
R12107 VSS.n7246 VSS.n7245 4.5005
R12108 VSS.n7246 VSS.n7126 4.5005
R12109 VSS.n7280 VSS.n7279 4.5005
R12110 VSS.n7279 VSS.n7278 4.5005
R12111 VSS.n141 VSS.n136 4.5005
R12112 VSS.n18684 VSS.n18683 4.5005
R12113 VSS.n18661 VSS.n151 4.5005
R12114 VSS.n179 VSS.n177 4.5005
R12115 VSS.n18600 VSS.n18598 4.5005
R12116 VSS.n18599 VSS.n184 4.5005
R12117 VSS.n18602 VSS.n18601 4.5005
R12118 VSS.n18660 VSS.n18659 4.5005
R12119 VSS.n153 VSS.n140 4.5005
R12120 VSS.n18650 VSS.n18649 4.5005
R12121 VSS.n162 VSS.n160 4.5005
R12122 VSS.n174 VSS.n173 4.5005
R12123 VSS.n18622 VSS.n18621 4.5005
R12124 VSS.n186 VSS.n176 4.5005
R12125 VSS.n18651 VSS.n155 4.5005
R12126 VSS.n18682 VSS.n135 4.5005
R12127 VSS.n18596 VSS.n18595 4.5005
R12128 VSS.n143 VSS.n142 4.5005
R12129 VSS.n18671 VSS.n143 4.5005
R12130 VSS.n172 VSS.n170 4.5005
R12131 VSS.n170 VSS.n169 4.5005
R12132 VSS.n18611 VSS.n185 4.5005
R12133 VSS.n18663 VSS.n18662 4.5005
R12134 VSS.n18663 VSS.n149 4.5005
R12135 VSS.n18718 VSS.n18717 4.5005
R12136 VSS.n18717 VSS.n18716 4.5005
R12137 VSS.n18841 VSS.n66 4.5005
R12138 VSS.n18782 VSS.n93 4.5005
R12139 VSS.n18745 VSS.n18744 4.5005
R12140 VSS.n18695 VSS.n18693 4.5005
R12141 VSS.n18724 VSS.n18723 4.5005
R12142 VSS.n18735 VSS.n18734 4.5005
R12143 VSS.n18736 VSS.n18735 4.5005
R12144 VSS.n18769 VSS.n18768 4.5005
R12145 VSS.n18742 VSS.n18741 4.5005
R12146 VSS.n102 VSS.n101 4.5005
R12147 VSS.n111 VSS.n102 4.5005
R12148 VSS.n18836 VSS.n18835 4.5005
R12149 VSS.n18809 VSS.n82 4.5005
R12150 VSS.n18809 VSS.n76 4.5005
R12151 VSS.n18816 VSS.n78 4.5005
R12152 VSS.n18787 VSS.n18783 4.5005
R12153 VSS.n18787 VSS.n18786 4.5005
R12154 VSS.n18790 VSS.n18781 4.5005
R12155 VSS.n18774 VSS.n18773 4.5005
R12156 VSS.n18773 VSS.n88 4.5005
R12157 VSS.n18840 VSS.n18839 4.5005
R12158 VSS.n67 VSS.n65 4.5005
R12159 VSS.n65 VSS.n64 4.5005
R12160 VSS.n18797 VSS.n18796 4.5005
R12161 VSS.n18798 VSS.n18797 4.5005
R12162 VSS.n79 VSS.n77 4.5005
R12163 VSS.n18855 VSS.n18854 4.5005
R12164 VSS.n18726 VSS.n18725 4.5005
R12165 VSS.n18727 VSS.n122 4.5005
R12166 VSS.n408 VSS.n407 4.5005
R12167 VSS.n410 VSS.n409 4.5005
R12168 VSS.n391 VSS.n390 4.5005
R12169 VSS.n367 VSS.n299 4.5005
R12170 VSS.n351 VSS.n345 4.5005
R12171 VSS.n354 VSS.n353 4.5005
R12172 VSS.n350 VSS.n349 4.5005
R12173 VSS.n321 VSS.n319 4.5005
R12174 VSS.n420 VSS.n419 4.5005
R12175 VSS.n427 VSS.n311 4.5005
R12176 VSS.n434 VSS.n433 4.5005
R12177 VSS.n435 VSS.n302 4.5005
R12178 VSS.n442 VSS.n441 4.5005
R12179 VSS.n426 VSS.n425 4.5005
R12180 VSS.n411 VSS.n324 4.5005
R12181 VSS.n450 VSS.n449 4.5005
R12182 VSS.n327 VSS.n326 4.5005
R12183 VSS.n328 VSS.n327 4.5005
R12184 VSS.n378 VSS.n307 4.5005
R12185 VSS.n369 VSS.n368 4.5005
R12186 VSS.n369 VSS.n342 4.5005
R12187 VSS.n352 VSS.n346 4.5005
R12188 VSS.n389 VSS.n388 4.5005
R12189 VSS.n388 VSS.n332 4.5005
R12190 VSS.n18592 VSS.n18591 4.5005
R12191 VSS.n18591 VSS.n18590 4.5005
R12192 VSS.n619 VSS.n618 4.5005
R12193 VSS.n622 VSS.n621 4.5005
R12194 VSS.n605 VSS.n604 4.5005
R12195 VSS.n580 VSS.n579 4.5005
R12196 VSS.n571 VSS.n570 4.5005
R12197 VSS.n572 VSS.n566 4.5005
R12198 VSS.n568 VSS.n567 4.5005
R12199 VSS.n526 VSS.n524 4.5005
R12200 VSS.n848 VSS.n847 4.5005
R12201 VSS.n855 VSS.n516 4.5005
R12202 VSS.n862 VSS.n861 4.5005
R12203 VSS.n863 VSS.n508 4.5005
R12204 VSS.n576 VSS.n505 4.5005
R12205 VSS.n870 VSS.n869 4.5005
R12206 VSS.n854 VSS.n853 4.5005
R12207 VSS.n620 VSS.n541 4.5005
R12208 VSS.n878 VSS.n877 4.5005
R12209 VSS.n617 VSS.n542 4.5005
R12210 VSS.n617 VSS.n616 4.5005
R12211 VSS.n578 VSS.n577 4.5005
R12212 VSS.n577 VSS.n552 4.5005
R12213 VSS.n574 VSS.n573 4.5005
R12214 VSS.n607 VSS.n606 4.5005
R12215 VSS.n607 VSS.n600 4.5005
R12216 VSS.n840 VSS.n534 4.5005
R12217 VSS.n840 VSS.n839 4.5005
R12218 VSS.n732 VSS.n49 4.5005
R12219 VSS.n739 VSS.n738 4.5005
R12220 VSS.n784 VSS.n713 4.5005
R12221 VSS.n805 VSS.n668 4.5005
R12222 VSS.n668 VSS.n666 4.5005
R12223 VSS.n655 VSS.n654 4.5005
R12224 VSS.n647 VSS.n631 4.5005
R12225 VSS.n673 VSS.n672 4.5005
R12226 VSS.n656 VSS.n644 4.5005
R12227 VSS.n821 VSS.n639 4.5005
R12228 VSS.n639 VSS.n637 4.5005
R12229 VSS.n702 VSS.n701 4.5005
R12230 VSS.n707 VSS.n706 4.5005
R12231 VSS.n706 VSS.n684 4.5005
R12232 VSS.n791 VSS.n790 4.5005
R12233 VSS.n792 VSS.n791 4.5005
R12234 VSS.n751 VSS.n750 4.5005
R12235 VSS.n751 VSS.n746 4.5005
R12236 VSS.n779 VSS.n778 4.5005
R12237 VSS.n780 VSS.n779 4.5005
R12238 VSS.n774 VSS.n720 4.5005
R12239 VSS.n766 VSS.n729 4.5005
R12240 VSS.n766 VSS.n765 4.5005
R12241 VSS.n50 VSS.n43 4.5005
R12242 VSS.n777 VSS.n718 4.5005
R12243 VSS.n640 VSS.n638 4.5005
R12244 VSS.n740 VSS.n731 4.5005
R12245 VSS.n749 VSS.n689 4.5005
R12246 VSS.n807 VSS.n806 4.5005
R12247 VSS.n963 VSS.n962 4.5005
R12248 VSS.n966 VSS.n965 4.5005
R12249 VSS.n948 VSS.n947 4.5005
R12250 VSS.n923 VSS.n465 4.5005
R12251 VSS.n916 VSS.n915 4.5005
R12252 VSS.n917 VSS.n909 4.5005
R12253 VSS.n913 VSS.n910 4.5005
R12254 VSS.n487 VSS.n485 4.5005
R12255 VSS.n985 VSS.n984 4.5005
R12256 VSS.n992 VSS.n477 4.5005
R12257 VSS.n999 VSS.n998 4.5005
R12258 VSS.n1000 VSS.n468 4.5005
R12259 VSS.n1007 VSS.n1006 4.5005
R12260 VSS.n991 VSS.n990 4.5005
R12261 VSS.n964 VSS.n888 4.5005
R12262 VSS.n1015 VSS.n1014 4.5005
R12263 VSS.n961 VSS.n889 4.5005
R12264 VSS.n961 VSS.n960 4.5005
R12265 VSS.n895 VSS.n473 4.5005
R12266 VSS.n922 VSS.n921 4.5005
R12267 VSS.n922 VSS.n900 4.5005
R12268 VSS.n919 VSS.n918 4.5005
R12269 VSS.n950 VSS.n949 4.5005
R12270 VSS.n950 VSS.n943 4.5005
R12271 VSS.n977 VSS.n881 4.5005
R12272 VSS.n977 VSS.n976 4.5005
R12273 VSS.n1429 VSS.n1428 4.5005
R12274 VSS.n1399 VSS.n1348 4.5005
R12275 VSS.n17921 VSS.n17920 4.5005
R12276 VSS.n1306 VSS.n1290 4.5005
R12277 VSS.n1314 VSS.n1313 4.5005
R12278 VSS.n17935 VSS.n1298 4.5005
R12279 VSS.n1298 VSS.n1296 4.5005
R12280 VSS.n1361 VSS.n1360 4.5005
R12281 VSS.n1332 VSS.n1331 4.5005
R12282 VSS.n17919 VSS.n1327 4.5005
R12283 VSS.n1327 VSS.n1325 4.5005
R12284 VSS.n1434 VSS.n1418 4.5005
R12285 VSS.n17893 VSS.n17892 4.5005
R12286 VSS.n17894 VSS.n17893 4.5005
R12287 VSS.n17888 VSS.n1379 4.5005
R12288 VSS.n1401 VSS.n1400 4.5005
R12289 VSS.n1401 VSS.n1396 4.5005
R12290 VSS.n17898 VSS.n1372 4.5005
R12291 VSS.n1366 VSS.n1365 4.5005
R12292 VSS.n1365 VSS.n1343 4.5005
R12293 VSS.n1430 VSS.n1426 4.5005
R12294 VSS.n17880 VSS.n1388 4.5005
R12295 VSS.n17880 VSS.n17879 4.5005
R12296 VSS.n17905 VSS.n17904 4.5005
R12297 VSS.n17906 VSS.n17905 4.5005
R12298 VSS.n17891 VSS.n1377 4.5005
R12299 VSS.n1419 VSS.n1417 4.5005
R12300 VSS.n1299 VSS.n1297 4.5005
R12301 VSS.n1315 VSS.n1303 4.5005
R12302 VSS.n17129 VSS.n16935 3.69976
R12303 VSS.n17721 VSS.n17349 3.69976
R12304 VSS.n9771 VSS.n9399 3.69976
R12305 VSS.n16714 VSS.n16341 3.69976
R12306 VSS.n16121 VSS.n1513 3.69976
R12307 VSS.n2306 VSS.n1977 3.69976
R12308 VSS.n3262 VSS.n2890 3.69976
R12309 VSS.n3854 VSS.n3482 3.69976
R12310 VSS.n4446 VSS.n4074 3.69976
R12311 VSS.n5038 VSS.n4666 3.69976
R12312 VSS.n5271 VSS.n2573 3.69976
R12313 VSS.n5844 VSS.n5534 3.69976
R12314 VSS.n6436 VSS.n6107 3.69976
R12315 VSS.n7995 VSS.n7623 3.69976
R12316 VSS.n8587 VSS.n8215 3.69976
R12317 VSS.n9179 VSS.n8807 3.69976
R12318 VSS.n10363 VSS.n9991 3.69976
R12319 VSS.n10955 VSS.n10583 3.69976
R12320 VSS.n11547 VSS.n11175 3.69976
R12321 VSS.n12139 VSS.n11767 3.69976
R12322 VSS.n12731 VSS.n12359 3.69976
R12323 VSS.n13323 VSS.n12951 3.69976
R12324 VSS.n13915 VSS.n13543 3.69976
R12325 VSS.n14507 VSS.n14135 3.69976
R12326 VSS.n15099 VSS.n14727 3.69976
R12327 VSS.n15691 VSS.n15319 3.69976
R12328 VSS.n15924 VSS.n6713 3.69976
R12329 VSS.n7403 VSS.n7030 3.69976
R12330 VSS.n18715 VSS.n128 3.69976
R12331 VSS.n18541 VSS.n18212 3.69976
R12332 VSS.n838 VSS.n533 3.69976
R12333 VSS.n17952 VSS.n1195 3.69976
R12334 VSS.n18172 VSS.n216 3.69922
R12335 VSS.n9645 VSS.n9474 3.69922
R12336 VSS.n16588 VSS.n16416 3.69922
R12337 VSS.n15995 VSS.n1581 3.69922
R12338 VSS.n1937 VSS.n1766 3.69922
R12339 VSS.n3136 VSS.n2965 3.69922
R12340 VSS.n3728 VSS.n3557 3.69922
R12341 VSS.n4320 VSS.n4149 3.69922
R12342 VSS.n4912 VSS.n4741 3.69922
R12343 VSS.n2533 VSS.n2362 3.69922
R12344 VSS.n5494 VSS.n5323 3.69922
R12345 VSS.n6067 VSS.n5896 3.69922
R12346 VSS.n7869 VSS.n7698 3.69922
R12347 VSS.n8461 VSS.n8290 3.69922
R12348 VSS.n9053 VSS.n8882 3.69922
R12349 VSS.n10237 VSS.n10066 3.69922
R12350 VSS.n10829 VSS.n10658 3.69922
R12351 VSS.n11421 VSS.n11250 3.69922
R12352 VSS.n12013 VSS.n11842 3.69922
R12353 VSS.n12605 VSS.n12434 3.69922
R12354 VSS.n13197 VSS.n13026 3.69922
R12355 VSS.n13789 VSS.n13618 3.69922
R12356 VSS.n14381 VSS.n14210 3.69922
R12357 VSS.n14973 VSS.n14802 3.69922
R12358 VSS.n15565 VSS.n15394 3.69922
R12359 VSS.n6673 VSS.n6502 3.69922
R12360 VSS.n7277 VSS.n7105 3.69922
R12361 VSS.n18589 VSS.n196 3.69922
R12362 VSS.n975 VSS.n494 3.69922
R12363 VSS.n18001 VSS.n1061 3.69922
R12364 VSS.n17595 VSS.n17424 3.69922
R12365 VSS.n17991 VSS.n1160 3.42389
R12366 VSS.n17007 VSS.n1062 3.42389
R12367 VSS.n17009 VSS.n17008 3.42389
R12368 VSS.n17599 VSS.n17598 3.42389
R12369 VSS.n17601 VSS.n17600 3.42389
R12370 VSS.n18580 VSS.n18177 3.42389
R12371 VSS.n18176 VSS.n18175 3.42389
R12372 VSS.n9651 VSS.n9650 3.42389
R12373 VSS.n9649 VSS.n9648 3.42389
R12374 VSS.n16594 VSS.n16593 3.42389
R12375 VSS.n16592 VSS.n16591 3.42389
R12376 VSS.n16001 VSS.n16000 3.42389
R12377 VSS.n15999 VSS.n15998 3.42389
R12378 VSS.n2345 VSS.n1942 3.42389
R12379 VSS.n1941 VSS.n1940 3.42389
R12380 VSS.n3142 VSS.n3141 3.42389
R12381 VSS.n3140 VSS.n3139 3.42389
R12382 VSS.n3734 VSS.n3733 3.42389
R12383 VSS.n3732 VSS.n3731 3.42389
R12384 VSS.n4326 VSS.n4325 3.42389
R12385 VSS.n4324 VSS.n4323 3.42389
R12386 VSS.n4918 VSS.n4917 3.42389
R12387 VSS.n4916 VSS.n4915 3.42389
R12388 VSS.n5310 VSS.n2538 3.42389
R12389 VSS.n2537 VSS.n2536 3.42389
R12390 VSS.n5883 VSS.n5499 3.42389
R12391 VSS.n5498 VSS.n5497 3.42389
R12392 VSS.n6475 VSS.n6072 3.42389
R12393 VSS.n6071 VSS.n6070 3.42389
R12394 VSS.n7875 VSS.n7874 3.42389
R12395 VSS.n7873 VSS.n7872 3.42389
R12396 VSS.n8467 VSS.n8466 3.42389
R12397 VSS.n8465 VSS.n8464 3.42389
R12398 VSS.n9059 VSS.n9058 3.42389
R12399 VSS.n9057 VSS.n9056 3.42389
R12400 VSS.n10243 VSS.n10242 3.42389
R12401 VSS.n10241 VSS.n10240 3.42389
R12402 VSS.n10835 VSS.n10834 3.42389
R12403 VSS.n10833 VSS.n10832 3.42389
R12404 VSS.n11427 VSS.n11426 3.42389
R12405 VSS.n11425 VSS.n11424 3.42389
R12406 VSS.n12019 VSS.n12018 3.42389
R12407 VSS.n12017 VSS.n12016 3.42389
R12408 VSS.n12611 VSS.n12610 3.42389
R12409 VSS.n12609 VSS.n12608 3.42389
R12410 VSS.n13203 VSS.n13202 3.42389
R12411 VSS.n13201 VSS.n13200 3.42389
R12412 VSS.n13795 VSS.n13794 3.42389
R12413 VSS.n13793 VSS.n13792 3.42389
R12414 VSS.n14387 VSS.n14386 3.42389
R12415 VSS.n14385 VSS.n14384 3.42389
R12416 VSS.n14979 VSS.n14978 3.42389
R12417 VSS.n14977 VSS.n14976 3.42389
R12418 VSS.n15571 VSS.n15570 3.42389
R12419 VSS.n15569 VSS.n15568 3.42389
R12420 VSS.n15963 VSS.n6678 3.42389
R12421 VSS.n6677 VSS.n6676 3.42389
R12422 VSS.n7283 VSS.n7282 3.42389
R12423 VSS.n7281 VSS.n7280 3.42389
R12424 VSS.n18595 VSS.n18594 3.42389
R12425 VSS.n18593 VSS.n18592 3.42389
R12426 VSS.n879 VSS.n878 3.42389
R12427 VSS.n881 VSS.n880 3.42389
R12428 VSS.n1309 VSS.n1196 3.423
R12429 VSS.n18040 VSS.n1025 3.423
R12430 VSS.n17133 VSS.n17132 3.423
R12431 VSS.n17503 VSS.n17502 3.423
R12432 VSS.n17725 VSS.n17724 3.423
R12433 VSS.n18327 VSS.n18213 3.423
R12434 VSS.n18080 VSS.n18079 3.423
R12435 VSS.n9775 VSS.n9774 3.423
R12436 VSS.n9553 VSS.n9552 3.423
R12437 VSS.n16718 VSS.n16717 3.423
R12438 VSS.n16489 VSS.n16488 3.423
R12439 VSS.n16125 VSS.n16124 3.423
R12440 VSS.n1654 VSS.n1653 3.423
R12441 VSS.n2091 VSS.n1978 3.423
R12442 VSS.n1845 VSS.n1844 3.423
R12443 VSS.n3266 VSS.n3265 3.423
R12444 VSS.n3044 VSS.n3043 3.423
R12445 VSS.n3858 VSS.n3857 3.423
R12446 VSS.n3636 VSS.n3635 3.423
R12447 VSS.n4450 VSS.n4449 3.423
R12448 VSS.n4228 VSS.n4227 3.423
R12449 VSS.n5042 VSS.n5041 3.423
R12450 VSS.n4820 VSS.n4819 3.423
R12451 VSS.n2687 VSS.n2574 3.423
R12452 VSS.n2441 VSS.n2440 3.423
R12453 VSS.n5648 VSS.n5535 3.423
R12454 VSS.n5402 VSS.n5401 3.423
R12455 VSS.n6221 VSS.n6108 3.423
R12456 VSS.n5975 VSS.n5974 3.423
R12457 VSS.n7999 VSS.n7998 3.423
R12458 VSS.n7777 VSS.n7776 3.423
R12459 VSS.n8591 VSS.n8590 3.423
R12460 VSS.n8369 VSS.n8368 3.423
R12461 VSS.n9183 VSS.n9182 3.423
R12462 VSS.n8961 VSS.n8960 3.423
R12463 VSS.n10367 VSS.n10366 3.423
R12464 VSS.n10145 VSS.n10144 3.423
R12465 VSS.n10959 VSS.n10958 3.423
R12466 VSS.n10737 VSS.n10736 3.423
R12467 VSS.n11551 VSS.n11550 3.423
R12468 VSS.n11329 VSS.n11328 3.423
R12469 VSS.n12143 VSS.n12142 3.423
R12470 VSS.n11921 VSS.n11920 3.423
R12471 VSS.n12735 VSS.n12734 3.423
R12472 VSS.n12513 VSS.n12512 3.423
R12473 VSS.n13327 VSS.n13326 3.423
R12474 VSS.n13105 VSS.n13104 3.423
R12475 VSS.n13919 VSS.n13918 3.423
R12476 VSS.n13697 VSS.n13696 3.423
R12477 VSS.n14511 VSS.n14510 3.423
R12478 VSS.n14289 VSS.n14288 3.423
R12479 VSS.n15103 VSS.n15102 3.423
R12480 VSS.n14881 VSS.n14880 3.423
R12481 VSS.n15695 VSS.n15694 3.423
R12482 VSS.n15473 VSS.n15472 3.423
R12483 VSS.n6827 VSS.n6714 3.423
R12484 VSS.n6581 VSS.n6580 3.423
R12485 VSS.n7407 VSS.n7406 3.423
R12486 VSS.n7178 VSS.n7177 3.423
R12487 VSS.n18719 VSS.n18718 3.423
R12488 VSS.n449 VSS.n292 3.423
R12489 VSS.n650 VSS.n534 3.423
R12490 VSS.n1014 VSS.n458 3.423
R12491 VSS.n17252 VSS.n17247 3.4105
R12492 VSS.n17252 VSS.n17251 3.4105
R12493 VSS.n17246 VSS.n16874 3.4105
R12494 VSS.n17271 VSS.n17270 3.4105
R12495 VSS.n17270 VSS.n17269 3.4105
R12496 VSS.n17229 VSS.n17227 3.4105
R12497 VSS.n17229 VSS.n17228 3.4105
R12498 VSS.n17245 VSS.n17244 3.4105
R12499 VSS.n17244 VSS.n17243 3.4105
R12500 VSS.n17207 VSS.n17206 3.4105
R12501 VSS.n17206 VSS.n17205 3.4105
R12502 VSS.n16888 VSS.n16887 3.4105
R12503 VSS.n17226 VSS.n17225 3.4105
R12504 VSS.n17225 VSS.n17224 3.4105
R12505 VSS.n17190 VSS.n17189 3.4105
R12506 VSS.n17209 VSS.n17208 3.4105
R12507 VSS.n17174 VSS.n17173 3.4105
R12508 VSS.n17173 VSS.n17172 3.4105
R12509 VSS.n17175 VSS.n16906 3.4105
R12510 VSS.n17178 VSS.n16901 3.4105
R12511 VSS.n17147 VSS.n17146 3.4105
R12512 VSS.n17147 VSS.n16924 3.4105
R12513 VSS.n16920 VSS.n16907 3.4105
R12514 VSS.n17154 VSS.n16920 3.4105
R12515 VSS.n18006 VSS.n18005 3.4105
R12516 VSS.n18005 VSS.n18004 3.4105
R12517 VSS.n18013 VSS.n18012 3.4105
R12518 VSS.n18008 VSS.n18007 3.4105
R12519 VSS.n18009 VSS.n18008 3.4105
R12520 VSS.n18021 VSS.n18020 3.4105
R12521 VSS.n18020 VSS.n18019 3.4105
R12522 VSS.n1047 VSS.n1042 3.4105
R12523 VSS.n18015 VSS.n18014 3.4105
R12524 VSS.n18015 VSS.n1046 3.4105
R12525 VSS.n18029 VSS.n18028 3.4105
R12526 VSS.n18028 VSS.n18027 3.4105
R12527 VSS.n1041 VSS.n1039 3.4105
R12528 VSS.n18023 VSS.n18022 3.4105
R12529 VSS.n18023 VSS.n1037 3.4105
R12530 VSS.n18036 VSS.n18035 3.4105
R12531 VSS.n18035 VSS.n18034 3.4105
R12532 VSS.n18031 VSS.n18030 3.4105
R12533 VSS.n18037 VSS.n1026 3.4105
R12534 VSS.n1026 VSS.n1024 3.4105
R12535 VSS.n17134 VSS.n16931 3.4105
R12536 VSS.n17108 VSS.n16931 3.4105
R12537 VSS.n16928 VSS.n16927 3.4105
R12538 VSS.n17144 VSS.n17143 3.4105
R12539 VSS.n17143 VSS.n17142 3.4105
R12540 VSS.n17093 VSS.n17092 3.4105
R12541 VSS.n17093 VSS.n16934 3.4105
R12542 VSS.n17070 VSS.n17069 3.4105
R12543 VSS.n17091 VSS.n17090 3.4105
R12544 VSS.n17090 VSS.n17089 3.4105
R12545 VSS.n17060 VSS.n16964 3.4105
R12546 VSS.n16964 VSS.n16963 3.4105
R12547 VSS.n17062 VSS.n17061 3.4105
R12548 VSS.n17068 VSS.n17067 3.4105
R12549 VSS.n17067 VSS.n17066 3.4105
R12550 VSS.n17043 VSS.n17042 3.4105
R12551 VSS.n17043 VSS.n16978 3.4105
R12552 VSS.n17039 VSS.n16966 3.4105
R12553 VSS.n17059 VSS.n17058 3.4105
R12554 VSS.n17058 VSS.n17057 3.4105
R12555 VSS.n17022 VSS.n17021 3.4105
R12556 VSS.n17022 VSS.n16994 3.4105
R12557 VSS.n17038 VSS.n17037 3.4105
R12558 VSS.n17020 VSS.n17019 3.4105
R12559 VSS.n17019 VSS.n17018 3.4105
R12560 VSS.n17844 VSS.n17839 3.4105
R12561 VSS.n17844 VSS.n17843 3.4105
R12562 VSS.n17838 VSS.n17288 3.4105
R12563 VSS.n17863 VSS.n17862 3.4105
R12564 VSS.n17862 VSS.n17861 3.4105
R12565 VSS.n17821 VSS.n17819 3.4105
R12566 VSS.n17821 VSS.n17820 3.4105
R12567 VSS.n17837 VSS.n17836 3.4105
R12568 VSS.n17836 VSS.n17835 3.4105
R12569 VSS.n17799 VSS.n17798 3.4105
R12570 VSS.n17798 VSS.n17797 3.4105
R12571 VSS.n17302 VSS.n17301 3.4105
R12572 VSS.n17818 VSS.n17817 3.4105
R12573 VSS.n17817 VSS.n17816 3.4105
R12574 VSS.n17782 VSS.n17781 3.4105
R12575 VSS.n17801 VSS.n17800 3.4105
R12576 VSS.n17766 VSS.n17765 3.4105
R12577 VSS.n17765 VSS.n17764 3.4105
R12578 VSS.n17767 VSS.n17320 3.4105
R12579 VSS.n17770 VSS.n17315 3.4105
R12580 VSS.n17739 VSS.n17738 3.4105
R12581 VSS.n17739 VSS.n17338 3.4105
R12582 VSS.n17334 VSS.n17321 3.4105
R12583 VSS.n17746 VSS.n17334 3.4105
R12584 VSS.n17578 VSS.n17577 3.4105
R12585 VSS.n17578 VSS.n17423 3.4105
R12586 VSS.n17571 VSS.n17570 3.4105
R12587 VSS.n17576 VSS.n17575 3.4105
R12588 VSS.n17575 VSS.n17574 3.4105
R12589 VSS.n17551 VSS.n17550 3.4105
R12590 VSS.n17551 VSS.n17463 3.4105
R12591 VSS.n17549 VSS.n17548 3.4105
R12592 VSS.n17569 VSS.n17568 3.4105
R12593 VSS.n17568 VSS.n17567 3.4105
R12594 VSS.n17538 VSS.n17469 3.4105
R12595 VSS.n17469 VSS.n17468 3.4105
R12596 VSS.n17467 VSS.n17466 3.4105
R12597 VSS.n17546 VSS.n17545 3.4105
R12598 VSS.n17545 VSS.n17461 3.4105
R12599 VSS.n17516 VSS.n17515 3.4105
R12600 VSS.n17516 VSS.n17488 3.4105
R12601 VSS.n17537 VSS.n17536 3.4105
R12602 VSS.n17514 VSS.n17513 3.4105
R12603 VSS.n17513 VSS.n17512 3.4105
R12604 VSS.n17726 VSS.n17345 3.4105
R12605 VSS.n17700 VSS.n17345 3.4105
R12606 VSS.n17342 VSS.n17341 3.4105
R12607 VSS.n17736 VSS.n17735 3.4105
R12608 VSS.n17735 VSS.n17734 3.4105
R12609 VSS.n17685 VSS.n17684 3.4105
R12610 VSS.n17685 VSS.n17348 3.4105
R12611 VSS.n17662 VSS.n17661 3.4105
R12612 VSS.n17683 VSS.n17682 3.4105
R12613 VSS.n17682 VSS.n17681 3.4105
R12614 VSS.n17652 VSS.n17378 3.4105
R12615 VSS.n17378 VSS.n17377 3.4105
R12616 VSS.n17654 VSS.n17653 3.4105
R12617 VSS.n17660 VSS.n17659 3.4105
R12618 VSS.n17659 VSS.n17658 3.4105
R12619 VSS.n17635 VSS.n17634 3.4105
R12620 VSS.n17635 VSS.n17392 3.4105
R12621 VSS.n17631 VSS.n17380 3.4105
R12622 VSS.n17651 VSS.n17650 3.4105
R12623 VSS.n17650 VSS.n17649 3.4105
R12624 VSS.n17614 VSS.n17613 3.4105
R12625 VSS.n17614 VSS.n17408 3.4105
R12626 VSS.n17630 VSS.n17629 3.4105
R12627 VSS.n17612 VSS.n17611 3.4105
R12628 VSS.n17611 VSS.n17610 3.4105
R12629 VSS.n18471 VSS.n18470 3.4105
R12630 VSS.n18472 VSS.n18471 3.4105
R12631 VSS.n18469 VSS.n18427 3.4105
R12632 VSS.n18466 VSS.n18430 3.4105
R12633 VSS.n18466 VSS.n18465 3.4105
R12634 VSS.n18485 VSS.n18484 3.4105
R12635 VSS.n18484 VSS.n18483 3.4105
R12636 VSS.n18428 VSS.n18424 3.4105
R12637 VSS.n18424 VSS.n18422 3.4105
R12638 VSS.n18410 VSS.n18392 3.4105
R12639 VSS.n18410 VSS.n18409 3.4105
R12640 VSS.n18414 VSS.n18390 3.4105
R12641 VSS.n18487 VSS.n18486 3.4105
R12642 VSS.n18488 VSS.n18487 3.4105
R12643 VSS.n18503 VSS.n18502 3.4105
R12644 VSS.n18399 VSS.n18398 3.4105
R12645 VSS.n18348 VSS.n18337 3.4105
R12646 VSS.n18348 VSS.n18342 3.4105
R12647 VSS.n18350 VSS.n18349 3.4105
R12648 VSS.n18505 VSS.n18504 3.4105
R12649 VSS.n18523 VSS.n18522 3.4105
R12650 VSS.n18523 VSS.n18316 3.4105
R12651 VSS.n18520 VSS.n18519 3.4105
R12652 VSS.n18519 VSS.n18518 3.4105
R12653 VSS.n18546 VSS.n18545 3.4105
R12654 VSS.n18545 VSS.n18544 3.4105
R12655 VSS.n18553 VSS.n18552 3.4105
R12656 VSS.n18548 VSS.n18547 3.4105
R12657 VSS.n18549 VSS.n18548 3.4105
R12658 VSS.n18561 VSS.n18560 3.4105
R12659 VSS.n18560 VSS.n18559 3.4105
R12660 VSS.n18198 VSS.n18194 3.4105
R12661 VSS.n18555 VSS.n18554 3.4105
R12662 VSS.n18555 VSS.n18197 3.4105
R12663 VSS.n18569 VSS.n18568 3.4105
R12664 VSS.n18568 VSS.n18567 3.4105
R12665 VSS.n18193 VSS.n18191 3.4105
R12666 VSS.n18563 VSS.n18562 3.4105
R12667 VSS.n18563 VSS.n18189 3.4105
R12668 VSS.n18576 VSS.n18575 3.4105
R12669 VSS.n18575 VSS.n18574 3.4105
R12670 VSS.n18571 VSS.n18570 3.4105
R12671 VSS.n18577 VSS.n18178 3.4105
R12672 VSS.n18178 VSS.n212 3.4105
R12673 VSS.n18328 VSS.n18326 3.4105
R12674 VSS.n18326 VSS.n18325 3.4105
R12675 VSS.n18319 VSS.n18318 3.4105
R12676 VSS.n18336 VSS.n18335 3.4105
R12677 VSS.n18335 VSS.n18334 3.4105
R12678 VSS.n18155 VSS.n18154 3.4105
R12679 VSS.n18155 VSS.n215 3.4105
R12680 VSS.n18148 VSS.n18147 3.4105
R12681 VSS.n18153 VSS.n18152 3.4105
R12682 VSS.n18152 VSS.n18151 3.4105
R12683 VSS.n18128 VSS.n18127 3.4105
R12684 VSS.n18128 VSS.n255 3.4105
R12685 VSS.n18126 VSS.n18125 3.4105
R12686 VSS.n18146 VSS.n18145 3.4105
R12687 VSS.n18145 VSS.n18144 3.4105
R12688 VSS.n18115 VSS.n261 3.4105
R12689 VSS.n261 VSS.n260 3.4105
R12690 VSS.n259 VSS.n258 3.4105
R12691 VSS.n18123 VSS.n18122 3.4105
R12692 VSS.n18122 VSS.n253 3.4105
R12693 VSS.n18093 VSS.n18092 3.4105
R12694 VSS.n18093 VSS.n280 3.4105
R12695 VSS.n18114 VSS.n18113 3.4105
R12696 VSS.n18091 VSS.n18090 3.4105
R12697 VSS.n18090 VSS.n18089 3.4105
R12698 VSS.n9888 VSS.n9339 3.4105
R12699 VSS.n9894 VSS.n9339 3.4105
R12700 VSS.n9890 VSS.n9889 3.4105
R12701 VSS.n9914 VSS.n9913 3.4105
R12702 VSS.n9913 VSS.n9912 3.4105
R12703 VSS.n9871 VSS.n9869 3.4105
R12704 VSS.n9871 VSS.n9870 3.4105
R12705 VSS.n9887 VSS.n9886 3.4105
R12706 VSS.n9886 VSS.n9885 3.4105
R12707 VSS.n9849 VSS.n9848 3.4105
R12708 VSS.n9848 VSS.n9847 3.4105
R12709 VSS.n9352 VSS.n9351 3.4105
R12710 VSS.n9868 VSS.n9867 3.4105
R12711 VSS.n9867 VSS.n9866 3.4105
R12712 VSS.n9832 VSS.n9831 3.4105
R12713 VSS.n9851 VSS.n9850 3.4105
R12714 VSS.n9816 VSS.n9815 3.4105
R12715 VSS.n9815 VSS.n9814 3.4105
R12716 VSS.n9817 VSS.n9370 3.4105
R12717 VSS.n9820 VSS.n9365 3.4105
R12718 VSS.n9789 VSS.n9788 3.4105
R12719 VSS.n9789 VSS.n9388 3.4105
R12720 VSS.n9384 VSS.n9371 3.4105
R12721 VSS.n9796 VSS.n9384 3.4105
R12722 VSS.n9735 VSS.n9734 3.4105
R12723 VSS.n9735 VSS.n9398 3.4105
R12724 VSS.n9712 VSS.n9711 3.4105
R12725 VSS.n9733 VSS.n9732 3.4105
R12726 VSS.n9732 VSS.n9731 3.4105
R12727 VSS.n9702 VSS.n9428 3.4105
R12728 VSS.n9428 VSS.n9427 3.4105
R12729 VSS.n9704 VSS.n9703 3.4105
R12730 VSS.n9710 VSS.n9709 3.4105
R12731 VSS.n9709 VSS.n9708 3.4105
R12732 VSS.n9685 VSS.n9684 3.4105
R12733 VSS.n9685 VSS.n9442 3.4105
R12734 VSS.n9681 VSS.n9430 3.4105
R12735 VSS.n9701 VSS.n9700 3.4105
R12736 VSS.n9700 VSS.n9699 3.4105
R12737 VSS.n9664 VSS.n9663 3.4105
R12738 VSS.n9664 VSS.n9458 3.4105
R12739 VSS.n9680 VSS.n9679 3.4105
R12740 VSS.n9662 VSS.n9661 3.4105
R12741 VSS.n9661 VSS.n9660 3.4105
R12742 VSS.n9776 VSS.n9395 3.4105
R12743 VSS.n9750 VSS.n9395 3.4105
R12744 VSS.n9392 VSS.n9391 3.4105
R12745 VSS.n9786 VSS.n9785 3.4105
R12746 VSS.n9785 VSS.n9784 3.4105
R12747 VSS.n9628 VSS.n9627 3.4105
R12748 VSS.n9628 VSS.n9473 3.4105
R12749 VSS.n9621 VSS.n9620 3.4105
R12750 VSS.n9626 VSS.n9625 3.4105
R12751 VSS.n9625 VSS.n9624 3.4105
R12752 VSS.n9601 VSS.n9600 3.4105
R12753 VSS.n9601 VSS.n9513 3.4105
R12754 VSS.n9599 VSS.n9598 3.4105
R12755 VSS.n9619 VSS.n9618 3.4105
R12756 VSS.n9618 VSS.n9617 3.4105
R12757 VSS.n9588 VSS.n9519 3.4105
R12758 VSS.n9519 VSS.n9518 3.4105
R12759 VSS.n9517 VSS.n9516 3.4105
R12760 VSS.n9596 VSS.n9595 3.4105
R12761 VSS.n9595 VSS.n9511 3.4105
R12762 VSS.n9566 VSS.n9565 3.4105
R12763 VSS.n9566 VSS.n9538 3.4105
R12764 VSS.n9587 VSS.n9586 3.4105
R12765 VSS.n9564 VSS.n9563 3.4105
R12766 VSS.n9563 VSS.n9562 3.4105
R12767 VSS.n16831 VSS.n16281 3.4105
R12768 VSS.n16837 VSS.n16281 3.4105
R12769 VSS.n16833 VSS.n16832 3.4105
R12770 VSS.n16857 VSS.n16856 3.4105
R12771 VSS.n16856 VSS.n16855 3.4105
R12772 VSS.n16814 VSS.n16812 3.4105
R12773 VSS.n16814 VSS.n16813 3.4105
R12774 VSS.n16830 VSS.n16829 3.4105
R12775 VSS.n16829 VSS.n16828 3.4105
R12776 VSS.n16792 VSS.n16791 3.4105
R12777 VSS.n16791 VSS.n16790 3.4105
R12778 VSS.n16294 VSS.n16293 3.4105
R12779 VSS.n16811 VSS.n16810 3.4105
R12780 VSS.n16810 VSS.n16809 3.4105
R12781 VSS.n16775 VSS.n16774 3.4105
R12782 VSS.n16794 VSS.n16793 3.4105
R12783 VSS.n16759 VSS.n16758 3.4105
R12784 VSS.n16758 VSS.n16757 3.4105
R12785 VSS.n16760 VSS.n16312 3.4105
R12786 VSS.n16763 VSS.n16307 3.4105
R12787 VSS.n16732 VSS.n16731 3.4105
R12788 VSS.n16732 VSS.n16330 3.4105
R12789 VSS.n16326 VSS.n16313 3.4105
R12790 VSS.n16739 VSS.n16326 3.4105
R12791 VSS.n16678 VSS.n16677 3.4105
R12792 VSS.n16678 VSS.n16340 3.4105
R12793 VSS.n16655 VSS.n16654 3.4105
R12794 VSS.n16676 VSS.n16675 3.4105
R12795 VSS.n16675 VSS.n16674 3.4105
R12796 VSS.n16645 VSS.n16370 3.4105
R12797 VSS.n16370 VSS.n16369 3.4105
R12798 VSS.n16647 VSS.n16646 3.4105
R12799 VSS.n16653 VSS.n16652 3.4105
R12800 VSS.n16652 VSS.n16651 3.4105
R12801 VSS.n16628 VSS.n16627 3.4105
R12802 VSS.n16628 VSS.n16384 3.4105
R12803 VSS.n16624 VSS.n16372 3.4105
R12804 VSS.n16644 VSS.n16643 3.4105
R12805 VSS.n16643 VSS.n16642 3.4105
R12806 VSS.n16607 VSS.n16606 3.4105
R12807 VSS.n16607 VSS.n16400 3.4105
R12808 VSS.n16623 VSS.n16622 3.4105
R12809 VSS.n16605 VSS.n16604 3.4105
R12810 VSS.n16604 VSS.n16603 3.4105
R12811 VSS.n16719 VSS.n16337 3.4105
R12812 VSS.n16693 VSS.n16337 3.4105
R12813 VSS.n16334 VSS.n16333 3.4105
R12814 VSS.n16729 VSS.n16728 3.4105
R12815 VSS.n16728 VSS.n16727 3.4105
R12816 VSS.n16574 VSS.n16573 3.4105
R12817 VSS.n16574 VSS.n16415 3.4105
R12818 VSS.n16550 VSS.n16549 3.4105
R12819 VSS.n16572 VSS.n16571 3.4105
R12820 VSS.n16571 VSS.n16570 3.4105
R12821 VSS.n16540 VSS.n16445 3.4105
R12822 VSS.n16445 VSS.n16444 3.4105
R12823 VSS.n16542 VSS.n16541 3.4105
R12824 VSS.n16548 VSS.n16547 3.4105
R12825 VSS.n16547 VSS.n16546 3.4105
R12826 VSS.n16523 VSS.n16522 3.4105
R12827 VSS.n16523 VSS.n16461 3.4105
R12828 VSS.n16519 VSS.n16447 3.4105
R12829 VSS.n16539 VSS.n16538 3.4105
R12830 VSS.n16538 VSS.n16537 3.4105
R12831 VSS.n16502 VSS.n16501 3.4105
R12832 VSS.n16502 VSS.n16475 3.4105
R12833 VSS.n16518 VSS.n16517 3.4105
R12834 VSS.n16500 VSS.n16499 3.4105
R12835 VSS.n16499 VSS.n16498 3.4105
R12836 VSS.n16238 VSS.n1453 3.4105
R12837 VSS.n16244 VSS.n1453 3.4105
R12838 VSS.n16240 VSS.n16239 3.4105
R12839 VSS.n16264 VSS.n16263 3.4105
R12840 VSS.n16263 VSS.n16262 3.4105
R12841 VSS.n16221 VSS.n16219 3.4105
R12842 VSS.n16221 VSS.n16220 3.4105
R12843 VSS.n16237 VSS.n16236 3.4105
R12844 VSS.n16236 VSS.n16235 3.4105
R12845 VSS.n16199 VSS.n16198 3.4105
R12846 VSS.n16198 VSS.n16197 3.4105
R12847 VSS.n1466 VSS.n1465 3.4105
R12848 VSS.n16218 VSS.n16217 3.4105
R12849 VSS.n16217 VSS.n16216 3.4105
R12850 VSS.n16182 VSS.n16181 3.4105
R12851 VSS.n16201 VSS.n16200 3.4105
R12852 VSS.n16166 VSS.n16165 3.4105
R12853 VSS.n16165 VSS.n16164 3.4105
R12854 VSS.n16167 VSS.n1484 3.4105
R12855 VSS.n16170 VSS.n1479 3.4105
R12856 VSS.n16139 VSS.n16138 3.4105
R12857 VSS.n16139 VSS.n1502 3.4105
R12858 VSS.n1498 VSS.n1485 3.4105
R12859 VSS.n16146 VSS.n1498 3.4105
R12860 VSS.n16085 VSS.n16084 3.4105
R12861 VSS.n16085 VSS.n1512 3.4105
R12862 VSS.n16062 VSS.n16061 3.4105
R12863 VSS.n16083 VSS.n16082 3.4105
R12864 VSS.n16082 VSS.n16081 3.4105
R12865 VSS.n16052 VSS.n1542 3.4105
R12866 VSS.n1542 VSS.n1541 3.4105
R12867 VSS.n16054 VSS.n16053 3.4105
R12868 VSS.n16060 VSS.n16059 3.4105
R12869 VSS.n16059 VSS.n16058 3.4105
R12870 VSS.n16035 VSS.n16034 3.4105
R12871 VSS.n16035 VSS.n1556 3.4105
R12872 VSS.n16031 VSS.n1544 3.4105
R12873 VSS.n16051 VSS.n16050 3.4105
R12874 VSS.n16050 VSS.n16049 3.4105
R12875 VSS.n16014 VSS.n16013 3.4105
R12876 VSS.n16014 VSS.n1572 3.4105
R12877 VSS.n16030 VSS.n16029 3.4105
R12878 VSS.n16012 VSS.n16011 3.4105
R12879 VSS.n16011 VSS.n16010 3.4105
R12880 VSS.n16126 VSS.n1509 3.4105
R12881 VSS.n16100 VSS.n1509 3.4105
R12882 VSS.n1506 VSS.n1505 3.4105
R12883 VSS.n16136 VSS.n16135 3.4105
R12884 VSS.n16135 VSS.n16134 3.4105
R12885 VSS.n1739 VSS.n1738 3.4105
R12886 VSS.n1739 VSS.n1580 3.4105
R12887 VSS.n1715 VSS.n1714 3.4105
R12888 VSS.n1737 VSS.n1736 3.4105
R12889 VSS.n1736 VSS.n1735 3.4105
R12890 VSS.n1705 VSS.n1610 3.4105
R12891 VSS.n1610 VSS.n1609 3.4105
R12892 VSS.n1707 VSS.n1706 3.4105
R12893 VSS.n1713 VSS.n1712 3.4105
R12894 VSS.n1712 VSS.n1711 3.4105
R12895 VSS.n1688 VSS.n1687 3.4105
R12896 VSS.n1688 VSS.n1626 3.4105
R12897 VSS.n1684 VSS.n1612 3.4105
R12898 VSS.n1704 VSS.n1703 3.4105
R12899 VSS.n1703 VSS.n1702 3.4105
R12900 VSS.n1667 VSS.n1666 3.4105
R12901 VSS.n1667 VSS.n1640 3.4105
R12902 VSS.n1683 VSS.n1682 3.4105
R12903 VSS.n1665 VSS.n1664 3.4105
R12904 VSS.n1664 VSS.n1663 3.4105
R12905 VSS.n2215 VSS.n2169 3.4105
R12906 VSS.n2215 VSS.n2214 3.4105
R12907 VSS.n2218 VSS.n2217 3.4105
R12908 VSS.n2222 VSS.n2221 3.4105
R12909 VSS.n2223 VSS.n2222 3.4105
R12910 VSS.n2240 VSS.n2239 3.4105
R12911 VSS.n2241 VSS.n2240 3.4105
R12912 VSS.n2237 VSS.n2236 3.4105
R12913 VSS.n2236 VSS.n2235 3.4105
R12914 VSS.n2255 VSS.n2254 3.4105
R12915 VSS.n2254 VSS.n2253 3.4105
R12916 VSS.n2167 VSS.n2166 3.4105
R12917 VSS.n2168 VSS.n2160 3.4105
R12918 VSS.n2160 VSS.n2156 3.4105
R12919 VSS.n2150 VSS.n2149 3.4105
R12920 VSS.n2257 VSS.n2256 3.4105
R12921 VSS.n2272 VSS.n2118 3.4105
R12922 VSS.n2272 VSS.n2271 3.4105
R12923 VSS.n2135 VSS.n2111 3.4105
R12924 VSS.n2138 VSS.n2131 3.4105
R12925 VSS.n2288 VSS.n2101 3.4105
R12926 VSS.n2288 VSS.n2287 3.4105
R12927 VSS.n2117 VSS.n2116 3.4105
R12928 VSS.n2116 VSS.n2115 3.4105
R12929 VSS.n2311 VSS.n2310 3.4105
R12930 VSS.n2310 VSS.n2309 3.4105
R12931 VSS.n2318 VSS.n2317 3.4105
R12932 VSS.n2313 VSS.n2312 3.4105
R12933 VSS.n2314 VSS.n2313 3.4105
R12934 VSS.n2326 VSS.n2325 3.4105
R12935 VSS.n2325 VSS.n2324 3.4105
R12936 VSS.n1963 VSS.n1959 3.4105
R12937 VSS.n2320 VSS.n2319 3.4105
R12938 VSS.n2320 VSS.n1962 3.4105
R12939 VSS.n2334 VSS.n2333 3.4105
R12940 VSS.n2333 VSS.n2332 3.4105
R12941 VSS.n1958 VSS.n1956 3.4105
R12942 VSS.n2328 VSS.n2327 3.4105
R12943 VSS.n2328 VSS.n1954 3.4105
R12944 VSS.n2341 VSS.n2340 3.4105
R12945 VSS.n2340 VSS.n2339 3.4105
R12946 VSS.n2336 VSS.n2335 3.4105
R12947 VSS.n2342 VSS.n1943 3.4105
R12948 VSS.n1943 VSS.n1762 3.4105
R12949 VSS.n2092 VSS.n2090 3.4105
R12950 VSS.n2090 VSS.n2089 3.4105
R12951 VSS.n2084 VSS.n2083 3.4105
R12952 VSS.n2100 VSS.n2099 3.4105
R12953 VSS.n2099 VSS.n2098 3.4105
R12954 VSS.n1920 VSS.n1919 3.4105
R12955 VSS.n1920 VSS.n1765 3.4105
R12956 VSS.n1913 VSS.n1912 3.4105
R12957 VSS.n1918 VSS.n1917 3.4105
R12958 VSS.n1917 VSS.n1916 3.4105
R12959 VSS.n1893 VSS.n1892 3.4105
R12960 VSS.n1893 VSS.n1805 3.4105
R12961 VSS.n1891 VSS.n1890 3.4105
R12962 VSS.n1911 VSS.n1910 3.4105
R12963 VSS.n1910 VSS.n1909 3.4105
R12964 VSS.n1880 VSS.n1811 3.4105
R12965 VSS.n1811 VSS.n1810 3.4105
R12966 VSS.n1809 VSS.n1808 3.4105
R12967 VSS.n1888 VSS.n1887 3.4105
R12968 VSS.n1887 VSS.n1803 3.4105
R12969 VSS.n1858 VSS.n1857 3.4105
R12970 VSS.n1858 VSS.n1830 3.4105
R12971 VSS.n1879 VSS.n1878 3.4105
R12972 VSS.n1856 VSS.n1855 3.4105
R12973 VSS.n1855 VSS.n1854 3.4105
R12974 VSS.n3379 VSS.n2830 3.4105
R12975 VSS.n3385 VSS.n2830 3.4105
R12976 VSS.n3381 VSS.n3380 3.4105
R12977 VSS.n3405 VSS.n3404 3.4105
R12978 VSS.n3404 VSS.n3403 3.4105
R12979 VSS.n3362 VSS.n3360 3.4105
R12980 VSS.n3362 VSS.n3361 3.4105
R12981 VSS.n3378 VSS.n3377 3.4105
R12982 VSS.n3377 VSS.n3376 3.4105
R12983 VSS.n3340 VSS.n3339 3.4105
R12984 VSS.n3339 VSS.n3338 3.4105
R12985 VSS.n2843 VSS.n2842 3.4105
R12986 VSS.n3359 VSS.n3358 3.4105
R12987 VSS.n3358 VSS.n3357 3.4105
R12988 VSS.n3323 VSS.n3322 3.4105
R12989 VSS.n3342 VSS.n3341 3.4105
R12990 VSS.n3307 VSS.n3306 3.4105
R12991 VSS.n3306 VSS.n3305 3.4105
R12992 VSS.n3308 VSS.n2861 3.4105
R12993 VSS.n3311 VSS.n2856 3.4105
R12994 VSS.n3280 VSS.n3279 3.4105
R12995 VSS.n3280 VSS.n2879 3.4105
R12996 VSS.n2875 VSS.n2862 3.4105
R12997 VSS.n3287 VSS.n2875 3.4105
R12998 VSS.n3226 VSS.n3225 3.4105
R12999 VSS.n3226 VSS.n2889 3.4105
R13000 VSS.n3203 VSS.n3202 3.4105
R13001 VSS.n3224 VSS.n3223 3.4105
R13002 VSS.n3223 VSS.n3222 3.4105
R13003 VSS.n3193 VSS.n2919 3.4105
R13004 VSS.n2919 VSS.n2918 3.4105
R13005 VSS.n3195 VSS.n3194 3.4105
R13006 VSS.n3201 VSS.n3200 3.4105
R13007 VSS.n3200 VSS.n3199 3.4105
R13008 VSS.n3176 VSS.n3175 3.4105
R13009 VSS.n3176 VSS.n2933 3.4105
R13010 VSS.n3172 VSS.n2921 3.4105
R13011 VSS.n3192 VSS.n3191 3.4105
R13012 VSS.n3191 VSS.n3190 3.4105
R13013 VSS.n3155 VSS.n3154 3.4105
R13014 VSS.n3155 VSS.n2949 3.4105
R13015 VSS.n3171 VSS.n3170 3.4105
R13016 VSS.n3153 VSS.n3152 3.4105
R13017 VSS.n3152 VSS.n3151 3.4105
R13018 VSS.n3267 VSS.n2886 3.4105
R13019 VSS.n3241 VSS.n2886 3.4105
R13020 VSS.n2883 VSS.n2882 3.4105
R13021 VSS.n3277 VSS.n3276 3.4105
R13022 VSS.n3276 VSS.n3275 3.4105
R13023 VSS.n3119 VSS.n3118 3.4105
R13024 VSS.n3119 VSS.n2964 3.4105
R13025 VSS.n3112 VSS.n3111 3.4105
R13026 VSS.n3117 VSS.n3116 3.4105
R13027 VSS.n3116 VSS.n3115 3.4105
R13028 VSS.n3092 VSS.n3091 3.4105
R13029 VSS.n3092 VSS.n3004 3.4105
R13030 VSS.n3090 VSS.n3089 3.4105
R13031 VSS.n3110 VSS.n3109 3.4105
R13032 VSS.n3109 VSS.n3108 3.4105
R13033 VSS.n3079 VSS.n3010 3.4105
R13034 VSS.n3010 VSS.n3009 3.4105
R13035 VSS.n3008 VSS.n3007 3.4105
R13036 VSS.n3087 VSS.n3086 3.4105
R13037 VSS.n3086 VSS.n3002 3.4105
R13038 VSS.n3057 VSS.n3056 3.4105
R13039 VSS.n3057 VSS.n3029 3.4105
R13040 VSS.n3078 VSS.n3077 3.4105
R13041 VSS.n3055 VSS.n3054 3.4105
R13042 VSS.n3054 VSS.n3053 3.4105
R13043 VSS.n3971 VSS.n3422 3.4105
R13044 VSS.n3977 VSS.n3422 3.4105
R13045 VSS.n3973 VSS.n3972 3.4105
R13046 VSS.n3997 VSS.n3996 3.4105
R13047 VSS.n3996 VSS.n3995 3.4105
R13048 VSS.n3954 VSS.n3952 3.4105
R13049 VSS.n3954 VSS.n3953 3.4105
R13050 VSS.n3970 VSS.n3969 3.4105
R13051 VSS.n3969 VSS.n3968 3.4105
R13052 VSS.n3932 VSS.n3931 3.4105
R13053 VSS.n3931 VSS.n3930 3.4105
R13054 VSS.n3435 VSS.n3434 3.4105
R13055 VSS.n3951 VSS.n3950 3.4105
R13056 VSS.n3950 VSS.n3949 3.4105
R13057 VSS.n3915 VSS.n3914 3.4105
R13058 VSS.n3934 VSS.n3933 3.4105
R13059 VSS.n3899 VSS.n3898 3.4105
R13060 VSS.n3898 VSS.n3897 3.4105
R13061 VSS.n3900 VSS.n3453 3.4105
R13062 VSS.n3903 VSS.n3448 3.4105
R13063 VSS.n3872 VSS.n3871 3.4105
R13064 VSS.n3872 VSS.n3471 3.4105
R13065 VSS.n3467 VSS.n3454 3.4105
R13066 VSS.n3879 VSS.n3467 3.4105
R13067 VSS.n3818 VSS.n3817 3.4105
R13068 VSS.n3818 VSS.n3481 3.4105
R13069 VSS.n3795 VSS.n3794 3.4105
R13070 VSS.n3816 VSS.n3815 3.4105
R13071 VSS.n3815 VSS.n3814 3.4105
R13072 VSS.n3785 VSS.n3511 3.4105
R13073 VSS.n3511 VSS.n3510 3.4105
R13074 VSS.n3787 VSS.n3786 3.4105
R13075 VSS.n3793 VSS.n3792 3.4105
R13076 VSS.n3792 VSS.n3791 3.4105
R13077 VSS.n3768 VSS.n3767 3.4105
R13078 VSS.n3768 VSS.n3525 3.4105
R13079 VSS.n3764 VSS.n3513 3.4105
R13080 VSS.n3784 VSS.n3783 3.4105
R13081 VSS.n3783 VSS.n3782 3.4105
R13082 VSS.n3747 VSS.n3746 3.4105
R13083 VSS.n3747 VSS.n3541 3.4105
R13084 VSS.n3763 VSS.n3762 3.4105
R13085 VSS.n3745 VSS.n3744 3.4105
R13086 VSS.n3744 VSS.n3743 3.4105
R13087 VSS.n3859 VSS.n3478 3.4105
R13088 VSS.n3833 VSS.n3478 3.4105
R13089 VSS.n3475 VSS.n3474 3.4105
R13090 VSS.n3869 VSS.n3868 3.4105
R13091 VSS.n3868 VSS.n3867 3.4105
R13092 VSS.n3711 VSS.n3710 3.4105
R13093 VSS.n3711 VSS.n3556 3.4105
R13094 VSS.n3704 VSS.n3703 3.4105
R13095 VSS.n3709 VSS.n3708 3.4105
R13096 VSS.n3708 VSS.n3707 3.4105
R13097 VSS.n3684 VSS.n3683 3.4105
R13098 VSS.n3684 VSS.n3596 3.4105
R13099 VSS.n3682 VSS.n3681 3.4105
R13100 VSS.n3702 VSS.n3701 3.4105
R13101 VSS.n3701 VSS.n3700 3.4105
R13102 VSS.n3671 VSS.n3602 3.4105
R13103 VSS.n3602 VSS.n3601 3.4105
R13104 VSS.n3600 VSS.n3599 3.4105
R13105 VSS.n3679 VSS.n3678 3.4105
R13106 VSS.n3678 VSS.n3594 3.4105
R13107 VSS.n3649 VSS.n3648 3.4105
R13108 VSS.n3649 VSS.n3621 3.4105
R13109 VSS.n3670 VSS.n3669 3.4105
R13110 VSS.n3647 VSS.n3646 3.4105
R13111 VSS.n3646 VSS.n3645 3.4105
R13112 VSS.n4563 VSS.n4014 3.4105
R13113 VSS.n4569 VSS.n4014 3.4105
R13114 VSS.n4565 VSS.n4564 3.4105
R13115 VSS.n4589 VSS.n4588 3.4105
R13116 VSS.n4588 VSS.n4587 3.4105
R13117 VSS.n4546 VSS.n4544 3.4105
R13118 VSS.n4546 VSS.n4545 3.4105
R13119 VSS.n4562 VSS.n4561 3.4105
R13120 VSS.n4561 VSS.n4560 3.4105
R13121 VSS.n4524 VSS.n4523 3.4105
R13122 VSS.n4523 VSS.n4522 3.4105
R13123 VSS.n4027 VSS.n4026 3.4105
R13124 VSS.n4543 VSS.n4542 3.4105
R13125 VSS.n4542 VSS.n4541 3.4105
R13126 VSS.n4507 VSS.n4506 3.4105
R13127 VSS.n4526 VSS.n4525 3.4105
R13128 VSS.n4491 VSS.n4490 3.4105
R13129 VSS.n4490 VSS.n4489 3.4105
R13130 VSS.n4492 VSS.n4045 3.4105
R13131 VSS.n4495 VSS.n4040 3.4105
R13132 VSS.n4464 VSS.n4463 3.4105
R13133 VSS.n4464 VSS.n4063 3.4105
R13134 VSS.n4059 VSS.n4046 3.4105
R13135 VSS.n4471 VSS.n4059 3.4105
R13136 VSS.n4410 VSS.n4409 3.4105
R13137 VSS.n4410 VSS.n4073 3.4105
R13138 VSS.n4387 VSS.n4386 3.4105
R13139 VSS.n4408 VSS.n4407 3.4105
R13140 VSS.n4407 VSS.n4406 3.4105
R13141 VSS.n4377 VSS.n4103 3.4105
R13142 VSS.n4103 VSS.n4102 3.4105
R13143 VSS.n4379 VSS.n4378 3.4105
R13144 VSS.n4385 VSS.n4384 3.4105
R13145 VSS.n4384 VSS.n4383 3.4105
R13146 VSS.n4360 VSS.n4359 3.4105
R13147 VSS.n4360 VSS.n4117 3.4105
R13148 VSS.n4356 VSS.n4105 3.4105
R13149 VSS.n4376 VSS.n4375 3.4105
R13150 VSS.n4375 VSS.n4374 3.4105
R13151 VSS.n4339 VSS.n4338 3.4105
R13152 VSS.n4339 VSS.n4133 3.4105
R13153 VSS.n4355 VSS.n4354 3.4105
R13154 VSS.n4337 VSS.n4336 3.4105
R13155 VSS.n4336 VSS.n4335 3.4105
R13156 VSS.n4451 VSS.n4070 3.4105
R13157 VSS.n4425 VSS.n4070 3.4105
R13158 VSS.n4067 VSS.n4066 3.4105
R13159 VSS.n4461 VSS.n4460 3.4105
R13160 VSS.n4460 VSS.n4459 3.4105
R13161 VSS.n4303 VSS.n4302 3.4105
R13162 VSS.n4303 VSS.n4148 3.4105
R13163 VSS.n4296 VSS.n4295 3.4105
R13164 VSS.n4301 VSS.n4300 3.4105
R13165 VSS.n4300 VSS.n4299 3.4105
R13166 VSS.n4276 VSS.n4275 3.4105
R13167 VSS.n4276 VSS.n4188 3.4105
R13168 VSS.n4274 VSS.n4273 3.4105
R13169 VSS.n4294 VSS.n4293 3.4105
R13170 VSS.n4293 VSS.n4292 3.4105
R13171 VSS.n4263 VSS.n4194 3.4105
R13172 VSS.n4194 VSS.n4193 3.4105
R13173 VSS.n4192 VSS.n4191 3.4105
R13174 VSS.n4271 VSS.n4270 3.4105
R13175 VSS.n4270 VSS.n4186 3.4105
R13176 VSS.n4241 VSS.n4240 3.4105
R13177 VSS.n4241 VSS.n4213 3.4105
R13178 VSS.n4262 VSS.n4261 3.4105
R13179 VSS.n4239 VSS.n4238 3.4105
R13180 VSS.n4238 VSS.n4237 3.4105
R13181 VSS.n5155 VSS.n4606 3.4105
R13182 VSS.n5161 VSS.n4606 3.4105
R13183 VSS.n5157 VSS.n5156 3.4105
R13184 VSS.n5181 VSS.n5180 3.4105
R13185 VSS.n5180 VSS.n5179 3.4105
R13186 VSS.n5138 VSS.n5136 3.4105
R13187 VSS.n5138 VSS.n5137 3.4105
R13188 VSS.n5154 VSS.n5153 3.4105
R13189 VSS.n5153 VSS.n5152 3.4105
R13190 VSS.n5116 VSS.n5115 3.4105
R13191 VSS.n5115 VSS.n5114 3.4105
R13192 VSS.n4619 VSS.n4618 3.4105
R13193 VSS.n5135 VSS.n5134 3.4105
R13194 VSS.n5134 VSS.n5133 3.4105
R13195 VSS.n5099 VSS.n5098 3.4105
R13196 VSS.n5118 VSS.n5117 3.4105
R13197 VSS.n5083 VSS.n5082 3.4105
R13198 VSS.n5082 VSS.n5081 3.4105
R13199 VSS.n5084 VSS.n4637 3.4105
R13200 VSS.n5087 VSS.n4632 3.4105
R13201 VSS.n5056 VSS.n5055 3.4105
R13202 VSS.n5056 VSS.n4655 3.4105
R13203 VSS.n4651 VSS.n4638 3.4105
R13204 VSS.n5063 VSS.n4651 3.4105
R13205 VSS.n5002 VSS.n5001 3.4105
R13206 VSS.n5002 VSS.n4665 3.4105
R13207 VSS.n4979 VSS.n4978 3.4105
R13208 VSS.n5000 VSS.n4999 3.4105
R13209 VSS.n4999 VSS.n4998 3.4105
R13210 VSS.n4969 VSS.n4695 3.4105
R13211 VSS.n4695 VSS.n4694 3.4105
R13212 VSS.n4971 VSS.n4970 3.4105
R13213 VSS.n4977 VSS.n4976 3.4105
R13214 VSS.n4976 VSS.n4975 3.4105
R13215 VSS.n4952 VSS.n4951 3.4105
R13216 VSS.n4952 VSS.n4709 3.4105
R13217 VSS.n4948 VSS.n4697 3.4105
R13218 VSS.n4968 VSS.n4967 3.4105
R13219 VSS.n4967 VSS.n4966 3.4105
R13220 VSS.n4931 VSS.n4930 3.4105
R13221 VSS.n4931 VSS.n4725 3.4105
R13222 VSS.n4947 VSS.n4946 3.4105
R13223 VSS.n4929 VSS.n4928 3.4105
R13224 VSS.n4928 VSS.n4927 3.4105
R13225 VSS.n5043 VSS.n4662 3.4105
R13226 VSS.n5017 VSS.n4662 3.4105
R13227 VSS.n4659 VSS.n4658 3.4105
R13228 VSS.n5053 VSS.n5052 3.4105
R13229 VSS.n5052 VSS.n5051 3.4105
R13230 VSS.n4895 VSS.n4894 3.4105
R13231 VSS.n4895 VSS.n4740 3.4105
R13232 VSS.n4888 VSS.n4887 3.4105
R13233 VSS.n4893 VSS.n4892 3.4105
R13234 VSS.n4892 VSS.n4891 3.4105
R13235 VSS.n4868 VSS.n4867 3.4105
R13236 VSS.n4868 VSS.n4780 3.4105
R13237 VSS.n4866 VSS.n4865 3.4105
R13238 VSS.n4886 VSS.n4885 3.4105
R13239 VSS.n4885 VSS.n4884 3.4105
R13240 VSS.n4855 VSS.n4786 3.4105
R13241 VSS.n4786 VSS.n4785 3.4105
R13242 VSS.n4784 VSS.n4783 3.4105
R13243 VSS.n4863 VSS.n4862 3.4105
R13244 VSS.n4862 VSS.n4778 3.4105
R13245 VSS.n4833 VSS.n4832 3.4105
R13246 VSS.n4833 VSS.n4805 3.4105
R13247 VSS.n4854 VSS.n4853 3.4105
R13248 VSS.n4831 VSS.n4830 3.4105
R13249 VSS.n4830 VSS.n4829 3.4105
R13250 VSS.n2811 VSS.n2765 3.4105
R13251 VSS.n2811 VSS.n2810 3.4105
R13252 VSS.n2814 VSS.n2813 3.4105
R13253 VSS.n5187 VSS.n5186 3.4105
R13254 VSS.n5188 VSS.n5187 3.4105
R13255 VSS.n5205 VSS.n5204 3.4105
R13256 VSS.n5206 VSS.n5205 3.4105
R13257 VSS.n5202 VSS.n5201 3.4105
R13258 VSS.n5201 VSS.n5200 3.4105
R13259 VSS.n5220 VSS.n5219 3.4105
R13260 VSS.n5219 VSS.n5218 3.4105
R13261 VSS.n2763 VSS.n2762 3.4105
R13262 VSS.n2764 VSS.n2756 3.4105
R13263 VSS.n2756 VSS.n2752 3.4105
R13264 VSS.n2746 VSS.n2745 3.4105
R13265 VSS.n5222 VSS.n5221 3.4105
R13266 VSS.n5237 VSS.n2714 3.4105
R13267 VSS.n5237 VSS.n5236 3.4105
R13268 VSS.n2731 VSS.n2707 3.4105
R13269 VSS.n2734 VSS.n2727 3.4105
R13270 VSS.n5253 VSS.n2697 3.4105
R13271 VSS.n5253 VSS.n5252 3.4105
R13272 VSS.n2713 VSS.n2712 3.4105
R13273 VSS.n2712 VSS.n2711 3.4105
R13274 VSS.n5276 VSS.n5275 3.4105
R13275 VSS.n5275 VSS.n5274 3.4105
R13276 VSS.n5283 VSS.n5282 3.4105
R13277 VSS.n5278 VSS.n5277 3.4105
R13278 VSS.n5279 VSS.n5278 3.4105
R13279 VSS.n5291 VSS.n5290 3.4105
R13280 VSS.n5290 VSS.n5289 3.4105
R13281 VSS.n2559 VSS.n2555 3.4105
R13282 VSS.n5285 VSS.n5284 3.4105
R13283 VSS.n5285 VSS.n2558 3.4105
R13284 VSS.n5299 VSS.n5298 3.4105
R13285 VSS.n5298 VSS.n5297 3.4105
R13286 VSS.n2554 VSS.n2552 3.4105
R13287 VSS.n5293 VSS.n5292 3.4105
R13288 VSS.n5293 VSS.n2550 3.4105
R13289 VSS.n5306 VSS.n5305 3.4105
R13290 VSS.n5305 VSS.n5304 3.4105
R13291 VSS.n5301 VSS.n5300 3.4105
R13292 VSS.n5307 VSS.n2539 3.4105
R13293 VSS.n2539 VSS.n2358 3.4105
R13294 VSS.n2688 VSS.n2686 3.4105
R13295 VSS.n2686 VSS.n2685 3.4105
R13296 VSS.n2680 VSS.n2679 3.4105
R13297 VSS.n2696 VSS.n2695 3.4105
R13298 VSS.n2695 VSS.n2694 3.4105
R13299 VSS.n2516 VSS.n2515 3.4105
R13300 VSS.n2516 VSS.n2361 3.4105
R13301 VSS.n2509 VSS.n2508 3.4105
R13302 VSS.n2514 VSS.n2513 3.4105
R13303 VSS.n2513 VSS.n2512 3.4105
R13304 VSS.n2489 VSS.n2488 3.4105
R13305 VSS.n2489 VSS.n2401 3.4105
R13306 VSS.n2487 VSS.n2486 3.4105
R13307 VSS.n2507 VSS.n2506 3.4105
R13308 VSS.n2506 VSS.n2505 3.4105
R13309 VSS.n2476 VSS.n2407 3.4105
R13310 VSS.n2407 VSS.n2406 3.4105
R13311 VSS.n2405 VSS.n2404 3.4105
R13312 VSS.n2484 VSS.n2483 3.4105
R13313 VSS.n2483 VSS.n2399 3.4105
R13314 VSS.n2454 VSS.n2453 3.4105
R13315 VSS.n2454 VSS.n2426 3.4105
R13316 VSS.n2475 VSS.n2474 3.4105
R13317 VSS.n2452 VSS.n2451 3.4105
R13318 VSS.n2451 VSS.n2450 3.4105
R13319 VSS.n5730 VSS.n5726 3.4105
R13320 VSS.n5736 VSS.n5730 3.4105
R13321 VSS.n5732 VSS.n5731 3.4105
R13322 VSS.n18887 VSS.n18886 3.4105
R13323 VSS.n18886 VSS.n18885 3.4105
R13324 VSS.n5778 VSS.n5777 3.4105
R13325 VSS.n5779 VSS.n5778 3.4105
R13326 VSS.n5775 VSS.n5774 3.4105
R13327 VSS.n5774 VSS.n5773 3.4105
R13328 VSS.n5793 VSS.n5792 3.4105
R13329 VSS.n5792 VSS.n5791 3.4105
R13330 VSS.n5724 VSS.n5723 3.4105
R13331 VSS.n5725 VSS.n5717 3.4105
R13332 VSS.n5717 VSS.n5713 3.4105
R13333 VSS.n5707 VSS.n5706 3.4105
R13334 VSS.n5795 VSS.n5794 3.4105
R13335 VSS.n5810 VSS.n5675 3.4105
R13336 VSS.n5810 VSS.n5809 3.4105
R13337 VSS.n5692 VSS.n5668 3.4105
R13338 VSS.n5695 VSS.n5688 3.4105
R13339 VSS.n5826 VSS.n5658 3.4105
R13340 VSS.n5826 VSS.n5825 3.4105
R13341 VSS.n5674 VSS.n5673 3.4105
R13342 VSS.n5673 VSS.n5672 3.4105
R13343 VSS.n5849 VSS.n5848 3.4105
R13344 VSS.n5848 VSS.n5847 3.4105
R13345 VSS.n5856 VSS.n5855 3.4105
R13346 VSS.n5851 VSS.n5850 3.4105
R13347 VSS.n5852 VSS.n5851 3.4105
R13348 VSS.n5864 VSS.n5863 3.4105
R13349 VSS.n5863 VSS.n5862 3.4105
R13350 VSS.n5520 VSS.n5516 3.4105
R13351 VSS.n5858 VSS.n5857 3.4105
R13352 VSS.n5858 VSS.n5519 3.4105
R13353 VSS.n5872 VSS.n5871 3.4105
R13354 VSS.n5871 VSS.n5870 3.4105
R13355 VSS.n5515 VSS.n5513 3.4105
R13356 VSS.n5866 VSS.n5865 3.4105
R13357 VSS.n5866 VSS.n5511 3.4105
R13358 VSS.n5879 VSS.n5878 3.4105
R13359 VSS.n5878 VSS.n5877 3.4105
R13360 VSS.n5874 VSS.n5873 3.4105
R13361 VSS.n5880 VSS.n5500 3.4105
R13362 VSS.n5500 VSS.n5319 3.4105
R13363 VSS.n5649 VSS.n5647 3.4105
R13364 VSS.n5647 VSS.n5646 3.4105
R13365 VSS.n5641 VSS.n5640 3.4105
R13366 VSS.n5657 VSS.n5656 3.4105
R13367 VSS.n5656 VSS.n5655 3.4105
R13368 VSS.n5477 VSS.n5476 3.4105
R13369 VSS.n5477 VSS.n5322 3.4105
R13370 VSS.n5470 VSS.n5469 3.4105
R13371 VSS.n5475 VSS.n5474 3.4105
R13372 VSS.n5474 VSS.n5473 3.4105
R13373 VSS.n5450 VSS.n5449 3.4105
R13374 VSS.n5450 VSS.n5362 3.4105
R13375 VSS.n5448 VSS.n5447 3.4105
R13376 VSS.n5468 VSS.n5467 3.4105
R13377 VSS.n5467 VSS.n5466 3.4105
R13378 VSS.n5437 VSS.n5368 3.4105
R13379 VSS.n5368 VSS.n5367 3.4105
R13380 VSS.n5366 VSS.n5365 3.4105
R13381 VSS.n5445 VSS.n5444 3.4105
R13382 VSS.n5444 VSS.n5360 3.4105
R13383 VSS.n5415 VSS.n5414 3.4105
R13384 VSS.n5415 VSS.n5387 3.4105
R13385 VSS.n5436 VSS.n5435 3.4105
R13386 VSS.n5413 VSS.n5412 3.4105
R13387 VSS.n5412 VSS.n5411 3.4105
R13388 VSS.n6345 VSS.n6299 3.4105
R13389 VSS.n6345 VSS.n6344 3.4105
R13390 VSS.n6348 VSS.n6347 3.4105
R13391 VSS.n6352 VSS.n6351 3.4105
R13392 VSS.n6353 VSS.n6352 3.4105
R13393 VSS.n6370 VSS.n6369 3.4105
R13394 VSS.n6371 VSS.n6370 3.4105
R13395 VSS.n6367 VSS.n6366 3.4105
R13396 VSS.n6366 VSS.n6365 3.4105
R13397 VSS.n6385 VSS.n6384 3.4105
R13398 VSS.n6384 VSS.n6383 3.4105
R13399 VSS.n6297 VSS.n6296 3.4105
R13400 VSS.n6298 VSS.n6290 3.4105
R13401 VSS.n6290 VSS.n6286 3.4105
R13402 VSS.n6280 VSS.n6279 3.4105
R13403 VSS.n6387 VSS.n6386 3.4105
R13404 VSS.n6402 VSS.n6248 3.4105
R13405 VSS.n6402 VSS.n6401 3.4105
R13406 VSS.n6265 VSS.n6241 3.4105
R13407 VSS.n6268 VSS.n6261 3.4105
R13408 VSS.n6418 VSS.n6231 3.4105
R13409 VSS.n6418 VSS.n6417 3.4105
R13410 VSS.n6247 VSS.n6246 3.4105
R13411 VSS.n6246 VSS.n6245 3.4105
R13412 VSS.n6441 VSS.n6440 3.4105
R13413 VSS.n6440 VSS.n6439 3.4105
R13414 VSS.n6448 VSS.n6447 3.4105
R13415 VSS.n6443 VSS.n6442 3.4105
R13416 VSS.n6444 VSS.n6443 3.4105
R13417 VSS.n6456 VSS.n6455 3.4105
R13418 VSS.n6455 VSS.n6454 3.4105
R13419 VSS.n6093 VSS.n6089 3.4105
R13420 VSS.n6450 VSS.n6449 3.4105
R13421 VSS.n6450 VSS.n6092 3.4105
R13422 VSS.n6464 VSS.n6463 3.4105
R13423 VSS.n6463 VSS.n6462 3.4105
R13424 VSS.n6088 VSS.n6086 3.4105
R13425 VSS.n6458 VSS.n6457 3.4105
R13426 VSS.n6458 VSS.n6084 3.4105
R13427 VSS.n6471 VSS.n6470 3.4105
R13428 VSS.n6470 VSS.n6469 3.4105
R13429 VSS.n6466 VSS.n6465 3.4105
R13430 VSS.n6472 VSS.n6073 3.4105
R13431 VSS.n6073 VSS.n5892 3.4105
R13432 VSS.n6222 VSS.n6220 3.4105
R13433 VSS.n6220 VSS.n6219 3.4105
R13434 VSS.n6214 VSS.n6213 3.4105
R13435 VSS.n6230 VSS.n6229 3.4105
R13436 VSS.n6229 VSS.n6228 3.4105
R13437 VSS.n6050 VSS.n6049 3.4105
R13438 VSS.n6050 VSS.n5895 3.4105
R13439 VSS.n6043 VSS.n6042 3.4105
R13440 VSS.n6048 VSS.n6047 3.4105
R13441 VSS.n6047 VSS.n6046 3.4105
R13442 VSS.n6023 VSS.n6022 3.4105
R13443 VSS.n6023 VSS.n5935 3.4105
R13444 VSS.n6021 VSS.n6020 3.4105
R13445 VSS.n6041 VSS.n6040 3.4105
R13446 VSS.n6040 VSS.n6039 3.4105
R13447 VSS.n6010 VSS.n5941 3.4105
R13448 VSS.n5941 VSS.n5940 3.4105
R13449 VSS.n5939 VSS.n5938 3.4105
R13450 VSS.n6018 VSS.n6017 3.4105
R13451 VSS.n6017 VSS.n5933 3.4105
R13452 VSS.n5988 VSS.n5987 3.4105
R13453 VSS.n5988 VSS.n5960 3.4105
R13454 VSS.n6009 VSS.n6008 3.4105
R13455 VSS.n5986 VSS.n5985 3.4105
R13456 VSS.n5985 VSS.n5984 3.4105
R13457 VSS.n8112 VSS.n7563 3.4105
R13458 VSS.n8118 VSS.n7563 3.4105
R13459 VSS.n8114 VSS.n8113 3.4105
R13460 VSS.n8138 VSS.n8137 3.4105
R13461 VSS.n8137 VSS.n8136 3.4105
R13462 VSS.n8095 VSS.n8093 3.4105
R13463 VSS.n8095 VSS.n8094 3.4105
R13464 VSS.n8111 VSS.n8110 3.4105
R13465 VSS.n8110 VSS.n8109 3.4105
R13466 VSS.n8073 VSS.n8072 3.4105
R13467 VSS.n8072 VSS.n8071 3.4105
R13468 VSS.n7576 VSS.n7575 3.4105
R13469 VSS.n8092 VSS.n8091 3.4105
R13470 VSS.n8091 VSS.n8090 3.4105
R13471 VSS.n8056 VSS.n8055 3.4105
R13472 VSS.n8075 VSS.n8074 3.4105
R13473 VSS.n8040 VSS.n8039 3.4105
R13474 VSS.n8039 VSS.n8038 3.4105
R13475 VSS.n8041 VSS.n7594 3.4105
R13476 VSS.n8044 VSS.n7589 3.4105
R13477 VSS.n8013 VSS.n8012 3.4105
R13478 VSS.n8013 VSS.n7612 3.4105
R13479 VSS.n7608 VSS.n7595 3.4105
R13480 VSS.n8020 VSS.n7608 3.4105
R13481 VSS.n7959 VSS.n7958 3.4105
R13482 VSS.n7959 VSS.n7622 3.4105
R13483 VSS.n7936 VSS.n7935 3.4105
R13484 VSS.n7957 VSS.n7956 3.4105
R13485 VSS.n7956 VSS.n7955 3.4105
R13486 VSS.n7926 VSS.n7652 3.4105
R13487 VSS.n7652 VSS.n7651 3.4105
R13488 VSS.n7928 VSS.n7927 3.4105
R13489 VSS.n7934 VSS.n7933 3.4105
R13490 VSS.n7933 VSS.n7932 3.4105
R13491 VSS.n7909 VSS.n7908 3.4105
R13492 VSS.n7909 VSS.n7666 3.4105
R13493 VSS.n7905 VSS.n7654 3.4105
R13494 VSS.n7925 VSS.n7924 3.4105
R13495 VSS.n7924 VSS.n7923 3.4105
R13496 VSS.n7888 VSS.n7887 3.4105
R13497 VSS.n7888 VSS.n7682 3.4105
R13498 VSS.n7904 VSS.n7903 3.4105
R13499 VSS.n7886 VSS.n7885 3.4105
R13500 VSS.n7885 VSS.n7884 3.4105
R13501 VSS.n8000 VSS.n7619 3.4105
R13502 VSS.n7974 VSS.n7619 3.4105
R13503 VSS.n7616 VSS.n7615 3.4105
R13504 VSS.n8010 VSS.n8009 3.4105
R13505 VSS.n8009 VSS.n8008 3.4105
R13506 VSS.n7852 VSS.n7851 3.4105
R13507 VSS.n7852 VSS.n7697 3.4105
R13508 VSS.n7845 VSS.n7844 3.4105
R13509 VSS.n7850 VSS.n7849 3.4105
R13510 VSS.n7849 VSS.n7848 3.4105
R13511 VSS.n7825 VSS.n7824 3.4105
R13512 VSS.n7825 VSS.n7737 3.4105
R13513 VSS.n7823 VSS.n7822 3.4105
R13514 VSS.n7843 VSS.n7842 3.4105
R13515 VSS.n7842 VSS.n7841 3.4105
R13516 VSS.n7812 VSS.n7743 3.4105
R13517 VSS.n7743 VSS.n7742 3.4105
R13518 VSS.n7741 VSS.n7740 3.4105
R13519 VSS.n7820 VSS.n7819 3.4105
R13520 VSS.n7819 VSS.n7735 3.4105
R13521 VSS.n7790 VSS.n7789 3.4105
R13522 VSS.n7790 VSS.n7762 3.4105
R13523 VSS.n7811 VSS.n7810 3.4105
R13524 VSS.n7788 VSS.n7787 3.4105
R13525 VSS.n7787 VSS.n7786 3.4105
R13526 VSS.n8704 VSS.n8155 3.4105
R13527 VSS.n8710 VSS.n8155 3.4105
R13528 VSS.n8706 VSS.n8705 3.4105
R13529 VSS.n8730 VSS.n8729 3.4105
R13530 VSS.n8729 VSS.n8728 3.4105
R13531 VSS.n8687 VSS.n8685 3.4105
R13532 VSS.n8687 VSS.n8686 3.4105
R13533 VSS.n8703 VSS.n8702 3.4105
R13534 VSS.n8702 VSS.n8701 3.4105
R13535 VSS.n8665 VSS.n8664 3.4105
R13536 VSS.n8664 VSS.n8663 3.4105
R13537 VSS.n8168 VSS.n8167 3.4105
R13538 VSS.n8684 VSS.n8683 3.4105
R13539 VSS.n8683 VSS.n8682 3.4105
R13540 VSS.n8648 VSS.n8647 3.4105
R13541 VSS.n8667 VSS.n8666 3.4105
R13542 VSS.n8632 VSS.n8631 3.4105
R13543 VSS.n8631 VSS.n8630 3.4105
R13544 VSS.n8633 VSS.n8186 3.4105
R13545 VSS.n8636 VSS.n8181 3.4105
R13546 VSS.n8605 VSS.n8604 3.4105
R13547 VSS.n8605 VSS.n8204 3.4105
R13548 VSS.n8200 VSS.n8187 3.4105
R13549 VSS.n8612 VSS.n8200 3.4105
R13550 VSS.n8551 VSS.n8550 3.4105
R13551 VSS.n8551 VSS.n8214 3.4105
R13552 VSS.n8528 VSS.n8527 3.4105
R13553 VSS.n8549 VSS.n8548 3.4105
R13554 VSS.n8548 VSS.n8547 3.4105
R13555 VSS.n8518 VSS.n8244 3.4105
R13556 VSS.n8244 VSS.n8243 3.4105
R13557 VSS.n8520 VSS.n8519 3.4105
R13558 VSS.n8526 VSS.n8525 3.4105
R13559 VSS.n8525 VSS.n8524 3.4105
R13560 VSS.n8501 VSS.n8500 3.4105
R13561 VSS.n8501 VSS.n8258 3.4105
R13562 VSS.n8497 VSS.n8246 3.4105
R13563 VSS.n8517 VSS.n8516 3.4105
R13564 VSS.n8516 VSS.n8515 3.4105
R13565 VSS.n8480 VSS.n8479 3.4105
R13566 VSS.n8480 VSS.n8274 3.4105
R13567 VSS.n8496 VSS.n8495 3.4105
R13568 VSS.n8478 VSS.n8477 3.4105
R13569 VSS.n8477 VSS.n8476 3.4105
R13570 VSS.n8592 VSS.n8211 3.4105
R13571 VSS.n8566 VSS.n8211 3.4105
R13572 VSS.n8208 VSS.n8207 3.4105
R13573 VSS.n8602 VSS.n8601 3.4105
R13574 VSS.n8601 VSS.n8600 3.4105
R13575 VSS.n8444 VSS.n8443 3.4105
R13576 VSS.n8444 VSS.n8289 3.4105
R13577 VSS.n8437 VSS.n8436 3.4105
R13578 VSS.n8442 VSS.n8441 3.4105
R13579 VSS.n8441 VSS.n8440 3.4105
R13580 VSS.n8417 VSS.n8416 3.4105
R13581 VSS.n8417 VSS.n8329 3.4105
R13582 VSS.n8415 VSS.n8414 3.4105
R13583 VSS.n8435 VSS.n8434 3.4105
R13584 VSS.n8434 VSS.n8433 3.4105
R13585 VSS.n8404 VSS.n8335 3.4105
R13586 VSS.n8335 VSS.n8334 3.4105
R13587 VSS.n8333 VSS.n8332 3.4105
R13588 VSS.n8412 VSS.n8411 3.4105
R13589 VSS.n8411 VSS.n8327 3.4105
R13590 VSS.n8382 VSS.n8381 3.4105
R13591 VSS.n8382 VSS.n8354 3.4105
R13592 VSS.n8403 VSS.n8402 3.4105
R13593 VSS.n8380 VSS.n8379 3.4105
R13594 VSS.n8379 VSS.n8378 3.4105
R13595 VSS.n9296 VSS.n8747 3.4105
R13596 VSS.n9302 VSS.n8747 3.4105
R13597 VSS.n9298 VSS.n9297 3.4105
R13598 VSS.n9322 VSS.n9321 3.4105
R13599 VSS.n9321 VSS.n9320 3.4105
R13600 VSS.n9279 VSS.n9277 3.4105
R13601 VSS.n9279 VSS.n9278 3.4105
R13602 VSS.n9295 VSS.n9294 3.4105
R13603 VSS.n9294 VSS.n9293 3.4105
R13604 VSS.n9257 VSS.n9256 3.4105
R13605 VSS.n9256 VSS.n9255 3.4105
R13606 VSS.n8760 VSS.n8759 3.4105
R13607 VSS.n9276 VSS.n9275 3.4105
R13608 VSS.n9275 VSS.n9274 3.4105
R13609 VSS.n9240 VSS.n9239 3.4105
R13610 VSS.n9259 VSS.n9258 3.4105
R13611 VSS.n9224 VSS.n9223 3.4105
R13612 VSS.n9223 VSS.n9222 3.4105
R13613 VSS.n9225 VSS.n8778 3.4105
R13614 VSS.n9228 VSS.n8773 3.4105
R13615 VSS.n9197 VSS.n9196 3.4105
R13616 VSS.n9197 VSS.n8796 3.4105
R13617 VSS.n8792 VSS.n8779 3.4105
R13618 VSS.n9204 VSS.n8792 3.4105
R13619 VSS.n9143 VSS.n9142 3.4105
R13620 VSS.n9143 VSS.n8806 3.4105
R13621 VSS.n9120 VSS.n9119 3.4105
R13622 VSS.n9141 VSS.n9140 3.4105
R13623 VSS.n9140 VSS.n9139 3.4105
R13624 VSS.n9110 VSS.n8836 3.4105
R13625 VSS.n8836 VSS.n8835 3.4105
R13626 VSS.n9112 VSS.n9111 3.4105
R13627 VSS.n9118 VSS.n9117 3.4105
R13628 VSS.n9117 VSS.n9116 3.4105
R13629 VSS.n9093 VSS.n9092 3.4105
R13630 VSS.n9093 VSS.n8850 3.4105
R13631 VSS.n9089 VSS.n8838 3.4105
R13632 VSS.n9109 VSS.n9108 3.4105
R13633 VSS.n9108 VSS.n9107 3.4105
R13634 VSS.n9072 VSS.n9071 3.4105
R13635 VSS.n9072 VSS.n8866 3.4105
R13636 VSS.n9088 VSS.n9087 3.4105
R13637 VSS.n9070 VSS.n9069 3.4105
R13638 VSS.n9069 VSS.n9068 3.4105
R13639 VSS.n9184 VSS.n8803 3.4105
R13640 VSS.n9158 VSS.n8803 3.4105
R13641 VSS.n8800 VSS.n8799 3.4105
R13642 VSS.n9194 VSS.n9193 3.4105
R13643 VSS.n9193 VSS.n9192 3.4105
R13644 VSS.n9036 VSS.n9035 3.4105
R13645 VSS.n9036 VSS.n8881 3.4105
R13646 VSS.n9029 VSS.n9028 3.4105
R13647 VSS.n9034 VSS.n9033 3.4105
R13648 VSS.n9033 VSS.n9032 3.4105
R13649 VSS.n9009 VSS.n9008 3.4105
R13650 VSS.n9009 VSS.n8921 3.4105
R13651 VSS.n9007 VSS.n9006 3.4105
R13652 VSS.n9027 VSS.n9026 3.4105
R13653 VSS.n9026 VSS.n9025 3.4105
R13654 VSS.n8996 VSS.n8927 3.4105
R13655 VSS.n8927 VSS.n8926 3.4105
R13656 VSS.n8925 VSS.n8924 3.4105
R13657 VSS.n9004 VSS.n9003 3.4105
R13658 VSS.n9003 VSS.n8919 3.4105
R13659 VSS.n8974 VSS.n8973 3.4105
R13660 VSS.n8974 VSS.n8946 3.4105
R13661 VSS.n8995 VSS.n8994 3.4105
R13662 VSS.n8972 VSS.n8971 3.4105
R13663 VSS.n8971 VSS.n8970 3.4105
R13664 VSS.n10480 VSS.n9931 3.4105
R13665 VSS.n10486 VSS.n9931 3.4105
R13666 VSS.n10482 VSS.n10481 3.4105
R13667 VSS.n10506 VSS.n10505 3.4105
R13668 VSS.n10505 VSS.n10504 3.4105
R13669 VSS.n10463 VSS.n10461 3.4105
R13670 VSS.n10463 VSS.n10462 3.4105
R13671 VSS.n10479 VSS.n10478 3.4105
R13672 VSS.n10478 VSS.n10477 3.4105
R13673 VSS.n10441 VSS.n10440 3.4105
R13674 VSS.n10440 VSS.n10439 3.4105
R13675 VSS.n9944 VSS.n9943 3.4105
R13676 VSS.n10460 VSS.n10459 3.4105
R13677 VSS.n10459 VSS.n10458 3.4105
R13678 VSS.n10424 VSS.n10423 3.4105
R13679 VSS.n10443 VSS.n10442 3.4105
R13680 VSS.n10408 VSS.n10407 3.4105
R13681 VSS.n10407 VSS.n10406 3.4105
R13682 VSS.n10409 VSS.n9962 3.4105
R13683 VSS.n10412 VSS.n9957 3.4105
R13684 VSS.n10381 VSS.n10380 3.4105
R13685 VSS.n10381 VSS.n9980 3.4105
R13686 VSS.n9976 VSS.n9963 3.4105
R13687 VSS.n10388 VSS.n9976 3.4105
R13688 VSS.n10327 VSS.n10326 3.4105
R13689 VSS.n10327 VSS.n9990 3.4105
R13690 VSS.n10304 VSS.n10303 3.4105
R13691 VSS.n10325 VSS.n10324 3.4105
R13692 VSS.n10324 VSS.n10323 3.4105
R13693 VSS.n10294 VSS.n10020 3.4105
R13694 VSS.n10020 VSS.n10019 3.4105
R13695 VSS.n10296 VSS.n10295 3.4105
R13696 VSS.n10302 VSS.n10301 3.4105
R13697 VSS.n10301 VSS.n10300 3.4105
R13698 VSS.n10277 VSS.n10276 3.4105
R13699 VSS.n10277 VSS.n10034 3.4105
R13700 VSS.n10273 VSS.n10022 3.4105
R13701 VSS.n10293 VSS.n10292 3.4105
R13702 VSS.n10292 VSS.n10291 3.4105
R13703 VSS.n10256 VSS.n10255 3.4105
R13704 VSS.n10256 VSS.n10050 3.4105
R13705 VSS.n10272 VSS.n10271 3.4105
R13706 VSS.n10254 VSS.n10253 3.4105
R13707 VSS.n10253 VSS.n10252 3.4105
R13708 VSS.n10368 VSS.n9987 3.4105
R13709 VSS.n10342 VSS.n9987 3.4105
R13710 VSS.n9984 VSS.n9983 3.4105
R13711 VSS.n10378 VSS.n10377 3.4105
R13712 VSS.n10377 VSS.n10376 3.4105
R13713 VSS.n10220 VSS.n10219 3.4105
R13714 VSS.n10220 VSS.n10065 3.4105
R13715 VSS.n10213 VSS.n10212 3.4105
R13716 VSS.n10218 VSS.n10217 3.4105
R13717 VSS.n10217 VSS.n10216 3.4105
R13718 VSS.n10193 VSS.n10192 3.4105
R13719 VSS.n10193 VSS.n10105 3.4105
R13720 VSS.n10191 VSS.n10190 3.4105
R13721 VSS.n10211 VSS.n10210 3.4105
R13722 VSS.n10210 VSS.n10209 3.4105
R13723 VSS.n10180 VSS.n10111 3.4105
R13724 VSS.n10111 VSS.n10110 3.4105
R13725 VSS.n10109 VSS.n10108 3.4105
R13726 VSS.n10188 VSS.n10187 3.4105
R13727 VSS.n10187 VSS.n10103 3.4105
R13728 VSS.n10158 VSS.n10157 3.4105
R13729 VSS.n10158 VSS.n10130 3.4105
R13730 VSS.n10179 VSS.n10178 3.4105
R13731 VSS.n10156 VSS.n10155 3.4105
R13732 VSS.n10155 VSS.n10154 3.4105
R13733 VSS.n11072 VSS.n10523 3.4105
R13734 VSS.n11078 VSS.n10523 3.4105
R13735 VSS.n11074 VSS.n11073 3.4105
R13736 VSS.n11098 VSS.n11097 3.4105
R13737 VSS.n11097 VSS.n11096 3.4105
R13738 VSS.n11055 VSS.n11053 3.4105
R13739 VSS.n11055 VSS.n11054 3.4105
R13740 VSS.n11071 VSS.n11070 3.4105
R13741 VSS.n11070 VSS.n11069 3.4105
R13742 VSS.n11033 VSS.n11032 3.4105
R13743 VSS.n11032 VSS.n11031 3.4105
R13744 VSS.n10536 VSS.n10535 3.4105
R13745 VSS.n11052 VSS.n11051 3.4105
R13746 VSS.n11051 VSS.n11050 3.4105
R13747 VSS.n11016 VSS.n11015 3.4105
R13748 VSS.n11035 VSS.n11034 3.4105
R13749 VSS.n11000 VSS.n10999 3.4105
R13750 VSS.n10999 VSS.n10998 3.4105
R13751 VSS.n11001 VSS.n10554 3.4105
R13752 VSS.n11004 VSS.n10549 3.4105
R13753 VSS.n10973 VSS.n10972 3.4105
R13754 VSS.n10973 VSS.n10572 3.4105
R13755 VSS.n10568 VSS.n10555 3.4105
R13756 VSS.n10980 VSS.n10568 3.4105
R13757 VSS.n10919 VSS.n10918 3.4105
R13758 VSS.n10919 VSS.n10582 3.4105
R13759 VSS.n10896 VSS.n10895 3.4105
R13760 VSS.n10917 VSS.n10916 3.4105
R13761 VSS.n10916 VSS.n10915 3.4105
R13762 VSS.n10886 VSS.n10612 3.4105
R13763 VSS.n10612 VSS.n10611 3.4105
R13764 VSS.n10888 VSS.n10887 3.4105
R13765 VSS.n10894 VSS.n10893 3.4105
R13766 VSS.n10893 VSS.n10892 3.4105
R13767 VSS.n10869 VSS.n10868 3.4105
R13768 VSS.n10869 VSS.n10626 3.4105
R13769 VSS.n10865 VSS.n10614 3.4105
R13770 VSS.n10885 VSS.n10884 3.4105
R13771 VSS.n10884 VSS.n10883 3.4105
R13772 VSS.n10848 VSS.n10847 3.4105
R13773 VSS.n10848 VSS.n10642 3.4105
R13774 VSS.n10864 VSS.n10863 3.4105
R13775 VSS.n10846 VSS.n10845 3.4105
R13776 VSS.n10845 VSS.n10844 3.4105
R13777 VSS.n10960 VSS.n10579 3.4105
R13778 VSS.n10934 VSS.n10579 3.4105
R13779 VSS.n10576 VSS.n10575 3.4105
R13780 VSS.n10970 VSS.n10969 3.4105
R13781 VSS.n10969 VSS.n10968 3.4105
R13782 VSS.n10812 VSS.n10811 3.4105
R13783 VSS.n10812 VSS.n10657 3.4105
R13784 VSS.n10805 VSS.n10804 3.4105
R13785 VSS.n10810 VSS.n10809 3.4105
R13786 VSS.n10809 VSS.n10808 3.4105
R13787 VSS.n10785 VSS.n10784 3.4105
R13788 VSS.n10785 VSS.n10697 3.4105
R13789 VSS.n10783 VSS.n10782 3.4105
R13790 VSS.n10803 VSS.n10802 3.4105
R13791 VSS.n10802 VSS.n10801 3.4105
R13792 VSS.n10772 VSS.n10703 3.4105
R13793 VSS.n10703 VSS.n10702 3.4105
R13794 VSS.n10701 VSS.n10700 3.4105
R13795 VSS.n10780 VSS.n10779 3.4105
R13796 VSS.n10779 VSS.n10695 3.4105
R13797 VSS.n10750 VSS.n10749 3.4105
R13798 VSS.n10750 VSS.n10722 3.4105
R13799 VSS.n10771 VSS.n10770 3.4105
R13800 VSS.n10748 VSS.n10747 3.4105
R13801 VSS.n10747 VSS.n10746 3.4105
R13802 VSS.n11664 VSS.n11115 3.4105
R13803 VSS.n11670 VSS.n11115 3.4105
R13804 VSS.n11666 VSS.n11665 3.4105
R13805 VSS.n11690 VSS.n11689 3.4105
R13806 VSS.n11689 VSS.n11688 3.4105
R13807 VSS.n11647 VSS.n11645 3.4105
R13808 VSS.n11647 VSS.n11646 3.4105
R13809 VSS.n11663 VSS.n11662 3.4105
R13810 VSS.n11662 VSS.n11661 3.4105
R13811 VSS.n11625 VSS.n11624 3.4105
R13812 VSS.n11624 VSS.n11623 3.4105
R13813 VSS.n11128 VSS.n11127 3.4105
R13814 VSS.n11644 VSS.n11643 3.4105
R13815 VSS.n11643 VSS.n11642 3.4105
R13816 VSS.n11608 VSS.n11607 3.4105
R13817 VSS.n11627 VSS.n11626 3.4105
R13818 VSS.n11592 VSS.n11591 3.4105
R13819 VSS.n11591 VSS.n11590 3.4105
R13820 VSS.n11593 VSS.n11146 3.4105
R13821 VSS.n11596 VSS.n11141 3.4105
R13822 VSS.n11565 VSS.n11564 3.4105
R13823 VSS.n11565 VSS.n11164 3.4105
R13824 VSS.n11160 VSS.n11147 3.4105
R13825 VSS.n11572 VSS.n11160 3.4105
R13826 VSS.n11511 VSS.n11510 3.4105
R13827 VSS.n11511 VSS.n11174 3.4105
R13828 VSS.n11488 VSS.n11487 3.4105
R13829 VSS.n11509 VSS.n11508 3.4105
R13830 VSS.n11508 VSS.n11507 3.4105
R13831 VSS.n11478 VSS.n11204 3.4105
R13832 VSS.n11204 VSS.n11203 3.4105
R13833 VSS.n11480 VSS.n11479 3.4105
R13834 VSS.n11486 VSS.n11485 3.4105
R13835 VSS.n11485 VSS.n11484 3.4105
R13836 VSS.n11461 VSS.n11460 3.4105
R13837 VSS.n11461 VSS.n11218 3.4105
R13838 VSS.n11457 VSS.n11206 3.4105
R13839 VSS.n11477 VSS.n11476 3.4105
R13840 VSS.n11476 VSS.n11475 3.4105
R13841 VSS.n11440 VSS.n11439 3.4105
R13842 VSS.n11440 VSS.n11234 3.4105
R13843 VSS.n11456 VSS.n11455 3.4105
R13844 VSS.n11438 VSS.n11437 3.4105
R13845 VSS.n11437 VSS.n11436 3.4105
R13846 VSS.n11552 VSS.n11171 3.4105
R13847 VSS.n11526 VSS.n11171 3.4105
R13848 VSS.n11168 VSS.n11167 3.4105
R13849 VSS.n11562 VSS.n11561 3.4105
R13850 VSS.n11561 VSS.n11560 3.4105
R13851 VSS.n11404 VSS.n11403 3.4105
R13852 VSS.n11404 VSS.n11249 3.4105
R13853 VSS.n11397 VSS.n11396 3.4105
R13854 VSS.n11402 VSS.n11401 3.4105
R13855 VSS.n11401 VSS.n11400 3.4105
R13856 VSS.n11377 VSS.n11376 3.4105
R13857 VSS.n11377 VSS.n11289 3.4105
R13858 VSS.n11375 VSS.n11374 3.4105
R13859 VSS.n11395 VSS.n11394 3.4105
R13860 VSS.n11394 VSS.n11393 3.4105
R13861 VSS.n11364 VSS.n11295 3.4105
R13862 VSS.n11295 VSS.n11294 3.4105
R13863 VSS.n11293 VSS.n11292 3.4105
R13864 VSS.n11372 VSS.n11371 3.4105
R13865 VSS.n11371 VSS.n11287 3.4105
R13866 VSS.n11342 VSS.n11341 3.4105
R13867 VSS.n11342 VSS.n11314 3.4105
R13868 VSS.n11363 VSS.n11362 3.4105
R13869 VSS.n11340 VSS.n11339 3.4105
R13870 VSS.n11339 VSS.n11338 3.4105
R13871 VSS.n12256 VSS.n11707 3.4105
R13872 VSS.n12262 VSS.n11707 3.4105
R13873 VSS.n12258 VSS.n12257 3.4105
R13874 VSS.n12282 VSS.n12281 3.4105
R13875 VSS.n12281 VSS.n12280 3.4105
R13876 VSS.n12239 VSS.n12237 3.4105
R13877 VSS.n12239 VSS.n12238 3.4105
R13878 VSS.n12255 VSS.n12254 3.4105
R13879 VSS.n12254 VSS.n12253 3.4105
R13880 VSS.n12217 VSS.n12216 3.4105
R13881 VSS.n12216 VSS.n12215 3.4105
R13882 VSS.n11720 VSS.n11719 3.4105
R13883 VSS.n12236 VSS.n12235 3.4105
R13884 VSS.n12235 VSS.n12234 3.4105
R13885 VSS.n12200 VSS.n12199 3.4105
R13886 VSS.n12219 VSS.n12218 3.4105
R13887 VSS.n12184 VSS.n12183 3.4105
R13888 VSS.n12183 VSS.n12182 3.4105
R13889 VSS.n12185 VSS.n11738 3.4105
R13890 VSS.n12188 VSS.n11733 3.4105
R13891 VSS.n12157 VSS.n12156 3.4105
R13892 VSS.n12157 VSS.n11756 3.4105
R13893 VSS.n11752 VSS.n11739 3.4105
R13894 VSS.n12164 VSS.n11752 3.4105
R13895 VSS.n12103 VSS.n12102 3.4105
R13896 VSS.n12103 VSS.n11766 3.4105
R13897 VSS.n12080 VSS.n12079 3.4105
R13898 VSS.n12101 VSS.n12100 3.4105
R13899 VSS.n12100 VSS.n12099 3.4105
R13900 VSS.n12070 VSS.n11796 3.4105
R13901 VSS.n11796 VSS.n11795 3.4105
R13902 VSS.n12072 VSS.n12071 3.4105
R13903 VSS.n12078 VSS.n12077 3.4105
R13904 VSS.n12077 VSS.n12076 3.4105
R13905 VSS.n12053 VSS.n12052 3.4105
R13906 VSS.n12053 VSS.n11810 3.4105
R13907 VSS.n12049 VSS.n11798 3.4105
R13908 VSS.n12069 VSS.n12068 3.4105
R13909 VSS.n12068 VSS.n12067 3.4105
R13910 VSS.n12032 VSS.n12031 3.4105
R13911 VSS.n12032 VSS.n11826 3.4105
R13912 VSS.n12048 VSS.n12047 3.4105
R13913 VSS.n12030 VSS.n12029 3.4105
R13914 VSS.n12029 VSS.n12028 3.4105
R13915 VSS.n12144 VSS.n11763 3.4105
R13916 VSS.n12118 VSS.n11763 3.4105
R13917 VSS.n11760 VSS.n11759 3.4105
R13918 VSS.n12154 VSS.n12153 3.4105
R13919 VSS.n12153 VSS.n12152 3.4105
R13920 VSS.n11996 VSS.n11995 3.4105
R13921 VSS.n11996 VSS.n11841 3.4105
R13922 VSS.n11989 VSS.n11988 3.4105
R13923 VSS.n11994 VSS.n11993 3.4105
R13924 VSS.n11993 VSS.n11992 3.4105
R13925 VSS.n11969 VSS.n11968 3.4105
R13926 VSS.n11969 VSS.n11881 3.4105
R13927 VSS.n11967 VSS.n11966 3.4105
R13928 VSS.n11987 VSS.n11986 3.4105
R13929 VSS.n11986 VSS.n11985 3.4105
R13930 VSS.n11956 VSS.n11887 3.4105
R13931 VSS.n11887 VSS.n11886 3.4105
R13932 VSS.n11885 VSS.n11884 3.4105
R13933 VSS.n11964 VSS.n11963 3.4105
R13934 VSS.n11963 VSS.n11879 3.4105
R13935 VSS.n11934 VSS.n11933 3.4105
R13936 VSS.n11934 VSS.n11906 3.4105
R13937 VSS.n11955 VSS.n11954 3.4105
R13938 VSS.n11932 VSS.n11931 3.4105
R13939 VSS.n11931 VSS.n11930 3.4105
R13940 VSS.n12848 VSS.n12299 3.4105
R13941 VSS.n12854 VSS.n12299 3.4105
R13942 VSS.n12850 VSS.n12849 3.4105
R13943 VSS.n12874 VSS.n12873 3.4105
R13944 VSS.n12873 VSS.n12872 3.4105
R13945 VSS.n12831 VSS.n12829 3.4105
R13946 VSS.n12831 VSS.n12830 3.4105
R13947 VSS.n12847 VSS.n12846 3.4105
R13948 VSS.n12846 VSS.n12845 3.4105
R13949 VSS.n12809 VSS.n12808 3.4105
R13950 VSS.n12808 VSS.n12807 3.4105
R13951 VSS.n12312 VSS.n12311 3.4105
R13952 VSS.n12828 VSS.n12827 3.4105
R13953 VSS.n12827 VSS.n12826 3.4105
R13954 VSS.n12792 VSS.n12791 3.4105
R13955 VSS.n12811 VSS.n12810 3.4105
R13956 VSS.n12776 VSS.n12775 3.4105
R13957 VSS.n12775 VSS.n12774 3.4105
R13958 VSS.n12777 VSS.n12330 3.4105
R13959 VSS.n12780 VSS.n12325 3.4105
R13960 VSS.n12749 VSS.n12748 3.4105
R13961 VSS.n12749 VSS.n12348 3.4105
R13962 VSS.n12344 VSS.n12331 3.4105
R13963 VSS.n12756 VSS.n12344 3.4105
R13964 VSS.n12695 VSS.n12694 3.4105
R13965 VSS.n12695 VSS.n12358 3.4105
R13966 VSS.n12672 VSS.n12671 3.4105
R13967 VSS.n12693 VSS.n12692 3.4105
R13968 VSS.n12692 VSS.n12691 3.4105
R13969 VSS.n12662 VSS.n12388 3.4105
R13970 VSS.n12388 VSS.n12387 3.4105
R13971 VSS.n12664 VSS.n12663 3.4105
R13972 VSS.n12670 VSS.n12669 3.4105
R13973 VSS.n12669 VSS.n12668 3.4105
R13974 VSS.n12645 VSS.n12644 3.4105
R13975 VSS.n12645 VSS.n12402 3.4105
R13976 VSS.n12641 VSS.n12390 3.4105
R13977 VSS.n12661 VSS.n12660 3.4105
R13978 VSS.n12660 VSS.n12659 3.4105
R13979 VSS.n12624 VSS.n12623 3.4105
R13980 VSS.n12624 VSS.n12418 3.4105
R13981 VSS.n12640 VSS.n12639 3.4105
R13982 VSS.n12622 VSS.n12621 3.4105
R13983 VSS.n12621 VSS.n12620 3.4105
R13984 VSS.n12736 VSS.n12355 3.4105
R13985 VSS.n12710 VSS.n12355 3.4105
R13986 VSS.n12352 VSS.n12351 3.4105
R13987 VSS.n12746 VSS.n12745 3.4105
R13988 VSS.n12745 VSS.n12744 3.4105
R13989 VSS.n12588 VSS.n12587 3.4105
R13990 VSS.n12588 VSS.n12433 3.4105
R13991 VSS.n12581 VSS.n12580 3.4105
R13992 VSS.n12586 VSS.n12585 3.4105
R13993 VSS.n12585 VSS.n12584 3.4105
R13994 VSS.n12561 VSS.n12560 3.4105
R13995 VSS.n12561 VSS.n12473 3.4105
R13996 VSS.n12559 VSS.n12558 3.4105
R13997 VSS.n12579 VSS.n12578 3.4105
R13998 VSS.n12578 VSS.n12577 3.4105
R13999 VSS.n12548 VSS.n12479 3.4105
R14000 VSS.n12479 VSS.n12478 3.4105
R14001 VSS.n12477 VSS.n12476 3.4105
R14002 VSS.n12556 VSS.n12555 3.4105
R14003 VSS.n12555 VSS.n12471 3.4105
R14004 VSS.n12526 VSS.n12525 3.4105
R14005 VSS.n12526 VSS.n12498 3.4105
R14006 VSS.n12547 VSS.n12546 3.4105
R14007 VSS.n12524 VSS.n12523 3.4105
R14008 VSS.n12523 VSS.n12522 3.4105
R14009 VSS.n13440 VSS.n12891 3.4105
R14010 VSS.n13446 VSS.n12891 3.4105
R14011 VSS.n13442 VSS.n13441 3.4105
R14012 VSS.n13466 VSS.n13465 3.4105
R14013 VSS.n13465 VSS.n13464 3.4105
R14014 VSS.n13423 VSS.n13421 3.4105
R14015 VSS.n13423 VSS.n13422 3.4105
R14016 VSS.n13439 VSS.n13438 3.4105
R14017 VSS.n13438 VSS.n13437 3.4105
R14018 VSS.n13401 VSS.n13400 3.4105
R14019 VSS.n13400 VSS.n13399 3.4105
R14020 VSS.n12904 VSS.n12903 3.4105
R14021 VSS.n13420 VSS.n13419 3.4105
R14022 VSS.n13419 VSS.n13418 3.4105
R14023 VSS.n13384 VSS.n13383 3.4105
R14024 VSS.n13403 VSS.n13402 3.4105
R14025 VSS.n13368 VSS.n13367 3.4105
R14026 VSS.n13367 VSS.n13366 3.4105
R14027 VSS.n13369 VSS.n12922 3.4105
R14028 VSS.n13372 VSS.n12917 3.4105
R14029 VSS.n13341 VSS.n13340 3.4105
R14030 VSS.n13341 VSS.n12940 3.4105
R14031 VSS.n12936 VSS.n12923 3.4105
R14032 VSS.n13348 VSS.n12936 3.4105
R14033 VSS.n13287 VSS.n13286 3.4105
R14034 VSS.n13287 VSS.n12950 3.4105
R14035 VSS.n13264 VSS.n13263 3.4105
R14036 VSS.n13285 VSS.n13284 3.4105
R14037 VSS.n13284 VSS.n13283 3.4105
R14038 VSS.n13254 VSS.n12980 3.4105
R14039 VSS.n12980 VSS.n12979 3.4105
R14040 VSS.n13256 VSS.n13255 3.4105
R14041 VSS.n13262 VSS.n13261 3.4105
R14042 VSS.n13261 VSS.n13260 3.4105
R14043 VSS.n13237 VSS.n13236 3.4105
R14044 VSS.n13237 VSS.n12994 3.4105
R14045 VSS.n13233 VSS.n12982 3.4105
R14046 VSS.n13253 VSS.n13252 3.4105
R14047 VSS.n13252 VSS.n13251 3.4105
R14048 VSS.n13216 VSS.n13215 3.4105
R14049 VSS.n13216 VSS.n13010 3.4105
R14050 VSS.n13232 VSS.n13231 3.4105
R14051 VSS.n13214 VSS.n13213 3.4105
R14052 VSS.n13213 VSS.n13212 3.4105
R14053 VSS.n13328 VSS.n12947 3.4105
R14054 VSS.n13302 VSS.n12947 3.4105
R14055 VSS.n12944 VSS.n12943 3.4105
R14056 VSS.n13338 VSS.n13337 3.4105
R14057 VSS.n13337 VSS.n13336 3.4105
R14058 VSS.n13180 VSS.n13179 3.4105
R14059 VSS.n13180 VSS.n13025 3.4105
R14060 VSS.n13173 VSS.n13172 3.4105
R14061 VSS.n13178 VSS.n13177 3.4105
R14062 VSS.n13177 VSS.n13176 3.4105
R14063 VSS.n13153 VSS.n13152 3.4105
R14064 VSS.n13153 VSS.n13065 3.4105
R14065 VSS.n13151 VSS.n13150 3.4105
R14066 VSS.n13171 VSS.n13170 3.4105
R14067 VSS.n13170 VSS.n13169 3.4105
R14068 VSS.n13140 VSS.n13071 3.4105
R14069 VSS.n13071 VSS.n13070 3.4105
R14070 VSS.n13069 VSS.n13068 3.4105
R14071 VSS.n13148 VSS.n13147 3.4105
R14072 VSS.n13147 VSS.n13063 3.4105
R14073 VSS.n13118 VSS.n13117 3.4105
R14074 VSS.n13118 VSS.n13090 3.4105
R14075 VSS.n13139 VSS.n13138 3.4105
R14076 VSS.n13116 VSS.n13115 3.4105
R14077 VSS.n13115 VSS.n13114 3.4105
R14078 VSS.n14032 VSS.n13483 3.4105
R14079 VSS.n14038 VSS.n13483 3.4105
R14080 VSS.n14034 VSS.n14033 3.4105
R14081 VSS.n14058 VSS.n14057 3.4105
R14082 VSS.n14057 VSS.n14056 3.4105
R14083 VSS.n14015 VSS.n14013 3.4105
R14084 VSS.n14015 VSS.n14014 3.4105
R14085 VSS.n14031 VSS.n14030 3.4105
R14086 VSS.n14030 VSS.n14029 3.4105
R14087 VSS.n13993 VSS.n13992 3.4105
R14088 VSS.n13992 VSS.n13991 3.4105
R14089 VSS.n13496 VSS.n13495 3.4105
R14090 VSS.n14012 VSS.n14011 3.4105
R14091 VSS.n14011 VSS.n14010 3.4105
R14092 VSS.n13976 VSS.n13975 3.4105
R14093 VSS.n13995 VSS.n13994 3.4105
R14094 VSS.n13960 VSS.n13959 3.4105
R14095 VSS.n13959 VSS.n13958 3.4105
R14096 VSS.n13961 VSS.n13514 3.4105
R14097 VSS.n13964 VSS.n13509 3.4105
R14098 VSS.n13933 VSS.n13932 3.4105
R14099 VSS.n13933 VSS.n13532 3.4105
R14100 VSS.n13528 VSS.n13515 3.4105
R14101 VSS.n13940 VSS.n13528 3.4105
R14102 VSS.n13879 VSS.n13878 3.4105
R14103 VSS.n13879 VSS.n13542 3.4105
R14104 VSS.n13856 VSS.n13855 3.4105
R14105 VSS.n13877 VSS.n13876 3.4105
R14106 VSS.n13876 VSS.n13875 3.4105
R14107 VSS.n13846 VSS.n13572 3.4105
R14108 VSS.n13572 VSS.n13571 3.4105
R14109 VSS.n13848 VSS.n13847 3.4105
R14110 VSS.n13854 VSS.n13853 3.4105
R14111 VSS.n13853 VSS.n13852 3.4105
R14112 VSS.n13829 VSS.n13828 3.4105
R14113 VSS.n13829 VSS.n13586 3.4105
R14114 VSS.n13825 VSS.n13574 3.4105
R14115 VSS.n13845 VSS.n13844 3.4105
R14116 VSS.n13844 VSS.n13843 3.4105
R14117 VSS.n13808 VSS.n13807 3.4105
R14118 VSS.n13808 VSS.n13602 3.4105
R14119 VSS.n13824 VSS.n13823 3.4105
R14120 VSS.n13806 VSS.n13805 3.4105
R14121 VSS.n13805 VSS.n13804 3.4105
R14122 VSS.n13920 VSS.n13539 3.4105
R14123 VSS.n13894 VSS.n13539 3.4105
R14124 VSS.n13536 VSS.n13535 3.4105
R14125 VSS.n13930 VSS.n13929 3.4105
R14126 VSS.n13929 VSS.n13928 3.4105
R14127 VSS.n13772 VSS.n13771 3.4105
R14128 VSS.n13772 VSS.n13617 3.4105
R14129 VSS.n13765 VSS.n13764 3.4105
R14130 VSS.n13770 VSS.n13769 3.4105
R14131 VSS.n13769 VSS.n13768 3.4105
R14132 VSS.n13745 VSS.n13744 3.4105
R14133 VSS.n13745 VSS.n13657 3.4105
R14134 VSS.n13743 VSS.n13742 3.4105
R14135 VSS.n13763 VSS.n13762 3.4105
R14136 VSS.n13762 VSS.n13761 3.4105
R14137 VSS.n13732 VSS.n13663 3.4105
R14138 VSS.n13663 VSS.n13662 3.4105
R14139 VSS.n13661 VSS.n13660 3.4105
R14140 VSS.n13740 VSS.n13739 3.4105
R14141 VSS.n13739 VSS.n13655 3.4105
R14142 VSS.n13710 VSS.n13709 3.4105
R14143 VSS.n13710 VSS.n13682 3.4105
R14144 VSS.n13731 VSS.n13730 3.4105
R14145 VSS.n13708 VSS.n13707 3.4105
R14146 VSS.n13707 VSS.n13706 3.4105
R14147 VSS.n14624 VSS.n14075 3.4105
R14148 VSS.n14630 VSS.n14075 3.4105
R14149 VSS.n14626 VSS.n14625 3.4105
R14150 VSS.n14650 VSS.n14649 3.4105
R14151 VSS.n14649 VSS.n14648 3.4105
R14152 VSS.n14607 VSS.n14605 3.4105
R14153 VSS.n14607 VSS.n14606 3.4105
R14154 VSS.n14623 VSS.n14622 3.4105
R14155 VSS.n14622 VSS.n14621 3.4105
R14156 VSS.n14585 VSS.n14584 3.4105
R14157 VSS.n14584 VSS.n14583 3.4105
R14158 VSS.n14088 VSS.n14087 3.4105
R14159 VSS.n14604 VSS.n14603 3.4105
R14160 VSS.n14603 VSS.n14602 3.4105
R14161 VSS.n14568 VSS.n14567 3.4105
R14162 VSS.n14587 VSS.n14586 3.4105
R14163 VSS.n14552 VSS.n14551 3.4105
R14164 VSS.n14551 VSS.n14550 3.4105
R14165 VSS.n14553 VSS.n14106 3.4105
R14166 VSS.n14556 VSS.n14101 3.4105
R14167 VSS.n14525 VSS.n14524 3.4105
R14168 VSS.n14525 VSS.n14124 3.4105
R14169 VSS.n14120 VSS.n14107 3.4105
R14170 VSS.n14532 VSS.n14120 3.4105
R14171 VSS.n14471 VSS.n14470 3.4105
R14172 VSS.n14471 VSS.n14134 3.4105
R14173 VSS.n14448 VSS.n14447 3.4105
R14174 VSS.n14469 VSS.n14468 3.4105
R14175 VSS.n14468 VSS.n14467 3.4105
R14176 VSS.n14438 VSS.n14164 3.4105
R14177 VSS.n14164 VSS.n14163 3.4105
R14178 VSS.n14440 VSS.n14439 3.4105
R14179 VSS.n14446 VSS.n14445 3.4105
R14180 VSS.n14445 VSS.n14444 3.4105
R14181 VSS.n14421 VSS.n14420 3.4105
R14182 VSS.n14421 VSS.n14178 3.4105
R14183 VSS.n14417 VSS.n14166 3.4105
R14184 VSS.n14437 VSS.n14436 3.4105
R14185 VSS.n14436 VSS.n14435 3.4105
R14186 VSS.n14400 VSS.n14399 3.4105
R14187 VSS.n14400 VSS.n14194 3.4105
R14188 VSS.n14416 VSS.n14415 3.4105
R14189 VSS.n14398 VSS.n14397 3.4105
R14190 VSS.n14397 VSS.n14396 3.4105
R14191 VSS.n14512 VSS.n14131 3.4105
R14192 VSS.n14486 VSS.n14131 3.4105
R14193 VSS.n14128 VSS.n14127 3.4105
R14194 VSS.n14522 VSS.n14521 3.4105
R14195 VSS.n14521 VSS.n14520 3.4105
R14196 VSS.n14364 VSS.n14363 3.4105
R14197 VSS.n14364 VSS.n14209 3.4105
R14198 VSS.n14357 VSS.n14356 3.4105
R14199 VSS.n14362 VSS.n14361 3.4105
R14200 VSS.n14361 VSS.n14360 3.4105
R14201 VSS.n14337 VSS.n14336 3.4105
R14202 VSS.n14337 VSS.n14249 3.4105
R14203 VSS.n14335 VSS.n14334 3.4105
R14204 VSS.n14355 VSS.n14354 3.4105
R14205 VSS.n14354 VSS.n14353 3.4105
R14206 VSS.n14324 VSS.n14255 3.4105
R14207 VSS.n14255 VSS.n14254 3.4105
R14208 VSS.n14253 VSS.n14252 3.4105
R14209 VSS.n14332 VSS.n14331 3.4105
R14210 VSS.n14331 VSS.n14247 3.4105
R14211 VSS.n14302 VSS.n14301 3.4105
R14212 VSS.n14302 VSS.n14274 3.4105
R14213 VSS.n14323 VSS.n14322 3.4105
R14214 VSS.n14300 VSS.n14299 3.4105
R14215 VSS.n14299 VSS.n14298 3.4105
R14216 VSS.n15216 VSS.n14667 3.4105
R14217 VSS.n15222 VSS.n14667 3.4105
R14218 VSS.n15218 VSS.n15217 3.4105
R14219 VSS.n15242 VSS.n15241 3.4105
R14220 VSS.n15241 VSS.n15240 3.4105
R14221 VSS.n15199 VSS.n15197 3.4105
R14222 VSS.n15199 VSS.n15198 3.4105
R14223 VSS.n15215 VSS.n15214 3.4105
R14224 VSS.n15214 VSS.n15213 3.4105
R14225 VSS.n15177 VSS.n15176 3.4105
R14226 VSS.n15176 VSS.n15175 3.4105
R14227 VSS.n14680 VSS.n14679 3.4105
R14228 VSS.n15196 VSS.n15195 3.4105
R14229 VSS.n15195 VSS.n15194 3.4105
R14230 VSS.n15160 VSS.n15159 3.4105
R14231 VSS.n15179 VSS.n15178 3.4105
R14232 VSS.n15144 VSS.n15143 3.4105
R14233 VSS.n15143 VSS.n15142 3.4105
R14234 VSS.n15145 VSS.n14698 3.4105
R14235 VSS.n15148 VSS.n14693 3.4105
R14236 VSS.n15117 VSS.n15116 3.4105
R14237 VSS.n15117 VSS.n14716 3.4105
R14238 VSS.n14712 VSS.n14699 3.4105
R14239 VSS.n15124 VSS.n14712 3.4105
R14240 VSS.n15063 VSS.n15062 3.4105
R14241 VSS.n15063 VSS.n14726 3.4105
R14242 VSS.n15040 VSS.n15039 3.4105
R14243 VSS.n15061 VSS.n15060 3.4105
R14244 VSS.n15060 VSS.n15059 3.4105
R14245 VSS.n15030 VSS.n14756 3.4105
R14246 VSS.n14756 VSS.n14755 3.4105
R14247 VSS.n15032 VSS.n15031 3.4105
R14248 VSS.n15038 VSS.n15037 3.4105
R14249 VSS.n15037 VSS.n15036 3.4105
R14250 VSS.n15013 VSS.n15012 3.4105
R14251 VSS.n15013 VSS.n14770 3.4105
R14252 VSS.n15009 VSS.n14758 3.4105
R14253 VSS.n15029 VSS.n15028 3.4105
R14254 VSS.n15028 VSS.n15027 3.4105
R14255 VSS.n14992 VSS.n14991 3.4105
R14256 VSS.n14992 VSS.n14786 3.4105
R14257 VSS.n15008 VSS.n15007 3.4105
R14258 VSS.n14990 VSS.n14989 3.4105
R14259 VSS.n14989 VSS.n14988 3.4105
R14260 VSS.n15104 VSS.n14723 3.4105
R14261 VSS.n15078 VSS.n14723 3.4105
R14262 VSS.n14720 VSS.n14719 3.4105
R14263 VSS.n15114 VSS.n15113 3.4105
R14264 VSS.n15113 VSS.n15112 3.4105
R14265 VSS.n14956 VSS.n14955 3.4105
R14266 VSS.n14956 VSS.n14801 3.4105
R14267 VSS.n14949 VSS.n14948 3.4105
R14268 VSS.n14954 VSS.n14953 3.4105
R14269 VSS.n14953 VSS.n14952 3.4105
R14270 VSS.n14929 VSS.n14928 3.4105
R14271 VSS.n14929 VSS.n14841 3.4105
R14272 VSS.n14927 VSS.n14926 3.4105
R14273 VSS.n14947 VSS.n14946 3.4105
R14274 VSS.n14946 VSS.n14945 3.4105
R14275 VSS.n14916 VSS.n14847 3.4105
R14276 VSS.n14847 VSS.n14846 3.4105
R14277 VSS.n14845 VSS.n14844 3.4105
R14278 VSS.n14924 VSS.n14923 3.4105
R14279 VSS.n14923 VSS.n14839 3.4105
R14280 VSS.n14894 VSS.n14893 3.4105
R14281 VSS.n14894 VSS.n14866 3.4105
R14282 VSS.n14915 VSS.n14914 3.4105
R14283 VSS.n14892 VSS.n14891 3.4105
R14284 VSS.n14891 VSS.n14890 3.4105
R14285 VSS.n15808 VSS.n15259 3.4105
R14286 VSS.n15814 VSS.n15259 3.4105
R14287 VSS.n15810 VSS.n15809 3.4105
R14288 VSS.n15834 VSS.n15833 3.4105
R14289 VSS.n15833 VSS.n15832 3.4105
R14290 VSS.n15791 VSS.n15789 3.4105
R14291 VSS.n15791 VSS.n15790 3.4105
R14292 VSS.n15807 VSS.n15806 3.4105
R14293 VSS.n15806 VSS.n15805 3.4105
R14294 VSS.n15769 VSS.n15768 3.4105
R14295 VSS.n15768 VSS.n15767 3.4105
R14296 VSS.n15272 VSS.n15271 3.4105
R14297 VSS.n15788 VSS.n15787 3.4105
R14298 VSS.n15787 VSS.n15786 3.4105
R14299 VSS.n15752 VSS.n15751 3.4105
R14300 VSS.n15771 VSS.n15770 3.4105
R14301 VSS.n15736 VSS.n15735 3.4105
R14302 VSS.n15735 VSS.n15734 3.4105
R14303 VSS.n15737 VSS.n15290 3.4105
R14304 VSS.n15740 VSS.n15285 3.4105
R14305 VSS.n15709 VSS.n15708 3.4105
R14306 VSS.n15709 VSS.n15308 3.4105
R14307 VSS.n15304 VSS.n15291 3.4105
R14308 VSS.n15716 VSS.n15304 3.4105
R14309 VSS.n15655 VSS.n15654 3.4105
R14310 VSS.n15655 VSS.n15318 3.4105
R14311 VSS.n15632 VSS.n15631 3.4105
R14312 VSS.n15653 VSS.n15652 3.4105
R14313 VSS.n15652 VSS.n15651 3.4105
R14314 VSS.n15622 VSS.n15348 3.4105
R14315 VSS.n15348 VSS.n15347 3.4105
R14316 VSS.n15624 VSS.n15623 3.4105
R14317 VSS.n15630 VSS.n15629 3.4105
R14318 VSS.n15629 VSS.n15628 3.4105
R14319 VSS.n15605 VSS.n15604 3.4105
R14320 VSS.n15605 VSS.n15362 3.4105
R14321 VSS.n15601 VSS.n15350 3.4105
R14322 VSS.n15621 VSS.n15620 3.4105
R14323 VSS.n15620 VSS.n15619 3.4105
R14324 VSS.n15584 VSS.n15583 3.4105
R14325 VSS.n15584 VSS.n15378 3.4105
R14326 VSS.n15600 VSS.n15599 3.4105
R14327 VSS.n15582 VSS.n15581 3.4105
R14328 VSS.n15581 VSS.n15580 3.4105
R14329 VSS.n15696 VSS.n15315 3.4105
R14330 VSS.n15670 VSS.n15315 3.4105
R14331 VSS.n15312 VSS.n15311 3.4105
R14332 VSS.n15706 VSS.n15705 3.4105
R14333 VSS.n15705 VSS.n15704 3.4105
R14334 VSS.n15548 VSS.n15547 3.4105
R14335 VSS.n15548 VSS.n15393 3.4105
R14336 VSS.n15541 VSS.n15540 3.4105
R14337 VSS.n15546 VSS.n15545 3.4105
R14338 VSS.n15545 VSS.n15544 3.4105
R14339 VSS.n15521 VSS.n15520 3.4105
R14340 VSS.n15521 VSS.n15433 3.4105
R14341 VSS.n15519 VSS.n15518 3.4105
R14342 VSS.n15539 VSS.n15538 3.4105
R14343 VSS.n15538 VSS.n15537 3.4105
R14344 VSS.n15508 VSS.n15439 3.4105
R14345 VSS.n15439 VSS.n15438 3.4105
R14346 VSS.n15437 VSS.n15436 3.4105
R14347 VSS.n15516 VSS.n15515 3.4105
R14348 VSS.n15515 VSS.n15431 3.4105
R14349 VSS.n15486 VSS.n15485 3.4105
R14350 VSS.n15486 VSS.n15458 3.4105
R14351 VSS.n15507 VSS.n15506 3.4105
R14352 VSS.n15484 VSS.n15483 3.4105
R14353 VSS.n15483 VSS.n15482 3.4105
R14354 VSS.n6951 VSS.n6905 3.4105
R14355 VSS.n6951 VSS.n6950 3.4105
R14356 VSS.n6954 VSS.n6953 3.4105
R14357 VSS.n15840 VSS.n15839 3.4105
R14358 VSS.n15841 VSS.n15840 3.4105
R14359 VSS.n15858 VSS.n15857 3.4105
R14360 VSS.n15859 VSS.n15858 3.4105
R14361 VSS.n15855 VSS.n15854 3.4105
R14362 VSS.n15854 VSS.n15853 3.4105
R14363 VSS.n15873 VSS.n15872 3.4105
R14364 VSS.n15872 VSS.n15871 3.4105
R14365 VSS.n6903 VSS.n6902 3.4105
R14366 VSS.n6904 VSS.n6896 3.4105
R14367 VSS.n6896 VSS.n6892 3.4105
R14368 VSS.n6886 VSS.n6885 3.4105
R14369 VSS.n15875 VSS.n15874 3.4105
R14370 VSS.n15890 VSS.n6854 3.4105
R14371 VSS.n15890 VSS.n15889 3.4105
R14372 VSS.n6871 VSS.n6847 3.4105
R14373 VSS.n6874 VSS.n6867 3.4105
R14374 VSS.n15906 VSS.n6837 3.4105
R14375 VSS.n15906 VSS.n15905 3.4105
R14376 VSS.n6853 VSS.n6852 3.4105
R14377 VSS.n6852 VSS.n6851 3.4105
R14378 VSS.n15929 VSS.n15928 3.4105
R14379 VSS.n15928 VSS.n15927 3.4105
R14380 VSS.n15936 VSS.n15935 3.4105
R14381 VSS.n15931 VSS.n15930 3.4105
R14382 VSS.n15932 VSS.n15931 3.4105
R14383 VSS.n15944 VSS.n15943 3.4105
R14384 VSS.n15943 VSS.n15942 3.4105
R14385 VSS.n6699 VSS.n6695 3.4105
R14386 VSS.n15938 VSS.n15937 3.4105
R14387 VSS.n15938 VSS.n6698 3.4105
R14388 VSS.n15952 VSS.n15951 3.4105
R14389 VSS.n15951 VSS.n15950 3.4105
R14390 VSS.n6694 VSS.n6692 3.4105
R14391 VSS.n15946 VSS.n15945 3.4105
R14392 VSS.n15946 VSS.n6690 3.4105
R14393 VSS.n15959 VSS.n15958 3.4105
R14394 VSS.n15958 VSS.n15957 3.4105
R14395 VSS.n15954 VSS.n15953 3.4105
R14396 VSS.n15960 VSS.n6679 3.4105
R14397 VSS.n6679 VSS.n6498 3.4105
R14398 VSS.n6828 VSS.n6826 3.4105
R14399 VSS.n6826 VSS.n6825 3.4105
R14400 VSS.n6820 VSS.n6819 3.4105
R14401 VSS.n6836 VSS.n6835 3.4105
R14402 VSS.n6835 VSS.n6834 3.4105
R14403 VSS.n6656 VSS.n6655 3.4105
R14404 VSS.n6656 VSS.n6501 3.4105
R14405 VSS.n6649 VSS.n6648 3.4105
R14406 VSS.n6654 VSS.n6653 3.4105
R14407 VSS.n6653 VSS.n6652 3.4105
R14408 VSS.n6629 VSS.n6628 3.4105
R14409 VSS.n6629 VSS.n6541 3.4105
R14410 VSS.n6627 VSS.n6626 3.4105
R14411 VSS.n6647 VSS.n6646 3.4105
R14412 VSS.n6646 VSS.n6645 3.4105
R14413 VSS.n6616 VSS.n6547 3.4105
R14414 VSS.n6547 VSS.n6546 3.4105
R14415 VSS.n6545 VSS.n6544 3.4105
R14416 VSS.n6624 VSS.n6623 3.4105
R14417 VSS.n6623 VSS.n6539 3.4105
R14418 VSS.n6594 VSS.n6593 3.4105
R14419 VSS.n6594 VSS.n6566 3.4105
R14420 VSS.n6615 VSS.n6614 3.4105
R14421 VSS.n6592 VSS.n6591 3.4105
R14422 VSS.n6591 VSS.n6590 3.4105
R14423 VSS.n7520 VSS.n6970 3.4105
R14424 VSS.n7526 VSS.n6970 3.4105
R14425 VSS.n7522 VSS.n7521 3.4105
R14426 VSS.n7546 VSS.n7545 3.4105
R14427 VSS.n7545 VSS.n7544 3.4105
R14428 VSS.n7503 VSS.n7501 3.4105
R14429 VSS.n7503 VSS.n7502 3.4105
R14430 VSS.n7519 VSS.n7518 3.4105
R14431 VSS.n7518 VSS.n7517 3.4105
R14432 VSS.n7481 VSS.n7480 3.4105
R14433 VSS.n7480 VSS.n7479 3.4105
R14434 VSS.n6983 VSS.n6982 3.4105
R14435 VSS.n7500 VSS.n7499 3.4105
R14436 VSS.n7499 VSS.n7498 3.4105
R14437 VSS.n7464 VSS.n7463 3.4105
R14438 VSS.n7483 VSS.n7482 3.4105
R14439 VSS.n7448 VSS.n7447 3.4105
R14440 VSS.n7447 VSS.n7446 3.4105
R14441 VSS.n7449 VSS.n7001 3.4105
R14442 VSS.n7452 VSS.n6996 3.4105
R14443 VSS.n7421 VSS.n7420 3.4105
R14444 VSS.n7421 VSS.n7019 3.4105
R14445 VSS.n7015 VSS.n7002 3.4105
R14446 VSS.n7428 VSS.n7015 3.4105
R14447 VSS.n7367 VSS.n7366 3.4105
R14448 VSS.n7367 VSS.n7029 3.4105
R14449 VSS.n7344 VSS.n7343 3.4105
R14450 VSS.n7365 VSS.n7364 3.4105
R14451 VSS.n7364 VSS.n7363 3.4105
R14452 VSS.n7334 VSS.n7059 3.4105
R14453 VSS.n7059 VSS.n7058 3.4105
R14454 VSS.n7336 VSS.n7335 3.4105
R14455 VSS.n7342 VSS.n7341 3.4105
R14456 VSS.n7341 VSS.n7340 3.4105
R14457 VSS.n7317 VSS.n7316 3.4105
R14458 VSS.n7317 VSS.n7073 3.4105
R14459 VSS.n7313 VSS.n7061 3.4105
R14460 VSS.n7333 VSS.n7332 3.4105
R14461 VSS.n7332 VSS.n7331 3.4105
R14462 VSS.n7296 VSS.n7295 3.4105
R14463 VSS.n7296 VSS.n7089 3.4105
R14464 VSS.n7312 VSS.n7311 3.4105
R14465 VSS.n7294 VSS.n7293 3.4105
R14466 VSS.n7293 VSS.n7292 3.4105
R14467 VSS.n7408 VSS.n7026 3.4105
R14468 VSS.n7382 VSS.n7026 3.4105
R14469 VSS.n7023 VSS.n7022 3.4105
R14470 VSS.n7418 VSS.n7417 3.4105
R14471 VSS.n7417 VSS.n7416 3.4105
R14472 VSS.n7263 VSS.n7262 3.4105
R14473 VSS.n7263 VSS.n7104 3.4105
R14474 VSS.n7239 VSS.n7238 3.4105
R14475 VSS.n7261 VSS.n7260 3.4105
R14476 VSS.n7260 VSS.n7259 3.4105
R14477 VSS.n7229 VSS.n7134 3.4105
R14478 VSS.n7134 VSS.n7133 3.4105
R14479 VSS.n7231 VSS.n7230 3.4105
R14480 VSS.n7237 VSS.n7236 3.4105
R14481 VSS.n7236 VSS.n7235 3.4105
R14482 VSS.n7212 VSS.n7211 3.4105
R14483 VSS.n7212 VSS.n7150 3.4105
R14484 VSS.n7208 VSS.n7136 3.4105
R14485 VSS.n7228 VSS.n7227 3.4105
R14486 VSS.n7227 VSS.n7226 3.4105
R14487 VSS.n7191 VSS.n7190 3.4105
R14488 VSS.n7191 VSS.n7164 3.4105
R14489 VSS.n7207 VSS.n7206 3.4105
R14490 VSS.n7189 VSS.n7188 3.4105
R14491 VSS.n7188 VSS.n7187 3.4105
R14492 VSS.n18832 VSS.n68 3.4105
R14493 VSS.n18838 VSS.n68 3.4105
R14494 VSS.n18834 VSS.n18833 3.4105
R14495 VSS.n18858 VSS.n18857 3.4105
R14496 VSS.n18857 VSS.n18856 3.4105
R14497 VSS.n18815 VSS.n18813 3.4105
R14498 VSS.n18815 VSS.n18814 3.4105
R14499 VSS.n18831 VSS.n18830 3.4105
R14500 VSS.n18830 VSS.n18829 3.4105
R14501 VSS.n18793 VSS.n18792 3.4105
R14502 VSS.n18792 VSS.n18791 3.4105
R14503 VSS.n81 VSS.n80 3.4105
R14504 VSS.n18812 VSS.n18811 3.4105
R14505 VSS.n18811 VSS.n18810 3.4105
R14506 VSS.n18776 VSS.n18775 3.4105
R14507 VSS.n18795 VSS.n18794 3.4105
R14508 VSS.n18760 VSS.n18759 3.4105
R14509 VSS.n18759 VSS.n18758 3.4105
R14510 VSS.n18761 VSS.n99 3.4105
R14511 VSS.n18764 VSS.n94 3.4105
R14512 VSS.n18733 VSS.n18732 3.4105
R14513 VSS.n18733 VSS.n117 3.4105
R14514 VSS.n113 VSS.n100 3.4105
R14515 VSS.n18740 VSS.n113 3.4105
R14516 VSS.n18679 VSS.n18678 3.4105
R14517 VSS.n18679 VSS.n127 3.4105
R14518 VSS.n18656 VSS.n18655 3.4105
R14519 VSS.n18677 VSS.n18676 3.4105
R14520 VSS.n18676 VSS.n18675 3.4105
R14521 VSS.n18646 VSS.n157 3.4105
R14522 VSS.n157 VSS.n156 3.4105
R14523 VSS.n18648 VSS.n18647 3.4105
R14524 VSS.n18654 VSS.n18653 3.4105
R14525 VSS.n18653 VSS.n18652 3.4105
R14526 VSS.n18629 VSS.n18628 3.4105
R14527 VSS.n18629 VSS.n171 3.4105
R14528 VSS.n18625 VSS.n159 3.4105
R14529 VSS.n18645 VSS.n18644 3.4105
R14530 VSS.n18644 VSS.n18643 3.4105
R14531 VSS.n18608 VSS.n18607 3.4105
R14532 VSS.n18608 VSS.n187 3.4105
R14533 VSS.n18624 VSS.n18623 3.4105
R14534 VSS.n18606 VSS.n18605 3.4105
R14535 VSS.n18605 VSS.n18604 3.4105
R14536 VSS.n18720 VSS.n124 3.4105
R14537 VSS.n18694 VSS.n124 3.4105
R14538 VSS.n121 VSS.n120 3.4105
R14539 VSS.n18730 VSS.n18729 3.4105
R14540 VSS.n18729 VSS.n18728 3.4105
R14541 VSS.n415 VSS.n414 3.4105
R14542 VSS.n414 VSS.n195 3.4105
R14543 VSS.n422 VSS.n421 3.4105
R14544 VSS.n417 VSS.n416 3.4105
R14545 VSS.n418 VSS.n417 3.4105
R14546 VSS.n430 VSS.n429 3.4105
R14547 VSS.n429 VSS.n428 3.4105
R14548 VSS.n314 VSS.n309 3.4105
R14549 VSS.n424 VSS.n423 3.4105
R14550 VSS.n424 VSS.n313 3.4105
R14551 VSS.n438 VSS.n437 3.4105
R14552 VSS.n437 VSS.n436 3.4105
R14553 VSS.n308 VSS.n306 3.4105
R14554 VSS.n432 VSS.n431 3.4105
R14555 VSS.n432 VSS.n304 3.4105
R14556 VSS.n445 VSS.n444 3.4105
R14557 VSS.n444 VSS.n443 3.4105
R14558 VSS.n440 VSS.n439 3.4105
R14559 VSS.n446 VSS.n293 3.4105
R14560 VSS.n293 VSS.n291 3.4105
R14561 VSS.n734 VSS.n733 3.4105
R14562 VSS.n772 VSS.n771 3.4105
R14563 VSS.n773 VSS.n772 3.4105
R14564 VSS.n769 VSS.n768 3.4105
R14565 VSS.n768 VSS.n767 3.4105
R14566 VSS.n787 VSS.n786 3.4105
R14567 VSS.n786 VSS.n785 3.4105
R14568 VSS.n726 VSS.n725 3.4105
R14569 VSS.n727 VSS.n719 3.4105
R14570 VSS.n719 VSS.n715 3.4105
R14571 VSS.n709 VSS.n708 3.4105
R14572 VSS.n789 VSS.n788 3.4105
R14573 VSS.n804 VSS.n677 3.4105
R14574 VSS.n804 VSS.n803 3.4105
R14575 VSS.n694 VSS.n670 3.4105
R14576 VSS.n697 VSS.n690 3.4105
R14577 VSS.n820 VSS.n660 3.4105
R14578 VSS.n820 VSS.n819 3.4105
R14579 VSS.n676 VSS.n675 3.4105
R14580 VSS.n675 VSS.n674 3.4105
R14581 VSS.n651 VSS.n649 3.4105
R14582 VSS.n649 VSS.n648 3.4105
R14583 VSS.n643 VSS.n642 3.4105
R14584 VSS.n659 VSS.n658 3.4105
R14585 VSS.n658 VSS.n657 3.4105
R14586 VSS.n735 VSS.n728 3.4105
R14587 VSS.n737 VSS.n735 3.4105
R14588 VSS.n843 VSS.n842 3.4105
R14589 VSS.n842 VSS.n841 3.4105
R14590 VSS.n850 VSS.n849 3.4105
R14591 VSS.n845 VSS.n844 3.4105
R14592 VSS.n846 VSS.n845 3.4105
R14593 VSS.n858 VSS.n857 3.4105
R14594 VSS.n857 VSS.n856 3.4105
R14595 VSS.n519 VSS.n515 3.4105
R14596 VSS.n852 VSS.n851 3.4105
R14597 VSS.n852 VSS.n518 3.4105
R14598 VSS.n866 VSS.n865 3.4105
R14599 VSS.n865 VSS.n864 3.4105
R14600 VSS.n514 VSS.n512 3.4105
R14601 VSS.n860 VSS.n859 3.4105
R14602 VSS.n860 VSS.n510 3.4105
R14603 VSS.n873 VSS.n872 3.4105
R14604 VSS.n872 VSS.n871 3.4105
R14605 VSS.n868 VSS.n867 3.4105
R14606 VSS.n875 VSS.n874 3.4105
R14607 VSS.n876 VSS.n875 3.4105
R14608 VSS.n18863 VSS.n18862 3.4105
R14609 VSS.n18864 VSS.n18863 3.4105
R14610 VSS.n980 VSS.n979 3.4105
R14611 VSS.n979 VSS.n978 3.4105
R14612 VSS.n987 VSS.n986 3.4105
R14613 VSS.n982 VSS.n981 3.4105
R14614 VSS.n983 VSS.n982 3.4105
R14615 VSS.n995 VSS.n994 3.4105
R14616 VSS.n994 VSS.n993 3.4105
R14617 VSS.n480 VSS.n475 3.4105
R14618 VSS.n989 VSS.n988 3.4105
R14619 VSS.n989 VSS.n479 3.4105
R14620 VSS.n1003 VSS.n1002 3.4105
R14621 VSS.n1002 VSS.n1001 3.4105
R14622 VSS.n474 VSS.n472 3.4105
R14623 VSS.n997 VSS.n996 3.4105
R14624 VSS.n997 VSS.n470 3.4105
R14625 VSS.n1010 VSS.n1009 3.4105
R14626 VSS.n1009 VSS.n1008 3.4105
R14627 VSS.n1005 VSS.n1004 3.4105
R14628 VSS.n1011 VSS.n459 3.4105
R14629 VSS.n459 VSS.n457 3.4105
R14630 VSS.n1433 VSS.n1387 3.4105
R14631 VSS.n1433 VSS.n1432 3.4105
R14632 VSS.n1436 VSS.n1435 3.4105
R14633 VSS.n17868 VSS.n17867 3.4105
R14634 VSS.n17869 VSS.n17868 3.4105
R14635 VSS.n17886 VSS.n17885 3.4105
R14636 VSS.n17887 VSS.n17886 3.4105
R14637 VSS.n17883 VSS.n17882 3.4105
R14638 VSS.n17882 VSS.n17881 3.4105
R14639 VSS.n17901 VSS.n17900 3.4105
R14640 VSS.n17900 VSS.n17899 3.4105
R14641 VSS.n1385 VSS.n1384 3.4105
R14642 VSS.n1386 VSS.n1378 3.4105
R14643 VSS.n1378 VSS.n1374 3.4105
R14644 VSS.n1368 VSS.n1367 3.4105
R14645 VSS.n17903 VSS.n17902 3.4105
R14646 VSS.n17918 VSS.n1336 3.4105
R14647 VSS.n17918 VSS.n17917 3.4105
R14648 VSS.n1353 VSS.n1329 3.4105
R14649 VSS.n1356 VSS.n1349 3.4105
R14650 VSS.n17934 VSS.n1319 3.4105
R14651 VSS.n17934 VSS.n17933 3.4105
R14652 VSS.n1335 VSS.n1334 3.4105
R14653 VSS.n1334 VSS.n1333 3.4105
R14654 VSS.n17957 VSS.n17956 3.4105
R14655 VSS.n17956 VSS.n17955 3.4105
R14656 VSS.n17964 VSS.n17963 3.4105
R14657 VSS.n17959 VSS.n17958 3.4105
R14658 VSS.n17960 VSS.n17959 3.4105
R14659 VSS.n17972 VSS.n17971 3.4105
R14660 VSS.n17971 VSS.n17970 3.4105
R14661 VSS.n1181 VSS.n1177 3.4105
R14662 VSS.n17966 VSS.n17965 3.4105
R14663 VSS.n17966 VSS.n1180 3.4105
R14664 VSS.n17980 VSS.n17979 3.4105
R14665 VSS.n17979 VSS.n17978 3.4105
R14666 VSS.n1176 VSS.n1174 3.4105
R14667 VSS.n17974 VSS.n17973 3.4105
R14668 VSS.n17974 VSS.n1172 3.4105
R14669 VSS.n17987 VSS.n17986 3.4105
R14670 VSS.n17986 VSS.n17985 3.4105
R14671 VSS.n17982 VSS.n17981 3.4105
R14672 VSS.n17988 VSS.n1161 3.4105
R14673 VSS.n1161 VSS.n1159 3.4105
R14674 VSS.n1310 VSS.n1308 3.4105
R14675 VSS.n1308 VSS.n1307 3.4105
R14676 VSS.n1302 VSS.n1301 3.4105
R14677 VSS.n1318 VSS.n1317 3.4105
R14678 VSS.n1317 VSS.n1316 3.4105
R14679 VSS.n1222 VSS.n1221 3.29193
R14680 VSS.n1242 VSS.n1241 3.29193
R14681 VSS.n1261 VSS.n1206 3.29193
R14682 VSS.n1089 VSS.n1088 3.29193
R14683 VSS.n1107 VSS.n1106 3.29193
R14684 VSS.n1126 VSS.n1072 3.29193
R14685 VSS.n17115 VSS.n17114 3.29193
R14686 VSS.n17258 VSS.n16864 3.29193
R14687 VSS.n17000 VSS.n16990 3.29193
R14688 VSS.n17033 VSS.n17032 3.29193
R14689 VSS.n17071 VSS.n16951 3.29193
R14690 VSS.n17494 VSS.n17483 3.29193
R14691 VSS.n17521 VSS.n17477 3.29193
R14692 VSS.n17456 VSS.n17455 3.29193
R14693 VSS.n17707 VSS.n17706 3.29193
R14694 VSS.n17850 VSS.n17278 3.29193
R14695 VSS.n17414 VSS.n17404 3.29193
R14696 VSS.n17625 VSS.n17624 3.29193
R14697 VSS.n17663 VSS.n17365 3.29193
R14698 VSS.n18239 VSS.n18238 3.29193
R14699 VSS.n18259 VSS.n18258 3.29193
R14700 VSS.n18278 VSS.n18223 3.29193
R14701 VSS.n18322 VSS.n18312 3.29193
R14702 VSS.n18454 VSS.n18435 3.29193
R14703 VSS.n286 VSS.n275 3.29193
R14704 VSS.n18098 VSS.n269 3.29193
R14705 VSS.n248 VSS.n247 3.29193
R14706 VSS.n9464 VSS.n9454 3.29193
R14707 VSS.n9675 VSS.n9674 3.29193
R14708 VSS.n9713 VSS.n9415 3.29193
R14709 VSS.n9757 VSS.n9756 3.29193
R14710 VSS.n9901 VSS.n9329 3.29193
R14711 VSS.n9544 VSS.n9533 3.29193
R14712 VSS.n9571 VSS.n9527 3.29193
R14713 VSS.n9506 VSS.n9505 3.29193
R14714 VSS.n16406 VSS.n16396 3.29193
R14715 VSS.n16618 VSS.n16617 3.29193
R14716 VSS.n16656 VSS.n16357 3.29193
R14717 VSS.n16700 VSS.n16699 3.29193
R14718 VSS.n16844 VSS.n16271 3.29193
R14719 VSS.n16481 VSS.n16471 3.29193
R14720 VSS.n16513 VSS.n16512 3.29193
R14721 VSS.n16551 VSS.n16432 3.29193
R14722 VSS.n1753 VSS.n1568 3.29193
R14723 VSS.n16025 VSS.n16024 3.29193
R14724 VSS.n16063 VSS.n1529 3.29193
R14725 VSS.n16107 VSS.n16106 3.29193
R14726 VSS.n16251 VSS.n1443 3.29193
R14727 VSS.n1646 VSS.n1636 3.29193
R14728 VSS.n1678 VSS.n1677 3.29193
R14729 VSS.n1716 VSS.n1597 3.29193
R14730 VSS.n2004 VSS.n2003 3.29193
R14731 VSS.n2024 VSS.n2023 3.29193
R14732 VSS.n2043 VSS.n1988 3.29193
R14733 VSS.n2086 VSS.n2077 3.29193
R14734 VSS.n2226 VSS.n2225 3.29193
R14735 VSS.n1836 VSS.n1825 3.29193
R14736 VSS.n1863 VSS.n1819 3.29193
R14737 VSS.n1798 VSS.n1797 3.29193
R14738 VSS.n2955 VSS.n2945 3.29193
R14739 VSS.n3166 VSS.n3165 3.29193
R14740 VSS.n3204 VSS.n2906 3.29193
R14741 VSS.n3248 VSS.n3247 3.29193
R14742 VSS.n3392 VSS.n2820 3.29193
R14743 VSS.n3035 VSS.n3024 3.29193
R14744 VSS.n3062 VSS.n3018 3.29193
R14745 VSS.n2997 VSS.n2996 3.29193
R14746 VSS.n3547 VSS.n3537 3.29193
R14747 VSS.n3758 VSS.n3757 3.29193
R14748 VSS.n3796 VSS.n3498 3.29193
R14749 VSS.n3840 VSS.n3839 3.29193
R14750 VSS.n3984 VSS.n3412 3.29193
R14751 VSS.n3627 VSS.n3616 3.29193
R14752 VSS.n3654 VSS.n3610 3.29193
R14753 VSS.n3589 VSS.n3588 3.29193
R14754 VSS.n4139 VSS.n4129 3.29193
R14755 VSS.n4350 VSS.n4349 3.29193
R14756 VSS.n4388 VSS.n4090 3.29193
R14757 VSS.n4432 VSS.n4431 3.29193
R14758 VSS.n4576 VSS.n4004 3.29193
R14759 VSS.n4219 VSS.n4208 3.29193
R14760 VSS.n4246 VSS.n4202 3.29193
R14761 VSS.n4181 VSS.n4180 3.29193
R14762 VSS.n4731 VSS.n4721 3.29193
R14763 VSS.n4942 VSS.n4941 3.29193
R14764 VSS.n4980 VSS.n4682 3.29193
R14765 VSS.n5024 VSS.n5023 3.29193
R14766 VSS.n5168 VSS.n4596 3.29193
R14767 VSS.n4811 VSS.n4800 3.29193
R14768 VSS.n4838 VSS.n4794 3.29193
R14769 VSS.n4773 VSS.n4772 3.29193
R14770 VSS.n2600 VSS.n2599 3.29193
R14771 VSS.n2620 VSS.n2619 3.29193
R14772 VSS.n2639 VSS.n2584 3.29193
R14773 VSS.n2682 VSS.n2673 3.29193
R14774 VSS.n5191 VSS.n5190 3.29193
R14775 VSS.n2432 VSS.n2421 3.29193
R14776 VSS.n2459 VSS.n2415 3.29193
R14777 VSS.n2394 VSS.n2393 3.29193
R14778 VSS.n5561 VSS.n5560 3.29193
R14779 VSS.n5581 VSS.n5580 3.29193
R14780 VSS.n5600 VSS.n5545 3.29193
R14781 VSS.n5643 VSS.n5634 3.29193
R14782 VSS.n5743 VSS.n5 3.29193
R14783 VSS.n5393 VSS.n5382 3.29193
R14784 VSS.n5420 VSS.n5376 3.29193
R14785 VSS.n5355 VSS.n5354 3.29193
R14786 VSS.n6134 VSS.n6133 3.29193
R14787 VSS.n6154 VSS.n6153 3.29193
R14788 VSS.n6173 VSS.n6118 3.29193
R14789 VSS.n6216 VSS.n6207 3.29193
R14790 VSS.n6356 VSS.n6355 3.29193
R14791 VSS.n5966 VSS.n5955 3.29193
R14792 VSS.n5993 VSS.n5949 3.29193
R14793 VSS.n5928 VSS.n5927 3.29193
R14794 VSS.n7688 VSS.n7678 3.29193
R14795 VSS.n7899 VSS.n7898 3.29193
R14796 VSS.n7937 VSS.n7639 3.29193
R14797 VSS.n7981 VSS.n7980 3.29193
R14798 VSS.n8125 VSS.n7553 3.29193
R14799 VSS.n7768 VSS.n7757 3.29193
R14800 VSS.n7795 VSS.n7751 3.29193
R14801 VSS.n7730 VSS.n7729 3.29193
R14802 VSS.n8280 VSS.n8270 3.29193
R14803 VSS.n8491 VSS.n8490 3.29193
R14804 VSS.n8529 VSS.n8231 3.29193
R14805 VSS.n8573 VSS.n8572 3.29193
R14806 VSS.n8717 VSS.n8145 3.29193
R14807 VSS.n8360 VSS.n8349 3.29193
R14808 VSS.n8387 VSS.n8343 3.29193
R14809 VSS.n8322 VSS.n8321 3.29193
R14810 VSS.n8872 VSS.n8862 3.29193
R14811 VSS.n9083 VSS.n9082 3.29193
R14812 VSS.n9121 VSS.n8823 3.29193
R14813 VSS.n9165 VSS.n9164 3.29193
R14814 VSS.n9309 VSS.n8737 3.29193
R14815 VSS.n8952 VSS.n8941 3.29193
R14816 VSS.n8979 VSS.n8935 3.29193
R14817 VSS.n8914 VSS.n8913 3.29193
R14818 VSS.n10056 VSS.n10046 3.29193
R14819 VSS.n10267 VSS.n10266 3.29193
R14820 VSS.n10305 VSS.n10007 3.29193
R14821 VSS.n10349 VSS.n10348 3.29193
R14822 VSS.n10493 VSS.n9921 3.29193
R14823 VSS.n10136 VSS.n10125 3.29193
R14824 VSS.n10163 VSS.n10119 3.29193
R14825 VSS.n10098 VSS.n10097 3.29193
R14826 VSS.n10648 VSS.n10638 3.29193
R14827 VSS.n10859 VSS.n10858 3.29193
R14828 VSS.n10897 VSS.n10599 3.29193
R14829 VSS.n10941 VSS.n10940 3.29193
R14830 VSS.n11085 VSS.n10513 3.29193
R14831 VSS.n10728 VSS.n10717 3.29193
R14832 VSS.n10755 VSS.n10711 3.29193
R14833 VSS.n10690 VSS.n10689 3.29193
R14834 VSS.n11240 VSS.n11230 3.29193
R14835 VSS.n11451 VSS.n11450 3.29193
R14836 VSS.n11489 VSS.n11191 3.29193
R14837 VSS.n11533 VSS.n11532 3.29193
R14838 VSS.n11677 VSS.n11105 3.29193
R14839 VSS.n11320 VSS.n11309 3.29193
R14840 VSS.n11347 VSS.n11303 3.29193
R14841 VSS.n11282 VSS.n11281 3.29193
R14842 VSS.n11832 VSS.n11822 3.29193
R14843 VSS.n12043 VSS.n12042 3.29193
R14844 VSS.n12081 VSS.n11783 3.29193
R14845 VSS.n12125 VSS.n12124 3.29193
R14846 VSS.n12269 VSS.n11697 3.29193
R14847 VSS.n11912 VSS.n11901 3.29193
R14848 VSS.n11939 VSS.n11895 3.29193
R14849 VSS.n11874 VSS.n11873 3.29193
R14850 VSS.n12424 VSS.n12414 3.29193
R14851 VSS.n12635 VSS.n12634 3.29193
R14852 VSS.n12673 VSS.n12375 3.29193
R14853 VSS.n12717 VSS.n12716 3.29193
R14854 VSS.n12861 VSS.n12289 3.29193
R14855 VSS.n12504 VSS.n12493 3.29193
R14856 VSS.n12531 VSS.n12487 3.29193
R14857 VSS.n12466 VSS.n12465 3.29193
R14858 VSS.n13016 VSS.n13006 3.29193
R14859 VSS.n13227 VSS.n13226 3.29193
R14860 VSS.n13265 VSS.n12967 3.29193
R14861 VSS.n13309 VSS.n13308 3.29193
R14862 VSS.n13453 VSS.n12881 3.29193
R14863 VSS.n13096 VSS.n13085 3.29193
R14864 VSS.n13123 VSS.n13079 3.29193
R14865 VSS.n13058 VSS.n13057 3.29193
R14866 VSS.n13608 VSS.n13598 3.29193
R14867 VSS.n13819 VSS.n13818 3.29193
R14868 VSS.n13857 VSS.n13559 3.29193
R14869 VSS.n13901 VSS.n13900 3.29193
R14870 VSS.n14045 VSS.n13473 3.29193
R14871 VSS.n13688 VSS.n13677 3.29193
R14872 VSS.n13715 VSS.n13671 3.29193
R14873 VSS.n13650 VSS.n13649 3.29193
R14874 VSS.n14200 VSS.n14190 3.29193
R14875 VSS.n14411 VSS.n14410 3.29193
R14876 VSS.n14449 VSS.n14151 3.29193
R14877 VSS.n14493 VSS.n14492 3.29193
R14878 VSS.n14637 VSS.n14065 3.29193
R14879 VSS.n14280 VSS.n14269 3.29193
R14880 VSS.n14307 VSS.n14263 3.29193
R14881 VSS.n14242 VSS.n14241 3.29193
R14882 VSS.n14792 VSS.n14782 3.29193
R14883 VSS.n15003 VSS.n15002 3.29193
R14884 VSS.n15041 VSS.n14743 3.29193
R14885 VSS.n15085 VSS.n15084 3.29193
R14886 VSS.n15229 VSS.n14657 3.29193
R14887 VSS.n14872 VSS.n14861 3.29193
R14888 VSS.n14899 VSS.n14855 3.29193
R14889 VSS.n14834 VSS.n14833 3.29193
R14890 VSS.n15384 VSS.n15374 3.29193
R14891 VSS.n15595 VSS.n15594 3.29193
R14892 VSS.n15633 VSS.n15335 3.29193
R14893 VSS.n15677 VSS.n15676 3.29193
R14894 VSS.n15821 VSS.n15249 3.29193
R14895 VSS.n15464 VSS.n15453 3.29193
R14896 VSS.n15491 VSS.n15447 3.29193
R14897 VSS.n15426 VSS.n15425 3.29193
R14898 VSS.n6740 VSS.n6739 3.29193
R14899 VSS.n6760 VSS.n6759 3.29193
R14900 VSS.n6779 VSS.n6724 3.29193
R14901 VSS.n6822 VSS.n6813 3.29193
R14902 VSS.n15844 VSS.n15843 3.29193
R14903 VSS.n6572 VSS.n6561 3.29193
R14904 VSS.n6599 VSS.n6555 3.29193
R14905 VSS.n6534 VSS.n6533 3.29193
R14906 VSS.n7095 VSS.n7085 3.29193
R14907 VSS.n7307 VSS.n7306 3.29193
R14908 VSS.n7345 VSS.n7046 3.29193
R14909 VSS.n7389 VSS.n7388 3.29193
R14910 VSS.n7533 VSS.n6960 3.29193
R14911 VSS.n7170 VSS.n7160 3.29193
R14912 VSS.n7202 VSS.n7201 3.29193
R14913 VSS.n7240 VSS.n7121 3.29193
R14914 VSS.n202 VSS.n183 3.29193
R14915 VSS.n18619 VSS.n18618 3.29193
R14916 VSS.n18657 VSS.n144 3.29193
R14917 VSS.n18701 VSS.n18700 3.29193
R14918 VSS.n18845 VSS.n58 3.29193
R14919 VSS.n357 VSS.n356 3.29193
R14920 VSS.n365 VSS.n364 3.29193
R14921 VSS.n394 VSS.n393 3.29193
R14922 VSS.n565 VSS.n564 3.29193
R14923 VSS.n583 VSS.n582 3.29193
R14924 VSS.n602 VSS.n544 3.29193
R14925 VSS.n645 VSS.n636 3.29193
R14926 VSS.n18867 VSS.n18866 3.29193
R14927 VSS.n908 VSS.n907 3.29193
R14928 VSS.n926 VSS.n925 3.29193
R14929 VSS.n945 VSS.n891 3.29193
R14930 VSS.n1304 VSS.n1295 3.29193
R14931 VSS.n17872 VSS.n17871 3.29193
R14932 VSS.n1284 VSS.n1283 3.2005
R14933 VSS.n1150 VSS.n1149 3.2005
R14934 VSS.n17101 VSS.n17100 3.2005
R14935 VSS.n17437 VSS.n17436 3.2005
R14936 VSS.n17693 VSS.n17692 3.2005
R14937 VSS.n18301 VSS.n18300 3.2005
R14938 VSS.n229 VSS.n228 3.2005
R14939 VSS.n9743 VSS.n9742 3.2005
R14940 VSS.n9487 VSS.n9486 3.2005
R14941 VSS.n16686 VSS.n16685 3.2005
R14942 VSS.n16582 VSS.n16581 3.2005
R14943 VSS.n16093 VSS.n16092 3.2005
R14944 VSS.n1747 VSS.n1746 3.2005
R14945 VSS.n2066 VSS.n2065 3.2005
R14946 VSS.n1779 VSS.n1778 3.2005
R14947 VSS.n3234 VSS.n3233 3.2005
R14948 VSS.n2978 VSS.n2977 3.2005
R14949 VSS.n3826 VSS.n3825 3.2005
R14950 VSS.n3570 VSS.n3569 3.2005
R14951 VSS.n4418 VSS.n4417 3.2005
R14952 VSS.n4162 VSS.n4161 3.2005
R14953 VSS.n5010 VSS.n5009 3.2005
R14954 VSS.n4754 VSS.n4753 3.2005
R14955 VSS.n2662 VSS.n2661 3.2005
R14956 VSS.n2375 VSS.n2374 3.2005
R14957 VSS.n5623 VSS.n5622 3.2005
R14958 VSS.n5336 VSS.n5335 3.2005
R14959 VSS.n6196 VSS.n6195 3.2005
R14960 VSS.n5909 VSS.n5908 3.2005
R14961 VSS.n7967 VSS.n7966 3.2005
R14962 VSS.n7711 VSS.n7710 3.2005
R14963 VSS.n8559 VSS.n8558 3.2005
R14964 VSS.n8303 VSS.n8302 3.2005
R14965 VSS.n9151 VSS.n9150 3.2005
R14966 VSS.n8895 VSS.n8894 3.2005
R14967 VSS.n10335 VSS.n10334 3.2005
R14968 VSS.n10079 VSS.n10078 3.2005
R14969 VSS.n10927 VSS.n10926 3.2005
R14970 VSS.n10671 VSS.n10670 3.2005
R14971 VSS.n11519 VSS.n11518 3.2005
R14972 VSS.n11263 VSS.n11262 3.2005
R14973 VSS.n12111 VSS.n12110 3.2005
R14974 VSS.n11855 VSS.n11854 3.2005
R14975 VSS.n12703 VSS.n12702 3.2005
R14976 VSS.n12447 VSS.n12446 3.2005
R14977 VSS.n13295 VSS.n13294 3.2005
R14978 VSS.n13039 VSS.n13038 3.2005
R14979 VSS.n13887 VSS.n13886 3.2005
R14980 VSS.n13631 VSS.n13630 3.2005
R14981 VSS.n14479 VSS.n14478 3.2005
R14982 VSS.n14223 VSS.n14222 3.2005
R14983 VSS.n15071 VSS.n15070 3.2005
R14984 VSS.n14815 VSS.n14814 3.2005
R14985 VSS.n15663 VSS.n15662 3.2005
R14986 VSS.n15407 VSS.n15406 3.2005
R14987 VSS.n6802 VSS.n6801 3.2005
R14988 VSS.n6515 VSS.n6514 3.2005
R14989 VSS.n7375 VSS.n7374 3.2005
R14990 VSS.n7271 VSS.n7270 3.2005
R14991 VSS.n18687 VSS.n18686 3.2005
R14992 VSS.n404 VSS.n403 3.2005
R14993 VSS.n625 VSS.n624 3.2005
R14994 VSS.n969 VSS.n968 3.2005
R14995 VSS.n17056 VSS.n17055 3.03311
R14996 VSS.n17026 VSS.n17025 3.03311
R14997 VSS.n17648 VSS.n17647 3.03311
R14998 VSS.n17618 VSS.n17617 3.03311
R14999 VSS.n18132 VSS.n18131 3.03311
R15000 VSS.n18097 VSS.n18096 3.03311
R15001 VSS.n9698 VSS.n9697 3.03311
R15002 VSS.n9668 VSS.n9667 3.03311
R15003 VSS.n9570 VSS.n9569 3.03311
R15004 VSS.n9605 VSS.n9604 3.03311
R15005 VSS.n16641 VSS.n16640 3.03311
R15006 VSS.n16611 VSS.n16610 3.03311
R15007 VSS.n16536 VSS.n16535 3.03311
R15008 VSS.n16506 VSS.n16505 3.03311
R15009 VSS.n16048 VSS.n16047 3.03311
R15010 VSS.n16018 VSS.n16017 3.03311
R15011 VSS.n1701 VSS.n1700 3.03311
R15012 VSS.n1671 VSS.n1670 3.03311
R15013 VSS.n1992 VSS.n1961 3.03311
R15014 VSS.n2016 VSS.n2015 3.03311
R15015 VSS.n1897 VSS.n1896 3.03311
R15016 VSS.n1862 VSS.n1861 3.03311
R15017 VSS.n3189 VSS.n3188 3.03311
R15018 VSS.n3159 VSS.n3158 3.03311
R15019 VSS.n3096 VSS.n3095 3.03311
R15020 VSS.n3061 VSS.n3060 3.03311
R15021 VSS.n3781 VSS.n3780 3.03311
R15022 VSS.n3751 VSS.n3750 3.03311
R15023 VSS.n3688 VSS.n3687 3.03311
R15024 VSS.n3653 VSS.n3652 3.03311
R15025 VSS.n4373 VSS.n4372 3.03311
R15026 VSS.n4343 VSS.n4342 3.03311
R15027 VSS.n4280 VSS.n4279 3.03311
R15028 VSS.n4245 VSS.n4244 3.03311
R15029 VSS.n4965 VSS.n4964 3.03311
R15030 VSS.n4935 VSS.n4934 3.03311
R15031 VSS.n4872 VSS.n4871 3.03311
R15032 VSS.n4837 VSS.n4836 3.03311
R15033 VSS.n2588 VSS.n2557 3.03311
R15034 VSS.n2612 VSS.n2611 3.03311
R15035 VSS.n2493 VSS.n2492 3.03311
R15036 VSS.n2458 VSS.n2457 3.03311
R15037 VSS.n5549 VSS.n5518 3.03311
R15038 VSS.n5573 VSS.n5572 3.03311
R15039 VSS.n5454 VSS.n5453 3.03311
R15040 VSS.n5419 VSS.n5418 3.03311
R15041 VSS.n6122 VSS.n6091 3.03311
R15042 VSS.n6146 VSS.n6145 3.03311
R15043 VSS.n6027 VSS.n6026 3.03311
R15044 VSS.n5992 VSS.n5991 3.03311
R15045 VSS.n7922 VSS.n7921 3.03311
R15046 VSS.n7892 VSS.n7891 3.03311
R15047 VSS.n7829 VSS.n7828 3.03311
R15048 VSS.n7794 VSS.n7793 3.03311
R15049 VSS.n8514 VSS.n8513 3.03311
R15050 VSS.n8484 VSS.n8483 3.03311
R15051 VSS.n8421 VSS.n8420 3.03311
R15052 VSS.n8386 VSS.n8385 3.03311
R15053 VSS.n9106 VSS.n9105 3.03311
R15054 VSS.n9076 VSS.n9075 3.03311
R15055 VSS.n9013 VSS.n9012 3.03311
R15056 VSS.n8978 VSS.n8977 3.03311
R15057 VSS.n10290 VSS.n10289 3.03311
R15058 VSS.n10260 VSS.n10259 3.03311
R15059 VSS.n10197 VSS.n10196 3.03311
R15060 VSS.n10162 VSS.n10161 3.03311
R15061 VSS.n10882 VSS.n10881 3.03311
R15062 VSS.n10852 VSS.n10851 3.03311
R15063 VSS.n10789 VSS.n10788 3.03311
R15064 VSS.n10754 VSS.n10753 3.03311
R15065 VSS.n11474 VSS.n11473 3.03311
R15066 VSS.n11444 VSS.n11443 3.03311
R15067 VSS.n11381 VSS.n11380 3.03311
R15068 VSS.n11346 VSS.n11345 3.03311
R15069 VSS.n12066 VSS.n12065 3.03311
R15070 VSS.n12036 VSS.n12035 3.03311
R15071 VSS.n11973 VSS.n11972 3.03311
R15072 VSS.n11938 VSS.n11937 3.03311
R15073 VSS.n12658 VSS.n12657 3.03311
R15074 VSS.n12628 VSS.n12627 3.03311
R15075 VSS.n12565 VSS.n12564 3.03311
R15076 VSS.n12530 VSS.n12529 3.03311
R15077 VSS.n13250 VSS.n13249 3.03311
R15078 VSS.n13220 VSS.n13219 3.03311
R15079 VSS.n13157 VSS.n13156 3.03311
R15080 VSS.n13122 VSS.n13121 3.03311
R15081 VSS.n13842 VSS.n13841 3.03311
R15082 VSS.n13812 VSS.n13811 3.03311
R15083 VSS.n13749 VSS.n13748 3.03311
R15084 VSS.n13714 VSS.n13713 3.03311
R15085 VSS.n14434 VSS.n14433 3.03311
R15086 VSS.n14404 VSS.n14403 3.03311
R15087 VSS.n14341 VSS.n14340 3.03311
R15088 VSS.n14306 VSS.n14305 3.03311
R15089 VSS.n15026 VSS.n15025 3.03311
R15090 VSS.n14996 VSS.n14995 3.03311
R15091 VSS.n14933 VSS.n14932 3.03311
R15092 VSS.n14898 VSS.n14897 3.03311
R15093 VSS.n15618 VSS.n15617 3.03311
R15094 VSS.n15588 VSS.n15587 3.03311
R15095 VSS.n15525 VSS.n15524 3.03311
R15096 VSS.n15490 VSS.n15489 3.03311
R15097 VSS.n6728 VSS.n6697 3.03311
R15098 VSS.n6752 VSS.n6751 3.03311
R15099 VSS.n6633 VSS.n6632 3.03311
R15100 VSS.n6598 VSS.n6597 3.03311
R15101 VSS.n7330 VSS.n7329 3.03311
R15102 VSS.n7300 VSS.n7299 3.03311
R15103 VSS.n7225 VSS.n7224 3.03311
R15104 VSS.n7195 VSS.n7194 3.03311
R15105 VSS.n18642 VSS.n18641 3.03311
R15106 VSS.n18612 VSS.n18611 3.03311
R15107 VSS.n379 VSS.n378 3.03311
R15108 VSS.n346 VSS.n343 3.03311
R15109 VSS.n18227 VSS.n18196 3.03311
R15110 VSS.n18251 VSS.n18250 3.03311
R15111 VSS.n548 VSS.n517 3.03311
R15112 VSS.n575 VSS.n574 3.03311
R15113 VSS.n896 VSS.n895 3.03311
R15114 VSS.n920 VSS.n919 3.03311
R15115 VSS.n1077 VSS.n1076 3.03311
R15116 VSS.n1101 VSS.n1100 3.03311
R15117 VSS.n17555 VSS.n17554 3.03311
R15118 VSS.n17520 VSS.n17519 3.03311
R15119 VSS.n1210 VSS.n1179 3.03311
R15120 VSS.n1234 VSS.n1233 3.03311
R15121 VSS.n1248 VSS.n1213 2.81479
R15122 VSS.n1269 VSS.n1209 2.81479
R15123 VSS.n17530 VSS.n17480 2.81479
R15124 VSS.n17563 VSS.n17450 2.81479
R15125 VSS.n1113 VSS.n1080 2.81479
R15126 VSS.n1134 VSS.n1075 2.81479
R15127 VSS.n932 VSS.n899 2.81479
R15128 VSS.n953 VSS.n894 2.81479
R15129 VSS.n17049 VSS.n16975 2.81479
R15130 VSS.n17080 VSS.n16954 2.81479
R15131 VSS.n17641 VSS.n17389 2.81479
R15132 VSS.n17672 VSS.n17368 2.81479
R15133 VSS.n18265 VSS.n18230 2.81479
R15134 VSS.n18286 VSS.n18226 2.81479
R15135 VSS.n18107 VSS.n272 2.81479
R15136 VSS.n18140 VSS.n242 2.81479
R15137 VSS.n9580 VSS.n9530 2.81479
R15138 VSS.n9613 VSS.n9500 2.81479
R15139 VSS.n9691 VSS.n9439 2.81479
R15140 VSS.n9722 VSS.n9418 2.81479
R15141 VSS.n16529 VSS.n16458 2.81479
R15142 VSS.n16560 VSS.n16435 2.81479
R15143 VSS.n16634 VSS.n16381 2.81479
R15144 VSS.n16665 VSS.n16360 2.81479
R15145 VSS.n1694 VSS.n1623 2.81479
R15146 VSS.n1725 VSS.n1600 2.81479
R15147 VSS.n16041 VSS.n1553 2.81479
R15148 VSS.n16072 VSS.n1532 2.81479
R15149 VSS.n1872 VSS.n1822 2.81479
R15150 VSS.n1905 VSS.n1792 2.81479
R15151 VSS.n2030 VSS.n1995 2.81479
R15152 VSS.n2051 VSS.n1991 2.81479
R15153 VSS.n3071 VSS.n3021 2.81479
R15154 VSS.n3104 VSS.n2991 2.81479
R15155 VSS.n3182 VSS.n2930 2.81479
R15156 VSS.n3213 VSS.n2909 2.81479
R15157 VSS.n3663 VSS.n3613 2.81479
R15158 VSS.n3696 VSS.n3583 2.81479
R15159 VSS.n3774 VSS.n3522 2.81479
R15160 VSS.n3805 VSS.n3501 2.81479
R15161 VSS.n4255 VSS.n4205 2.81479
R15162 VSS.n4288 VSS.n4175 2.81479
R15163 VSS.n4366 VSS.n4114 2.81479
R15164 VSS.n4397 VSS.n4093 2.81479
R15165 VSS.n4847 VSS.n4797 2.81479
R15166 VSS.n4880 VSS.n4767 2.81479
R15167 VSS.n4958 VSS.n4706 2.81479
R15168 VSS.n4989 VSS.n4685 2.81479
R15169 VSS.n2468 VSS.n2418 2.81479
R15170 VSS.n2501 VSS.n2388 2.81479
R15171 VSS.n2626 VSS.n2591 2.81479
R15172 VSS.n2647 VSS.n2587 2.81479
R15173 VSS.n5429 VSS.n5379 2.81479
R15174 VSS.n5462 VSS.n5349 2.81479
R15175 VSS.n5587 VSS.n5552 2.81479
R15176 VSS.n5608 VSS.n5548 2.81479
R15177 VSS.n6002 VSS.n5952 2.81479
R15178 VSS.n6035 VSS.n5922 2.81479
R15179 VSS.n6160 VSS.n6125 2.81479
R15180 VSS.n6181 VSS.n6121 2.81479
R15181 VSS.n7804 VSS.n7754 2.81479
R15182 VSS.n7837 VSS.n7724 2.81479
R15183 VSS.n7915 VSS.n7663 2.81479
R15184 VSS.n7946 VSS.n7642 2.81479
R15185 VSS.n8396 VSS.n8346 2.81479
R15186 VSS.n8429 VSS.n8316 2.81479
R15187 VSS.n8507 VSS.n8255 2.81479
R15188 VSS.n8538 VSS.n8234 2.81479
R15189 VSS.n8988 VSS.n8938 2.81479
R15190 VSS.n9021 VSS.n8908 2.81479
R15191 VSS.n9099 VSS.n8847 2.81479
R15192 VSS.n9130 VSS.n8826 2.81479
R15193 VSS.n10172 VSS.n10122 2.81479
R15194 VSS.n10205 VSS.n10092 2.81479
R15195 VSS.n10283 VSS.n10031 2.81479
R15196 VSS.n10314 VSS.n10010 2.81479
R15197 VSS.n10764 VSS.n10714 2.81479
R15198 VSS.n10797 VSS.n10684 2.81479
R15199 VSS.n10875 VSS.n10623 2.81479
R15200 VSS.n10906 VSS.n10602 2.81479
R15201 VSS.n11356 VSS.n11306 2.81479
R15202 VSS.n11389 VSS.n11276 2.81479
R15203 VSS.n11467 VSS.n11215 2.81479
R15204 VSS.n11498 VSS.n11194 2.81479
R15205 VSS.n11948 VSS.n11898 2.81479
R15206 VSS.n11981 VSS.n11868 2.81479
R15207 VSS.n12059 VSS.n11807 2.81479
R15208 VSS.n12090 VSS.n11786 2.81479
R15209 VSS.n12540 VSS.n12490 2.81479
R15210 VSS.n12573 VSS.n12460 2.81479
R15211 VSS.n12651 VSS.n12399 2.81479
R15212 VSS.n12682 VSS.n12378 2.81479
R15213 VSS.n13132 VSS.n13082 2.81479
R15214 VSS.n13165 VSS.n13052 2.81479
R15215 VSS.n13243 VSS.n12991 2.81479
R15216 VSS.n13274 VSS.n12970 2.81479
R15217 VSS.n13724 VSS.n13674 2.81479
R15218 VSS.n13757 VSS.n13644 2.81479
R15219 VSS.n13835 VSS.n13583 2.81479
R15220 VSS.n13866 VSS.n13562 2.81479
R15221 VSS.n14316 VSS.n14266 2.81479
R15222 VSS.n14349 VSS.n14236 2.81479
R15223 VSS.n14427 VSS.n14175 2.81479
R15224 VSS.n14458 VSS.n14154 2.81479
R15225 VSS.n14908 VSS.n14858 2.81479
R15226 VSS.n14941 VSS.n14828 2.81479
R15227 VSS.n15019 VSS.n14767 2.81479
R15228 VSS.n15050 VSS.n14746 2.81479
R15229 VSS.n15500 VSS.n15450 2.81479
R15230 VSS.n15533 VSS.n15420 2.81479
R15231 VSS.n15611 VSS.n15359 2.81479
R15232 VSS.n15642 VSS.n15338 2.81479
R15233 VSS.n6608 VSS.n6558 2.81479
R15234 VSS.n6641 VSS.n6528 2.81479
R15235 VSS.n6766 VSS.n6731 2.81479
R15236 VSS.n6787 VSS.n6727 2.81479
R15237 VSS.n7218 VSS.n7147 2.81479
R15238 VSS.n7249 VSS.n7124 2.81479
R15239 VSS.n7323 VSS.n7070 2.81479
R15240 VSS.n7354 VSS.n7049 2.81479
R15241 VSS.n372 VSS.n339 2.81479
R15242 VSS.n385 VSS.n335 2.81479
R15243 VSS.n18635 VSS.n168 2.81479
R15244 VSS.n18666 VSS.n147 2.81479
R15245 VSS.n589 VSS.n551 2.81479
R15246 VSS.n610 VSS.n547 2.81479
R15247 VSS.n17221 VSS.n17220 2.5605
R15248 VSS.n17813 VSS.n17812 2.5605
R15249 VSS.n18491 VSS.n18490 2.5605
R15250 VSS.n9863 VSS.n9862 2.5605
R15251 VSS.n16806 VSS.n16805 2.5605
R15252 VSS.n16213 VSS.n16212 2.5605
R15253 VSS.n2250 VSS.n2157 2.5605
R15254 VSS.n3354 VSS.n3353 2.5605
R15255 VSS.n3946 VSS.n3945 2.5605
R15256 VSS.n4538 VSS.n4537 2.5605
R15257 VSS.n5130 VSS.n5129 2.5605
R15258 VSS.n5215 VSS.n2753 2.5605
R15259 VSS.n5788 VSS.n5714 2.5605
R15260 VSS.n6380 VSS.n6287 2.5605
R15261 VSS.n8087 VSS.n8086 2.5605
R15262 VSS.n8679 VSS.n8678 2.5605
R15263 VSS.n9271 VSS.n9270 2.5605
R15264 VSS.n10455 VSS.n10454 2.5605
R15265 VSS.n11047 VSS.n11046 2.5605
R15266 VSS.n11639 VSS.n11638 2.5605
R15267 VSS.n12231 VSS.n12230 2.5605
R15268 VSS.n12823 VSS.n12822 2.5605
R15269 VSS.n13415 VSS.n13414 2.5605
R15270 VSS.n14007 VSS.n14006 2.5605
R15271 VSS.n14599 VSS.n14598 2.5605
R15272 VSS.n15191 VSS.n15190 2.5605
R15273 VSS.n15783 VSS.n15782 2.5605
R15274 VSS.n15868 VSS.n6893 2.5605
R15275 VSS.n7495 VSS.n7494 2.5605
R15276 VSS.n18807 VSS.n18806 2.5605
R15277 VSS.n782 VSS.n716 2.5605
R15278 VSS.n17896 VSS.n1375 2.5605
R15279 VSS.n17170 VSS.n17169 2.46907
R15280 VSS.n17762 VSS.n17761 2.46907
R15281 VSS.n18509 VSS.n18344 2.46907
R15282 VSS.n9812 VSS.n9811 2.46907
R15283 VSS.n16755 VSS.n16754 2.46907
R15284 VSS.n16162 VSS.n16161 2.46907
R15285 VSS.n2269 VSS.n2268 2.46907
R15286 VSS.n3303 VSS.n3302 2.46907
R15287 VSS.n3895 VSS.n3894 2.46907
R15288 VSS.n4487 VSS.n4486 2.46907
R15289 VSS.n5079 VSS.n5078 2.46907
R15290 VSS.n5234 VSS.n5233 2.46907
R15291 VSS.n5807 VSS.n5806 2.46907
R15292 VSS.n6399 VSS.n6398 2.46907
R15293 VSS.n8036 VSS.n8035 2.46907
R15294 VSS.n8628 VSS.n8627 2.46907
R15295 VSS.n9220 VSS.n9219 2.46907
R15296 VSS.n10404 VSS.n10403 2.46907
R15297 VSS.n10996 VSS.n10995 2.46907
R15298 VSS.n11588 VSS.n11587 2.46907
R15299 VSS.n12180 VSS.n12179 2.46907
R15300 VSS.n12772 VSS.n12771 2.46907
R15301 VSS.n13364 VSS.n13363 2.46907
R15302 VSS.n13956 VSS.n13955 2.46907
R15303 VSS.n14548 VSS.n14547 2.46907
R15304 VSS.n15140 VSS.n15139 2.46907
R15305 VSS.n15732 VSS.n15731 2.46907
R15306 VSS.n15887 VSS.n15886 2.46907
R15307 VSS.n7444 VSS.n7443 2.46907
R15308 VSS.n18756 VSS.n18755 2.46907
R15309 VSS.n801 VSS.n800 2.46907
R15310 VSS.n17915 VSS.n17914 2.46907
R15311 VSS.n17560 VSS.t409 2.42341
R15312 VSS.n17240 VSS.n17239 2.37764
R15313 VSS.n17832 VSS.n17831 2.37764
R15314 VSS.n18481 VSS.n18420 2.37764
R15315 VSS.n9882 VSS.n9881 2.37764
R15316 VSS.n16825 VSS.n16824 2.37764
R15317 VSS.n16232 VSS.n16231 2.37764
R15318 VSS.n2193 VSS.n2192 2.37764
R15319 VSS.n3373 VSS.n3372 2.37764
R15320 VSS.n3965 VSS.n3964 2.37764
R15321 VSS.n4557 VSS.n4556 2.37764
R15322 VSS.n5149 VSS.n5148 2.37764
R15323 VSS.n2789 VSS.n2788 2.37764
R15324 VSS.n5763 VSS.n5762 2.37764
R15325 VSS.n6323 VSS.n6322 2.37764
R15326 VSS.n8106 VSS.n8105 2.37764
R15327 VSS.n8698 VSS.n8697 2.37764
R15328 VSS.n9290 VSS.n9289 2.37764
R15329 VSS.n10474 VSS.n10473 2.37764
R15330 VSS.n11066 VSS.n11065 2.37764
R15331 VSS.n11658 VSS.n11657 2.37764
R15332 VSS.n12250 VSS.n12249 2.37764
R15333 VSS.n12842 VSS.n12841 2.37764
R15334 VSS.n13434 VSS.n13433 2.37764
R15335 VSS.n14026 VSS.n14025 2.37764
R15336 VSS.n14618 VSS.n14617 2.37764
R15337 VSS.n15210 VSS.n15209 2.37764
R15338 VSS.n15802 VSS.n15801 2.37764
R15339 VSS.n6929 VSS.n6928 2.37764
R15340 VSS.n7514 VSS.n7513 2.37764
R15341 VSS.n18826 VSS.n18825 2.37764
R15342 VSS.n763 VSS.n762 2.37764
R15343 VSS.n1411 VSS.n1410 2.37764
R15344 VSS.n17152 VSS.n16917 2.28621
R15345 VSS.n17744 VSS.n17331 2.28621
R15346 VSS.n18367 VSS.n18365 2.28621
R15347 VSS.n9794 VSS.n9381 2.28621
R15348 VSS.n16737 VSS.n16323 2.28621
R15349 VSS.n16144 VSS.n1495 2.28621
R15350 VSS.n2284 VSS.n2283 2.28621
R15351 VSS.n3285 VSS.n2872 2.28621
R15352 VSS.n3877 VSS.n3464 2.28621
R15353 VSS.n4469 VSS.n4056 2.28621
R15354 VSS.n5061 VSS.n4648 2.28621
R15355 VSS.n5249 VSS.n5248 2.28621
R15356 VSS.n5822 VSS.n5821 2.28621
R15357 VSS.n6414 VSS.n6413 2.28621
R15358 VSS.n8018 VSS.n7605 2.28621
R15359 VSS.n8610 VSS.n8197 2.28621
R15360 VSS.n9202 VSS.n8789 2.28621
R15361 VSS.n10386 VSS.n9973 2.28621
R15362 VSS.n10978 VSS.n10565 2.28621
R15363 VSS.n11570 VSS.n11157 2.28621
R15364 VSS.n12162 VSS.n11749 2.28621
R15365 VSS.n12754 VSS.n12341 2.28621
R15366 VSS.n13346 VSS.n12933 2.28621
R15367 VSS.n13938 VSS.n13525 2.28621
R15368 VSS.n14530 VSS.n14117 2.28621
R15369 VSS.n15122 VSS.n14709 2.28621
R15370 VSS.n15714 VSS.n15301 2.28621
R15371 VSS.n15902 VSS.n15901 2.28621
R15372 VSS.n7426 VSS.n7012 2.28621
R15373 VSS.n18738 VSS.n110 2.28621
R15374 VSS.n816 VSS.n815 2.28621
R15375 VSS.n17930 VSS.n17929 2.28621
R15376 VSS.n17866 VSS.n17865 2.27261
R15377 VSS.n7548 VSS.n53 2.27256
R15378 VSS.n15244 VSS.n14652 2.27256
R15379 VSS.n12876 VSS.n12284 2.27256
R15380 VSS.n10508 VSS.n9916 2.27256
R15381 VSS.n8140 VSS.n0 2.27256
R15382 VSS.n5183 VSS.n4591 2.27256
R15383 VSS.n16266 VSS.n1438 2.27256
R15384 VSS.n1194 VSS.n1192 2.2505
R15385 VSS.n1260 VSS.n1183 2.2505
R15386 VSS.n1190 VSS.n1189 2.2505
R15387 VSS.n1165 VSS.n1163 2.2505
R15388 VSS.n1171 VSS.n1169 2.2505
R15389 VSS.n1226 VSS.n1225 2.2505
R15390 VSS.n1060 VSS.n1058 2.2505
R15391 VSS.n1125 VSS.n1049 2.2505
R15392 VSS.n1056 VSS.n1055 2.2505
R15393 VSS.n1030 VSS.n1028 2.2505
R15394 VSS.n1036 VSS.n1034 2.2505
R15395 VSS.n1093 VSS.n1092 2.2505
R15396 VSS.n17256 VSS.n16872 2.2505
R15397 VSS.n17203 VSS.n17193 2.2505
R15398 VSS.n17232 VSS.n17231 2.2505
R15399 VSS.n17157 VSS.n16919 2.2505
R15400 VSS.n17180 VSS.n17179 2.2505
R15401 VSS.n17182 VSS.n16902 2.2505
R15402 VSS.n16925 VSS.n16923 2.2505
R15403 VSS.n17095 VSS.n17094 2.2505
R15404 VSS.n16959 VSS.n16957 2.2505
R15405 VSS.n17088 VSS.n16946 2.2505
R15406 VSS.n17024 VSS.n17023 2.2505
R15407 VSS.n17045 VSS.n17044 2.2505
R15408 VSS.n17017 VSS.n16998 2.2505
R15409 VSS.n17580 VSS.n17579 2.2505
R15410 VSS.n17566 VSS.n17445 2.2505
R15411 VSS.n17432 VSS.n17430 2.2505
R15412 VSS.n17518 VSS.n17517 2.2505
R15413 VSS.n17475 VSS.n17474 2.2505
R15414 VSS.n17511 VSS.n17492 2.2505
R15415 VSS.n17848 VSS.n17286 2.2505
R15416 VSS.n17795 VSS.n17785 2.2505
R15417 VSS.n17824 VSS.n17823 2.2505
R15418 VSS.n17749 VSS.n17333 2.2505
R15419 VSS.n17772 VSS.n17771 2.2505
R15420 VSS.n17774 VSS.n17316 2.2505
R15421 VSS.n17339 VSS.n17337 2.2505
R15422 VSS.n17687 VSS.n17686 2.2505
R15423 VSS.n17373 VSS.n17371 2.2505
R15424 VSS.n17680 VSS.n17360 2.2505
R15425 VSS.n17616 VSS.n17615 2.2505
R15426 VSS.n17637 VSS.n17636 2.2505
R15427 VSS.n17609 VSS.n17412 2.2505
R15428 VSS.n18211 VSS.n18209 2.2505
R15429 VSS.n18277 VSS.n18200 2.2505
R15430 VSS.n18207 VSS.n18206 2.2505
R15431 VSS.n18182 VSS.n18180 2.2505
R15432 VSS.n18188 VSS.n18186 2.2505
R15433 VSS.n18243 VSS.n18242 2.2505
R15434 VSS.n18476 VSS.n18423 2.2505
R15435 VSS.n18408 VSS.n18393 2.2505
R15436 VSS.n18446 VSS.n18445 2.2505
R15437 VSS.n18516 VSS.n18515 2.2505
R15438 VSS.n18347 VSS.n18345 2.2505
R15439 VSS.n18377 VSS.n18353 2.2505
R15440 VSS.n18526 VSS.n18315 2.2505
R15441 VSS.n18157 VSS.n18156 2.2505
R15442 VSS.n18143 VSS.n237 2.2505
R15443 VSS.n224 VSS.n222 2.2505
R15444 VSS.n18095 VSS.n18094 2.2505
R15445 VSS.n267 VSS.n266 2.2505
R15446 VSS.n18088 VSS.n284 2.2505
R15447 VSS.n9737 VSS.n9736 2.2505
R15448 VSS.n9423 VSS.n9421 2.2505
R15449 VSS.n9730 VSS.n9410 2.2505
R15450 VSS.n9666 VSS.n9665 2.2505
R15451 VSS.n9687 VSS.n9686 2.2505
R15452 VSS.n9659 VSS.n9462 2.2505
R15453 VSS.n9899 VSS.n9898 2.2505
R15454 VSS.n9845 VSS.n9835 2.2505
R15455 VSS.n9874 VSS.n9873 2.2505
R15456 VSS.n9799 VSS.n9383 2.2505
R15457 VSS.n9822 VSS.n9821 2.2505
R15458 VSS.n9824 VSS.n9366 2.2505
R15459 VSS.n9389 VSS.n9387 2.2505
R15460 VSS.n9630 VSS.n9629 2.2505
R15461 VSS.n9482 VSS.n9480 2.2505
R15462 VSS.n9616 VSS.n9495 2.2505
R15463 VSS.n9561 VSS.n9542 2.2505
R15464 VSS.n9568 VSS.n9567 2.2505
R15465 VSS.n9525 VSS.n9524 2.2505
R15466 VSS.n16680 VSS.n16679 2.2505
R15467 VSS.n16365 VSS.n16363 2.2505
R15468 VSS.n16673 VSS.n16352 2.2505
R15469 VSS.n16609 VSS.n16608 2.2505
R15470 VSS.n16630 VSS.n16629 2.2505
R15471 VSS.n16602 VSS.n16404 2.2505
R15472 VSS.n16842 VSS.n16841 2.2505
R15473 VSS.n16788 VSS.n16778 2.2505
R15474 VSS.n16817 VSS.n16816 2.2505
R15475 VSS.n16742 VSS.n16325 2.2505
R15476 VSS.n16765 VSS.n16764 2.2505
R15477 VSS.n16767 VSS.n16308 2.2505
R15478 VSS.n16331 VSS.n16329 2.2505
R15479 VSS.n16576 VSS.n16575 2.2505
R15480 VSS.n16440 VSS.n16438 2.2505
R15481 VSS.n16569 VSS.n16427 2.2505
R15482 VSS.n16504 VSS.n16503 2.2505
R15483 VSS.n16525 VSS.n16524 2.2505
R15484 VSS.n16497 VSS.n16479 2.2505
R15485 VSS.n16087 VSS.n16086 2.2505
R15486 VSS.n1537 VSS.n1535 2.2505
R15487 VSS.n16080 VSS.n1524 2.2505
R15488 VSS.n16016 VSS.n16015 2.2505
R15489 VSS.n16037 VSS.n16036 2.2505
R15490 VSS.n16009 VSS.n1576 2.2505
R15491 VSS.n16249 VSS.n16248 2.2505
R15492 VSS.n16195 VSS.n16185 2.2505
R15493 VSS.n16224 VSS.n16223 2.2505
R15494 VSS.n16149 VSS.n1497 2.2505
R15495 VSS.n16172 VSS.n16171 2.2505
R15496 VSS.n16174 VSS.n1480 2.2505
R15497 VSS.n1503 VSS.n1501 2.2505
R15498 VSS.n1741 VSS.n1740 2.2505
R15499 VSS.n1605 VSS.n1603 2.2505
R15500 VSS.n1734 VSS.n1592 2.2505
R15501 VSS.n1669 VSS.n1668 2.2505
R15502 VSS.n1690 VSS.n1689 2.2505
R15503 VSS.n1662 VSS.n1644 2.2505
R15504 VSS.n1976 VSS.n1974 2.2505
R15505 VSS.n2042 VSS.n1965 2.2505
R15506 VSS.n1972 VSS.n1971 2.2505
R15507 VSS.n1947 VSS.n1945 2.2505
R15508 VSS.n1953 VSS.n1951 2.2505
R15509 VSS.n2008 VSS.n2007 2.2505
R15510 VSS.n2209 VSS.n2172 2.2505
R15511 VSS.n2155 VSS.n2153 2.2505
R15512 VSS.n2244 VSS.n2243 2.2505
R15513 VSS.n2110 VSS.n2108 2.2505
R15514 VSS.n2140 VSS.n2139 2.2505
R15515 VSS.n2142 VSS.n2132 2.2505
R15516 VSS.n2291 VSS.n2290 2.2505
R15517 VSS.n1922 VSS.n1921 2.2505
R15518 VSS.n1908 VSS.n1787 2.2505
R15519 VSS.n1774 VSS.n1772 2.2505
R15520 VSS.n1860 VSS.n1859 2.2505
R15521 VSS.n1817 VSS.n1816 2.2505
R15522 VSS.n1853 VSS.n1834 2.2505
R15523 VSS.n3228 VSS.n3227 2.2505
R15524 VSS.n2914 VSS.n2912 2.2505
R15525 VSS.n3221 VSS.n2901 2.2505
R15526 VSS.n3157 VSS.n3156 2.2505
R15527 VSS.n3178 VSS.n3177 2.2505
R15528 VSS.n3150 VSS.n2953 2.2505
R15529 VSS.n3390 VSS.n3389 2.2505
R15530 VSS.n3336 VSS.n3326 2.2505
R15531 VSS.n3365 VSS.n3364 2.2505
R15532 VSS.n3290 VSS.n2874 2.2505
R15533 VSS.n3313 VSS.n3312 2.2505
R15534 VSS.n3315 VSS.n2857 2.2505
R15535 VSS.n2880 VSS.n2878 2.2505
R15536 VSS.n3121 VSS.n3120 2.2505
R15537 VSS.n3107 VSS.n2986 2.2505
R15538 VSS.n2973 VSS.n2971 2.2505
R15539 VSS.n3059 VSS.n3058 2.2505
R15540 VSS.n3016 VSS.n3015 2.2505
R15541 VSS.n3052 VSS.n3033 2.2505
R15542 VSS.n3820 VSS.n3819 2.2505
R15543 VSS.n3506 VSS.n3504 2.2505
R15544 VSS.n3813 VSS.n3493 2.2505
R15545 VSS.n3749 VSS.n3748 2.2505
R15546 VSS.n3770 VSS.n3769 2.2505
R15547 VSS.n3742 VSS.n3545 2.2505
R15548 VSS.n3982 VSS.n3981 2.2505
R15549 VSS.n3928 VSS.n3918 2.2505
R15550 VSS.n3957 VSS.n3956 2.2505
R15551 VSS.n3882 VSS.n3466 2.2505
R15552 VSS.n3905 VSS.n3904 2.2505
R15553 VSS.n3907 VSS.n3449 2.2505
R15554 VSS.n3472 VSS.n3470 2.2505
R15555 VSS.n3713 VSS.n3712 2.2505
R15556 VSS.n3699 VSS.n3578 2.2505
R15557 VSS.n3565 VSS.n3563 2.2505
R15558 VSS.n3651 VSS.n3650 2.2505
R15559 VSS.n3608 VSS.n3607 2.2505
R15560 VSS.n3644 VSS.n3625 2.2505
R15561 VSS.n4412 VSS.n4411 2.2505
R15562 VSS.n4098 VSS.n4096 2.2505
R15563 VSS.n4405 VSS.n4085 2.2505
R15564 VSS.n4341 VSS.n4340 2.2505
R15565 VSS.n4362 VSS.n4361 2.2505
R15566 VSS.n4334 VSS.n4137 2.2505
R15567 VSS.n4574 VSS.n4573 2.2505
R15568 VSS.n4520 VSS.n4510 2.2505
R15569 VSS.n4549 VSS.n4548 2.2505
R15570 VSS.n4474 VSS.n4058 2.2505
R15571 VSS.n4497 VSS.n4496 2.2505
R15572 VSS.n4499 VSS.n4041 2.2505
R15573 VSS.n4064 VSS.n4062 2.2505
R15574 VSS.n4305 VSS.n4304 2.2505
R15575 VSS.n4291 VSS.n4170 2.2505
R15576 VSS.n4157 VSS.n4155 2.2505
R15577 VSS.n4243 VSS.n4242 2.2505
R15578 VSS.n4200 VSS.n4199 2.2505
R15579 VSS.n4236 VSS.n4217 2.2505
R15580 VSS.n5004 VSS.n5003 2.2505
R15581 VSS.n4690 VSS.n4688 2.2505
R15582 VSS.n4997 VSS.n4677 2.2505
R15583 VSS.n4933 VSS.n4932 2.2505
R15584 VSS.n4954 VSS.n4953 2.2505
R15585 VSS.n4926 VSS.n4729 2.2505
R15586 VSS.n5166 VSS.n5165 2.2505
R15587 VSS.n5112 VSS.n5102 2.2505
R15588 VSS.n5141 VSS.n5140 2.2505
R15589 VSS.n5066 VSS.n4650 2.2505
R15590 VSS.n5089 VSS.n5088 2.2505
R15591 VSS.n5091 VSS.n4633 2.2505
R15592 VSS.n4656 VSS.n4654 2.2505
R15593 VSS.n4897 VSS.n4896 2.2505
R15594 VSS.n4883 VSS.n4762 2.2505
R15595 VSS.n4749 VSS.n4747 2.2505
R15596 VSS.n4835 VSS.n4834 2.2505
R15597 VSS.n4792 VSS.n4791 2.2505
R15598 VSS.n4828 VSS.n4809 2.2505
R15599 VSS.n2572 VSS.n2570 2.2505
R15600 VSS.n2638 VSS.n2561 2.2505
R15601 VSS.n2568 VSS.n2567 2.2505
R15602 VSS.n2543 VSS.n2541 2.2505
R15603 VSS.n2549 VSS.n2547 2.2505
R15604 VSS.n2604 VSS.n2603 2.2505
R15605 VSS.n2805 VSS.n2768 2.2505
R15606 VSS.n2751 VSS.n2749 2.2505
R15607 VSS.n5209 VSS.n5208 2.2505
R15608 VSS.n2706 VSS.n2704 2.2505
R15609 VSS.n2736 VSS.n2735 2.2505
R15610 VSS.n2738 VSS.n2728 2.2505
R15611 VSS.n5256 VSS.n5255 2.2505
R15612 VSS.n2518 VSS.n2517 2.2505
R15613 VSS.n2504 VSS.n2383 2.2505
R15614 VSS.n2370 VSS.n2368 2.2505
R15615 VSS.n2456 VSS.n2455 2.2505
R15616 VSS.n2413 VSS.n2412 2.2505
R15617 VSS.n2449 VSS.n2430 2.2505
R15618 VSS.n5533 VSS.n5531 2.2505
R15619 VSS.n5599 VSS.n5522 2.2505
R15620 VSS.n5529 VSS.n5528 2.2505
R15621 VSS.n5504 VSS.n5502 2.2505
R15622 VSS.n5510 VSS.n5508 2.2505
R15623 VSS.n5565 VSS.n5564 2.2505
R15624 VSS.n5741 VSS.n5740 2.2505
R15625 VSS.n5712 VSS.n5710 2.2505
R15626 VSS.n5782 VSS.n5781 2.2505
R15627 VSS.n5667 VSS.n5665 2.2505
R15628 VSS.n5697 VSS.n5696 2.2505
R15629 VSS.n5699 VSS.n5689 2.2505
R15630 VSS.n5829 VSS.n5828 2.2505
R15631 VSS.n5479 VSS.n5478 2.2505
R15632 VSS.n5465 VSS.n5344 2.2505
R15633 VSS.n5331 VSS.n5329 2.2505
R15634 VSS.n5417 VSS.n5416 2.2505
R15635 VSS.n5374 VSS.n5373 2.2505
R15636 VSS.n5410 VSS.n5391 2.2505
R15637 VSS.n6106 VSS.n6104 2.2505
R15638 VSS.n6172 VSS.n6095 2.2505
R15639 VSS.n6102 VSS.n6101 2.2505
R15640 VSS.n6077 VSS.n6075 2.2505
R15641 VSS.n6083 VSS.n6081 2.2505
R15642 VSS.n6138 VSS.n6137 2.2505
R15643 VSS.n6339 VSS.n6302 2.2505
R15644 VSS.n6285 VSS.n6283 2.2505
R15645 VSS.n6374 VSS.n6373 2.2505
R15646 VSS.n6240 VSS.n6238 2.2505
R15647 VSS.n6270 VSS.n6269 2.2505
R15648 VSS.n6272 VSS.n6262 2.2505
R15649 VSS.n6421 VSS.n6420 2.2505
R15650 VSS.n6052 VSS.n6051 2.2505
R15651 VSS.n6038 VSS.n5917 2.2505
R15652 VSS.n5904 VSS.n5902 2.2505
R15653 VSS.n5990 VSS.n5989 2.2505
R15654 VSS.n5947 VSS.n5946 2.2505
R15655 VSS.n5983 VSS.n5964 2.2505
R15656 VSS.n7961 VSS.n7960 2.2505
R15657 VSS.n7647 VSS.n7645 2.2505
R15658 VSS.n7954 VSS.n7634 2.2505
R15659 VSS.n7890 VSS.n7889 2.2505
R15660 VSS.n7911 VSS.n7910 2.2505
R15661 VSS.n7883 VSS.n7686 2.2505
R15662 VSS.n8123 VSS.n8122 2.2505
R15663 VSS.n8069 VSS.n8059 2.2505
R15664 VSS.n8098 VSS.n8097 2.2505
R15665 VSS.n8023 VSS.n7607 2.2505
R15666 VSS.n8046 VSS.n8045 2.2505
R15667 VSS.n8048 VSS.n7590 2.2505
R15668 VSS.n7613 VSS.n7611 2.2505
R15669 VSS.n7854 VSS.n7853 2.2505
R15670 VSS.n7840 VSS.n7719 2.2505
R15671 VSS.n7706 VSS.n7704 2.2505
R15672 VSS.n7792 VSS.n7791 2.2505
R15673 VSS.n7749 VSS.n7748 2.2505
R15674 VSS.n7785 VSS.n7766 2.2505
R15675 VSS.n8553 VSS.n8552 2.2505
R15676 VSS.n8239 VSS.n8237 2.2505
R15677 VSS.n8546 VSS.n8226 2.2505
R15678 VSS.n8482 VSS.n8481 2.2505
R15679 VSS.n8503 VSS.n8502 2.2505
R15680 VSS.n8475 VSS.n8278 2.2505
R15681 VSS.n8715 VSS.n8714 2.2505
R15682 VSS.n8661 VSS.n8651 2.2505
R15683 VSS.n8690 VSS.n8689 2.2505
R15684 VSS.n8615 VSS.n8199 2.2505
R15685 VSS.n8638 VSS.n8637 2.2505
R15686 VSS.n8640 VSS.n8182 2.2505
R15687 VSS.n8205 VSS.n8203 2.2505
R15688 VSS.n8446 VSS.n8445 2.2505
R15689 VSS.n8432 VSS.n8311 2.2505
R15690 VSS.n8298 VSS.n8296 2.2505
R15691 VSS.n8384 VSS.n8383 2.2505
R15692 VSS.n8341 VSS.n8340 2.2505
R15693 VSS.n8377 VSS.n8358 2.2505
R15694 VSS.n9145 VSS.n9144 2.2505
R15695 VSS.n8831 VSS.n8829 2.2505
R15696 VSS.n9138 VSS.n8818 2.2505
R15697 VSS.n9074 VSS.n9073 2.2505
R15698 VSS.n9095 VSS.n9094 2.2505
R15699 VSS.n9067 VSS.n8870 2.2505
R15700 VSS.n9307 VSS.n9306 2.2505
R15701 VSS.n9253 VSS.n9243 2.2505
R15702 VSS.n9282 VSS.n9281 2.2505
R15703 VSS.n9207 VSS.n8791 2.2505
R15704 VSS.n9230 VSS.n9229 2.2505
R15705 VSS.n9232 VSS.n8774 2.2505
R15706 VSS.n8797 VSS.n8795 2.2505
R15707 VSS.n9038 VSS.n9037 2.2505
R15708 VSS.n9024 VSS.n8903 2.2505
R15709 VSS.n8890 VSS.n8888 2.2505
R15710 VSS.n8976 VSS.n8975 2.2505
R15711 VSS.n8933 VSS.n8932 2.2505
R15712 VSS.n8969 VSS.n8950 2.2505
R15713 VSS.n10329 VSS.n10328 2.2505
R15714 VSS.n10015 VSS.n10013 2.2505
R15715 VSS.n10322 VSS.n10002 2.2505
R15716 VSS.n10258 VSS.n10257 2.2505
R15717 VSS.n10279 VSS.n10278 2.2505
R15718 VSS.n10251 VSS.n10054 2.2505
R15719 VSS.n10491 VSS.n10490 2.2505
R15720 VSS.n10437 VSS.n10427 2.2505
R15721 VSS.n10466 VSS.n10465 2.2505
R15722 VSS.n10391 VSS.n9975 2.2505
R15723 VSS.n10414 VSS.n10413 2.2505
R15724 VSS.n10416 VSS.n9958 2.2505
R15725 VSS.n9981 VSS.n9979 2.2505
R15726 VSS.n10222 VSS.n10221 2.2505
R15727 VSS.n10208 VSS.n10087 2.2505
R15728 VSS.n10074 VSS.n10072 2.2505
R15729 VSS.n10160 VSS.n10159 2.2505
R15730 VSS.n10117 VSS.n10116 2.2505
R15731 VSS.n10153 VSS.n10134 2.2505
R15732 VSS.n10921 VSS.n10920 2.2505
R15733 VSS.n10607 VSS.n10605 2.2505
R15734 VSS.n10914 VSS.n10594 2.2505
R15735 VSS.n10850 VSS.n10849 2.2505
R15736 VSS.n10871 VSS.n10870 2.2505
R15737 VSS.n10843 VSS.n10646 2.2505
R15738 VSS.n11083 VSS.n11082 2.2505
R15739 VSS.n11029 VSS.n11019 2.2505
R15740 VSS.n11058 VSS.n11057 2.2505
R15741 VSS.n10983 VSS.n10567 2.2505
R15742 VSS.n11006 VSS.n11005 2.2505
R15743 VSS.n11008 VSS.n10550 2.2505
R15744 VSS.n10573 VSS.n10571 2.2505
R15745 VSS.n10814 VSS.n10813 2.2505
R15746 VSS.n10800 VSS.n10679 2.2505
R15747 VSS.n10666 VSS.n10664 2.2505
R15748 VSS.n10752 VSS.n10751 2.2505
R15749 VSS.n10709 VSS.n10708 2.2505
R15750 VSS.n10745 VSS.n10726 2.2505
R15751 VSS.n11513 VSS.n11512 2.2505
R15752 VSS.n11199 VSS.n11197 2.2505
R15753 VSS.n11506 VSS.n11186 2.2505
R15754 VSS.n11442 VSS.n11441 2.2505
R15755 VSS.n11463 VSS.n11462 2.2505
R15756 VSS.n11435 VSS.n11238 2.2505
R15757 VSS.n11675 VSS.n11674 2.2505
R15758 VSS.n11621 VSS.n11611 2.2505
R15759 VSS.n11650 VSS.n11649 2.2505
R15760 VSS.n11575 VSS.n11159 2.2505
R15761 VSS.n11598 VSS.n11597 2.2505
R15762 VSS.n11600 VSS.n11142 2.2505
R15763 VSS.n11165 VSS.n11163 2.2505
R15764 VSS.n11406 VSS.n11405 2.2505
R15765 VSS.n11392 VSS.n11271 2.2505
R15766 VSS.n11258 VSS.n11256 2.2505
R15767 VSS.n11344 VSS.n11343 2.2505
R15768 VSS.n11301 VSS.n11300 2.2505
R15769 VSS.n11337 VSS.n11318 2.2505
R15770 VSS.n12105 VSS.n12104 2.2505
R15771 VSS.n11791 VSS.n11789 2.2505
R15772 VSS.n12098 VSS.n11778 2.2505
R15773 VSS.n12034 VSS.n12033 2.2505
R15774 VSS.n12055 VSS.n12054 2.2505
R15775 VSS.n12027 VSS.n11830 2.2505
R15776 VSS.n12267 VSS.n12266 2.2505
R15777 VSS.n12213 VSS.n12203 2.2505
R15778 VSS.n12242 VSS.n12241 2.2505
R15779 VSS.n12167 VSS.n11751 2.2505
R15780 VSS.n12190 VSS.n12189 2.2505
R15781 VSS.n12192 VSS.n11734 2.2505
R15782 VSS.n11757 VSS.n11755 2.2505
R15783 VSS.n11998 VSS.n11997 2.2505
R15784 VSS.n11984 VSS.n11863 2.2505
R15785 VSS.n11850 VSS.n11848 2.2505
R15786 VSS.n11936 VSS.n11935 2.2505
R15787 VSS.n11893 VSS.n11892 2.2505
R15788 VSS.n11929 VSS.n11910 2.2505
R15789 VSS.n12697 VSS.n12696 2.2505
R15790 VSS.n12383 VSS.n12381 2.2505
R15791 VSS.n12690 VSS.n12370 2.2505
R15792 VSS.n12626 VSS.n12625 2.2505
R15793 VSS.n12647 VSS.n12646 2.2505
R15794 VSS.n12619 VSS.n12422 2.2505
R15795 VSS.n12859 VSS.n12858 2.2505
R15796 VSS.n12805 VSS.n12795 2.2505
R15797 VSS.n12834 VSS.n12833 2.2505
R15798 VSS.n12759 VSS.n12343 2.2505
R15799 VSS.n12782 VSS.n12781 2.2505
R15800 VSS.n12784 VSS.n12326 2.2505
R15801 VSS.n12349 VSS.n12347 2.2505
R15802 VSS.n12590 VSS.n12589 2.2505
R15803 VSS.n12576 VSS.n12455 2.2505
R15804 VSS.n12442 VSS.n12440 2.2505
R15805 VSS.n12528 VSS.n12527 2.2505
R15806 VSS.n12485 VSS.n12484 2.2505
R15807 VSS.n12521 VSS.n12502 2.2505
R15808 VSS.n13289 VSS.n13288 2.2505
R15809 VSS.n12975 VSS.n12973 2.2505
R15810 VSS.n13282 VSS.n12962 2.2505
R15811 VSS.n13218 VSS.n13217 2.2505
R15812 VSS.n13239 VSS.n13238 2.2505
R15813 VSS.n13211 VSS.n13014 2.2505
R15814 VSS.n13451 VSS.n13450 2.2505
R15815 VSS.n13397 VSS.n13387 2.2505
R15816 VSS.n13426 VSS.n13425 2.2505
R15817 VSS.n13351 VSS.n12935 2.2505
R15818 VSS.n13374 VSS.n13373 2.2505
R15819 VSS.n13376 VSS.n12918 2.2505
R15820 VSS.n12941 VSS.n12939 2.2505
R15821 VSS.n13182 VSS.n13181 2.2505
R15822 VSS.n13168 VSS.n13047 2.2505
R15823 VSS.n13034 VSS.n13032 2.2505
R15824 VSS.n13120 VSS.n13119 2.2505
R15825 VSS.n13077 VSS.n13076 2.2505
R15826 VSS.n13113 VSS.n13094 2.2505
R15827 VSS.n13881 VSS.n13880 2.2505
R15828 VSS.n13567 VSS.n13565 2.2505
R15829 VSS.n13874 VSS.n13554 2.2505
R15830 VSS.n13810 VSS.n13809 2.2505
R15831 VSS.n13831 VSS.n13830 2.2505
R15832 VSS.n13803 VSS.n13606 2.2505
R15833 VSS.n14043 VSS.n14042 2.2505
R15834 VSS.n13989 VSS.n13979 2.2505
R15835 VSS.n14018 VSS.n14017 2.2505
R15836 VSS.n13943 VSS.n13527 2.2505
R15837 VSS.n13966 VSS.n13965 2.2505
R15838 VSS.n13968 VSS.n13510 2.2505
R15839 VSS.n13533 VSS.n13531 2.2505
R15840 VSS.n13774 VSS.n13773 2.2505
R15841 VSS.n13760 VSS.n13639 2.2505
R15842 VSS.n13626 VSS.n13624 2.2505
R15843 VSS.n13712 VSS.n13711 2.2505
R15844 VSS.n13669 VSS.n13668 2.2505
R15845 VSS.n13705 VSS.n13686 2.2505
R15846 VSS.n14473 VSS.n14472 2.2505
R15847 VSS.n14159 VSS.n14157 2.2505
R15848 VSS.n14466 VSS.n14146 2.2505
R15849 VSS.n14402 VSS.n14401 2.2505
R15850 VSS.n14423 VSS.n14422 2.2505
R15851 VSS.n14395 VSS.n14198 2.2505
R15852 VSS.n14635 VSS.n14634 2.2505
R15853 VSS.n14581 VSS.n14571 2.2505
R15854 VSS.n14610 VSS.n14609 2.2505
R15855 VSS.n14535 VSS.n14119 2.2505
R15856 VSS.n14558 VSS.n14557 2.2505
R15857 VSS.n14560 VSS.n14102 2.2505
R15858 VSS.n14125 VSS.n14123 2.2505
R15859 VSS.n14366 VSS.n14365 2.2505
R15860 VSS.n14352 VSS.n14231 2.2505
R15861 VSS.n14218 VSS.n14216 2.2505
R15862 VSS.n14304 VSS.n14303 2.2505
R15863 VSS.n14261 VSS.n14260 2.2505
R15864 VSS.n14297 VSS.n14278 2.2505
R15865 VSS.n15065 VSS.n15064 2.2505
R15866 VSS.n14751 VSS.n14749 2.2505
R15867 VSS.n15058 VSS.n14738 2.2505
R15868 VSS.n14994 VSS.n14993 2.2505
R15869 VSS.n15015 VSS.n15014 2.2505
R15870 VSS.n14987 VSS.n14790 2.2505
R15871 VSS.n15227 VSS.n15226 2.2505
R15872 VSS.n15173 VSS.n15163 2.2505
R15873 VSS.n15202 VSS.n15201 2.2505
R15874 VSS.n15127 VSS.n14711 2.2505
R15875 VSS.n15150 VSS.n15149 2.2505
R15876 VSS.n15152 VSS.n14694 2.2505
R15877 VSS.n14717 VSS.n14715 2.2505
R15878 VSS.n14958 VSS.n14957 2.2505
R15879 VSS.n14944 VSS.n14823 2.2505
R15880 VSS.n14810 VSS.n14808 2.2505
R15881 VSS.n14896 VSS.n14895 2.2505
R15882 VSS.n14853 VSS.n14852 2.2505
R15883 VSS.n14889 VSS.n14870 2.2505
R15884 VSS.n15657 VSS.n15656 2.2505
R15885 VSS.n15343 VSS.n15341 2.2505
R15886 VSS.n15650 VSS.n15330 2.2505
R15887 VSS.n15586 VSS.n15585 2.2505
R15888 VSS.n15607 VSS.n15606 2.2505
R15889 VSS.n15579 VSS.n15382 2.2505
R15890 VSS.n15819 VSS.n15818 2.2505
R15891 VSS.n15765 VSS.n15755 2.2505
R15892 VSS.n15794 VSS.n15793 2.2505
R15893 VSS.n15719 VSS.n15303 2.2505
R15894 VSS.n15742 VSS.n15741 2.2505
R15895 VSS.n15744 VSS.n15286 2.2505
R15896 VSS.n15309 VSS.n15307 2.2505
R15897 VSS.n15550 VSS.n15549 2.2505
R15898 VSS.n15536 VSS.n15415 2.2505
R15899 VSS.n15402 VSS.n15400 2.2505
R15900 VSS.n15488 VSS.n15487 2.2505
R15901 VSS.n15445 VSS.n15444 2.2505
R15902 VSS.n15481 VSS.n15462 2.2505
R15903 VSS.n6712 VSS.n6710 2.2505
R15904 VSS.n6778 VSS.n6701 2.2505
R15905 VSS.n6708 VSS.n6707 2.2505
R15906 VSS.n6683 VSS.n6681 2.2505
R15907 VSS.n6689 VSS.n6687 2.2505
R15908 VSS.n6744 VSS.n6743 2.2505
R15909 VSS.n6945 VSS.n6908 2.2505
R15910 VSS.n6891 VSS.n6889 2.2505
R15911 VSS.n15862 VSS.n15861 2.2505
R15912 VSS.n6846 VSS.n6844 2.2505
R15913 VSS.n6876 VSS.n6875 2.2505
R15914 VSS.n6878 VSS.n6868 2.2505
R15915 VSS.n15909 VSS.n15908 2.2505
R15916 VSS.n6658 VSS.n6657 2.2505
R15917 VSS.n6644 VSS.n6523 2.2505
R15918 VSS.n6510 VSS.n6508 2.2505
R15919 VSS.n6596 VSS.n6595 2.2505
R15920 VSS.n6553 VSS.n6552 2.2505
R15921 VSS.n6589 VSS.n6570 2.2505
R15922 VSS.n7369 VSS.n7368 2.2505
R15923 VSS.n7054 VSS.n7052 2.2505
R15924 VSS.n7362 VSS.n7041 2.2505
R15925 VSS.n7298 VSS.n7297 2.2505
R15926 VSS.n7319 VSS.n7318 2.2505
R15927 VSS.n7291 VSS.n7093 2.2505
R15928 VSS.n7531 VSS.n7530 2.2505
R15929 VSS.n7477 VSS.n7467 2.2505
R15930 VSS.n7506 VSS.n7505 2.2505
R15931 VSS.n7431 VSS.n7014 2.2505
R15932 VSS.n7454 VSS.n7453 2.2505
R15933 VSS.n7456 VSS.n6997 2.2505
R15934 VSS.n7020 VSS.n7018 2.2505
R15935 VSS.n7265 VSS.n7264 2.2505
R15936 VSS.n7129 VSS.n7127 2.2505
R15937 VSS.n7258 VSS.n7116 2.2505
R15938 VSS.n7193 VSS.n7192 2.2505
R15939 VSS.n7214 VSS.n7213 2.2505
R15940 VSS.n7186 VSS.n7168 2.2505
R15941 VSS.n18681 VSS.n18680 2.2505
R15942 VSS.n152 VSS.n150 2.2505
R15943 VSS.n18674 VSS.n139 2.2505
R15944 VSS.n18610 VSS.n18609 2.2505
R15945 VSS.n18631 VSS.n18630 2.2505
R15946 VSS.n18603 VSS.n191 2.2505
R15947 VSS.n18843 VSS.n18842 2.2505
R15948 VSS.n18789 VSS.n18779 2.2505
R15949 VSS.n18818 VSS.n18817 2.2505
R15950 VSS.n18743 VSS.n112 2.2505
R15951 VSS.n18766 VSS.n18765 2.2505
R15952 VSS.n18768 VSS.n95 2.2505
R15953 VSS.n118 VSS.n116 2.2505
R15954 VSS.n413 VSS.n412 2.2505
R15955 VSS.n333 VSS.n316 2.2505
R15956 VSS.n323 VSS.n322 2.2505
R15957 VSS.n297 VSS.n295 2.2505
R15958 VSS.n303 VSS.n301 2.2505
R15959 VSS.n348 VSS.n347 2.2505
R15960 VSS.n532 VSS.n530 2.2505
R15961 VSS.n601 VSS.n521 2.2505
R15962 VSS.n528 VSS.n527 2.2505
R15963 VSS.n503 VSS.n501 2.2505
R15964 VSS.n509 VSS.n507 2.2505
R15965 VSS.n499 VSS.n498 2.2505
R15966 VSS.n823 VSS.n822 2.2505
R15967 VSS.n669 VSS.n667 2.2505
R15968 VSS.n699 VSS.n698 2.2505
R15969 VSS.n714 VSS.n712 2.2505
R15970 VSS.n776 VSS.n775 2.2505
R15971 VSS.n742 VSS.n741 2.2505
R15972 VSS.n701 VSS.n691 2.2505
R15973 VSS.n493 VSS.n491 2.2505
R15974 VSS.n944 VSS.n482 2.2505
R15975 VSS.n489 VSS.n488 2.2505
R15976 VSS.n463 VSS.n461 2.2505
R15977 VSS.n469 VSS.n467 2.2505
R15978 VSS.n912 VSS.n911 2.2505
R15979 VSS.n1427 VSS.n1390 2.2505
R15980 VSS.n1373 VSS.n1371 2.2505
R15981 VSS.n17890 VSS.n17889 2.2505
R15982 VSS.n1328 VSS.n1326 2.2505
R15983 VSS.n1358 VSS.n1357 2.2505
R15984 VSS.n1360 VSS.n1350 2.2505
R15985 VSS.n17937 VSS.n17936 2.2505
R15986 VSS.n18860 VSS.n53 2.24315
R15987 VSS.n15836 VSS.n15244 2.24315
R15988 VSS.n13468 VSS.n12876 2.24315
R15989 VSS.n11100 VSS.n10508 2.24315
R15990 VSS.n8732 VSS.n8140 2.24315
R15991 VSS.n5184 VSS.n5183 2.24315
R15992 VSS.n3407 VSS.n1438 2.24315
R15993 VSS.n17865 VSS.n17273 2.24315
R15994 VSS.n17213 VSS.n17212 2.10336
R15995 VSS.n17805 VSS.n17804 2.10336
R15996 VSS.n18498 VSS.n18358 2.10336
R15997 VSS.n9855 VSS.n9854 2.10336
R15998 VSS.n16798 VSS.n16797 2.10336
R15999 VSS.n16205 VSS.n16204 2.10336
R16000 VSS.n2261 VSS.n2260 2.10336
R16001 VSS.n3346 VSS.n3345 2.10336
R16002 VSS.n3938 VSS.n3937 2.10336
R16003 VSS.n4530 VSS.n4529 2.10336
R16004 VSS.n5122 VSS.n5121 2.10336
R16005 VSS.n5226 VSS.n5225 2.10336
R16006 VSS.n5799 VSS.n5798 2.10336
R16007 VSS.n6391 VSS.n6390 2.10336
R16008 VSS.n8079 VSS.n8078 2.10336
R16009 VSS.n8671 VSS.n8670 2.10336
R16010 VSS.n9263 VSS.n9262 2.10336
R16011 VSS.n10447 VSS.n10446 2.10336
R16012 VSS.n11039 VSS.n11038 2.10336
R16013 VSS.n11631 VSS.n11630 2.10336
R16014 VSS.n12223 VSS.n12222 2.10336
R16015 VSS.n12815 VSS.n12814 2.10336
R16016 VSS.n13407 VSS.n13406 2.10336
R16017 VSS.n13999 VSS.n13998 2.10336
R16018 VSS.n14591 VSS.n14590 2.10336
R16019 VSS.n15183 VSS.n15182 2.10336
R16020 VSS.n15775 VSS.n15774 2.10336
R16021 VSS.n15879 VSS.n15878 2.10336
R16022 VSS.n7487 VSS.n7486 2.10336
R16023 VSS.n18799 VSS.n18798 2.10336
R16024 VSS.n793 VSS.n792 2.10336
R16025 VSS.n17907 VSS.n17906 2.10336
R16026 VSS.n17213 VSS.n16895 2.01193
R16027 VSS.n17805 VSS.n17309 2.01193
R16028 VSS.n18499 VSS.n18498 2.01193
R16029 VSS.n9855 VSS.n9359 2.01193
R16030 VSS.n16798 VSS.n16301 2.01193
R16031 VSS.n16205 VSS.n1473 2.01193
R16032 VSS.n2261 VSS.n2125 2.01193
R16033 VSS.n3346 VSS.n2850 2.01193
R16034 VSS.n3938 VSS.n3442 2.01193
R16035 VSS.n4530 VSS.n4034 2.01193
R16036 VSS.n5122 VSS.n4626 2.01193
R16037 VSS.n5226 VSS.n2721 2.01193
R16038 VSS.n5799 VSS.n5682 2.01193
R16039 VSS.n6391 VSS.n6255 2.01193
R16040 VSS.n8079 VSS.n7583 2.01193
R16041 VSS.n8671 VSS.n8175 2.01193
R16042 VSS.n9263 VSS.n8767 2.01193
R16043 VSS.n10447 VSS.n9951 2.01193
R16044 VSS.n11039 VSS.n10543 2.01193
R16045 VSS.n11631 VSS.n11135 2.01193
R16046 VSS.n12223 VSS.n11727 2.01193
R16047 VSS.n12815 VSS.n12319 2.01193
R16048 VSS.n13407 VSS.n12911 2.01193
R16049 VSS.n13999 VSS.n13503 2.01193
R16050 VSS.n14591 VSS.n14095 2.01193
R16051 VSS.n15183 VSS.n14687 2.01193
R16052 VSS.n15775 VSS.n15279 2.01193
R16053 VSS.n15879 VSS.n6861 2.01193
R16054 VSS.n7487 VSS.n6990 2.01193
R16055 VSS.n18799 VSS.n88 2.01193
R16056 VSS.n793 VSS.n684 2.01193
R16057 VSS.n17907 VSS.n1343 2.01193
R16058 VSS.n17993 VSS.n17992 1.98071
R16059 VSS.n1016 VSS.n1015 1.98071
R16060 VSS.n17010 VSS.n17006 1.98071
R16061 VSS.n18042 VSS.n18041 1.98071
R16062 VSS.n17602 VSS.n17420 1.98071
R16063 VSS.n17504 VSS.n17501 1.98071
R16064 VSS.n18081 VSS.n18078 1.98071
R16065 VSS.n18582 VSS.n18581 1.98071
R16066 VSS.n9554 VSS.n9551 1.98071
R16067 VSS.n9652 VSS.n9470 1.98071
R16068 VSS.n16490 VSS.n16487 1.98071
R16069 VSS.n16595 VSS.n16412 1.98071
R16070 VSS.n1655 VSS.n1652 1.98071
R16071 VSS.n16002 VSS.n1577 1.98071
R16072 VSS.n1846 VSS.n1843 1.98071
R16073 VSS.n2347 VSS.n2346 1.98071
R16074 VSS.n3045 VSS.n3042 1.98071
R16075 VSS.n3143 VSS.n2961 1.98071
R16076 VSS.n3637 VSS.n3634 1.98071
R16077 VSS.n3735 VSS.n3553 1.98071
R16078 VSS.n4229 VSS.n4226 1.98071
R16079 VSS.n4327 VSS.n4145 1.98071
R16080 VSS.n4821 VSS.n4818 1.98071
R16081 VSS.n4919 VSS.n4737 1.98071
R16082 VSS.n2442 VSS.n2439 1.98071
R16083 VSS.n5312 VSS.n5311 1.98071
R16084 VSS.n5403 VSS.n5400 1.98071
R16085 VSS.n5885 VSS.n5884 1.98071
R16086 VSS.n5976 VSS.n5973 1.98071
R16087 VSS.n6477 VSS.n6476 1.98071
R16088 VSS.n7778 VSS.n7775 1.98071
R16089 VSS.n7876 VSS.n7694 1.98071
R16090 VSS.n8370 VSS.n8367 1.98071
R16091 VSS.n8468 VSS.n8286 1.98071
R16092 VSS.n8962 VSS.n8959 1.98071
R16093 VSS.n9060 VSS.n8878 1.98071
R16094 VSS.n10146 VSS.n10143 1.98071
R16095 VSS.n10244 VSS.n10062 1.98071
R16096 VSS.n10738 VSS.n10735 1.98071
R16097 VSS.n10836 VSS.n10654 1.98071
R16098 VSS.n11330 VSS.n11327 1.98071
R16099 VSS.n11428 VSS.n11246 1.98071
R16100 VSS.n11922 VSS.n11919 1.98071
R16101 VSS.n12020 VSS.n11838 1.98071
R16102 VSS.n12514 VSS.n12511 1.98071
R16103 VSS.n12612 VSS.n12430 1.98071
R16104 VSS.n13106 VSS.n13103 1.98071
R16105 VSS.n13204 VSS.n13022 1.98071
R16106 VSS.n13698 VSS.n13695 1.98071
R16107 VSS.n13796 VSS.n13614 1.98071
R16108 VSS.n14290 VSS.n14287 1.98071
R16109 VSS.n14388 VSS.n14206 1.98071
R16110 VSS.n14882 VSS.n14879 1.98071
R16111 VSS.n14980 VSS.n14798 1.98071
R16112 VSS.n15474 VSS.n15471 1.98071
R16113 VSS.n15572 VSS.n15390 1.98071
R16114 VSS.n6582 VSS.n6579 1.98071
R16115 VSS.n15965 VSS.n15964 1.98071
R16116 VSS.n7179 VSS.n7176 1.98071
R16117 VSS.n7284 VSS.n7101 1.98071
R16118 VSS.n451 VSS.n450 1.98071
R16119 VSS.n18596 VSS.n192 1.98071
R16120 VSS.n877 VSS.n497 1.98071
R16121 VSS.n17178 VSS.n16905 1.94045
R16122 VSS.n17770 VSS.n17319 1.94045
R16123 VSS.n18506 VSS.n18505 1.94045
R16124 VSS.n9820 VSS.n9369 1.94045
R16125 VSS.n16763 VSS.n16311 1.94045
R16126 VSS.n16170 VSS.n1483 1.94045
R16127 VSS.n2138 VSS.n2134 1.94045
R16128 VSS.n3311 VSS.n2860 1.94045
R16129 VSS.n3903 VSS.n3452 1.94045
R16130 VSS.n4495 VSS.n4044 1.94045
R16131 VSS.n5087 VSS.n4636 1.94045
R16132 VSS.n2734 VSS.n2730 1.94045
R16133 VSS.n5695 VSS.n5691 1.94045
R16134 VSS.n6268 VSS.n6264 1.94045
R16135 VSS.n8044 VSS.n7593 1.94045
R16136 VSS.n8636 VSS.n8185 1.94045
R16137 VSS.n9228 VSS.n8777 1.94045
R16138 VSS.n10412 VSS.n9961 1.94045
R16139 VSS.n11004 VSS.n10553 1.94045
R16140 VSS.n11596 VSS.n11145 1.94045
R16141 VSS.n12188 VSS.n11737 1.94045
R16142 VSS.n12780 VSS.n12329 1.94045
R16143 VSS.n13372 VSS.n12921 1.94045
R16144 VSS.n13964 VSS.n13513 1.94045
R16145 VSS.n14556 VSS.n14105 1.94045
R16146 VSS.n15148 VSS.n14697 1.94045
R16147 VSS.n15740 VSS.n15289 1.94045
R16148 VSS.n6874 VSS.n6870 1.94045
R16149 VSS.n7452 VSS.n7000 1.94045
R16150 VSS.n18764 VSS.n98 1.94045
R16151 VSS.n697 VSS.n693 1.94045
R16152 VSS.n1356 VSS.n1352 1.94045
R16153 VSS VSS.n14060 1.86079
R16154 VSS VSS.n3999 1.86079
R16155 VSS VSS.n18860 1.85712
R16156 VSS VSS.n15836 1.85712
R16157 VSS VSS.n13468 1.85712
R16158 VSS VSS.n11100 1.85712
R16159 VSS VSS.n8732 1.85712
R16160 VSS.n5184 VSS 1.85712
R16161 VSS VSS.n3407 1.85712
R16162 VSS.n17273 VSS 1.85712
R16163 VSS VSS.n9324 1.71006
R16164 VSS.n15837 VSS 1.563
R16165 VSS VSS.n11692 1.563
R16166 VSS VSS.n18889 1.563
R16167 VSS.n16859 VSS 1.563
R16168 VSS.n1234 VSS.n1222 1.55479
R16169 VSS.n1101 VSS.n1089 1.55479
R16170 VSS.n17026 VSS.n16990 1.55479
R16171 VSS.n17520 VSS.n17483 1.55479
R16172 VSS.n17618 VSS.n17404 1.55479
R16173 VSS.n18251 VSS.n18239 1.55479
R16174 VSS.n18097 VSS.n275 1.55479
R16175 VSS.n9668 VSS.n9454 1.55479
R16176 VSS.n9570 VSS.n9533 1.55479
R16177 VSS.n16611 VSS.n16396 1.55479
R16178 VSS.n16506 VSS.n16471 1.55479
R16179 VSS.n16018 VSS.n1568 1.55479
R16180 VSS.n1671 VSS.n1636 1.55479
R16181 VSS.n2016 VSS.n2004 1.55479
R16182 VSS.n1862 VSS.n1825 1.55479
R16183 VSS.n3159 VSS.n2945 1.55479
R16184 VSS.n3061 VSS.n3024 1.55479
R16185 VSS.n3751 VSS.n3537 1.55479
R16186 VSS.n3653 VSS.n3616 1.55479
R16187 VSS.n4343 VSS.n4129 1.55479
R16188 VSS.n4245 VSS.n4208 1.55479
R16189 VSS.n4935 VSS.n4721 1.55479
R16190 VSS.n4837 VSS.n4800 1.55479
R16191 VSS.n2612 VSS.n2600 1.55479
R16192 VSS.n2458 VSS.n2421 1.55479
R16193 VSS.n5573 VSS.n5561 1.55479
R16194 VSS.n5419 VSS.n5382 1.55479
R16195 VSS.n6146 VSS.n6134 1.55479
R16196 VSS.n5992 VSS.n5955 1.55479
R16197 VSS.n7892 VSS.n7678 1.55479
R16198 VSS.n7794 VSS.n7757 1.55479
R16199 VSS.n8484 VSS.n8270 1.55479
R16200 VSS.n8386 VSS.n8349 1.55479
R16201 VSS.n9076 VSS.n8862 1.55479
R16202 VSS.n8978 VSS.n8941 1.55479
R16203 VSS.n10260 VSS.n10046 1.55479
R16204 VSS.n10162 VSS.n10125 1.55479
R16205 VSS.n10852 VSS.n10638 1.55479
R16206 VSS.n10754 VSS.n10717 1.55479
R16207 VSS.n11444 VSS.n11230 1.55479
R16208 VSS.n11346 VSS.n11309 1.55479
R16209 VSS.n12036 VSS.n11822 1.55479
R16210 VSS.n11938 VSS.n11901 1.55479
R16211 VSS.n12628 VSS.n12414 1.55479
R16212 VSS.n12530 VSS.n12493 1.55479
R16213 VSS.n13220 VSS.n13006 1.55479
R16214 VSS.n13122 VSS.n13085 1.55479
R16215 VSS.n13812 VSS.n13598 1.55479
R16216 VSS.n13714 VSS.n13677 1.55479
R16217 VSS.n14404 VSS.n14190 1.55479
R16218 VSS.n14306 VSS.n14269 1.55479
R16219 VSS.n14996 VSS.n14782 1.55479
R16220 VSS.n14898 VSS.n14861 1.55479
R16221 VSS.n15588 VSS.n15374 1.55479
R16222 VSS.n15490 VSS.n15453 1.55479
R16223 VSS.n6752 VSS.n6740 1.55479
R16224 VSS.n6598 VSS.n6561 1.55479
R16225 VSS.n7300 VSS.n7085 1.55479
R16226 VSS.n7195 VSS.n7160 1.55479
R16227 VSS.n18612 VSS.n183 1.55479
R16228 VSS.n356 VSS.n343 1.55479
R16229 VSS.n575 VSS.n565 1.55479
R16230 VSS.n920 VSS.n908 1.55479
R16231 VSS.n17168 VSS.n16914 1.53956
R16232 VSS.n17218 VSS.n16882 1.53956
R16233 VSS.n17760 VSS.n17328 1.53956
R16234 VSS.n17810 VSS.n17296 1.53956
R16235 VSS.n18381 VSS.n18373 1.53956
R16236 VSS.n18493 VSS.n18385 1.53956
R16237 VSS.n9810 VSS.n9378 1.53956
R16238 VSS.n9860 VSS.n9346 1.53956
R16239 VSS.n16753 VSS.n16320 1.53956
R16240 VSS.n16803 VSS.n16288 1.53956
R16241 VSS.n16160 VSS.n1492 1.53956
R16242 VSS.n16210 VSS.n1460 1.53956
R16243 VSS.n2266 VSS.n2106 1.53956
R16244 VSS.n2190 VSS.n2187 1.53956
R16245 VSS.n3301 VSS.n2869 1.53956
R16246 VSS.n3351 VSS.n2837 1.53956
R16247 VSS.n3893 VSS.n3461 1.53956
R16248 VSS.n3943 VSS.n3429 1.53956
R16249 VSS.n4485 VSS.n4053 1.53956
R16250 VSS.n4535 VSS.n4021 1.53956
R16251 VSS.n5077 VSS.n4645 1.53956
R16252 VSS.n5127 VSS.n4613 1.53956
R16253 VSS.n5231 VSS.n2702 1.53956
R16254 VSS.n2786 VSS.n2783 1.53956
R16255 VSS.n5804 VSS.n5663 1.53956
R16256 VSS.n5760 VSS.n5757 1.53956
R16257 VSS.n6396 VSS.n6236 1.53956
R16258 VSS.n6320 VSS.n6317 1.53956
R16259 VSS.n8034 VSS.n7602 1.53956
R16260 VSS.n8084 VSS.n7570 1.53956
R16261 VSS.n8626 VSS.n8194 1.53956
R16262 VSS.n8676 VSS.n8162 1.53956
R16263 VSS.n9218 VSS.n8786 1.53956
R16264 VSS.n9268 VSS.n8754 1.53956
R16265 VSS.n10402 VSS.n9970 1.53956
R16266 VSS.n10452 VSS.n9938 1.53956
R16267 VSS.n10994 VSS.n10562 1.53956
R16268 VSS.n11044 VSS.n10530 1.53956
R16269 VSS.n11586 VSS.n11154 1.53956
R16270 VSS.n11636 VSS.n11122 1.53956
R16271 VSS.n12178 VSS.n11746 1.53956
R16272 VSS.n12228 VSS.n11714 1.53956
R16273 VSS.n12770 VSS.n12338 1.53956
R16274 VSS.n12820 VSS.n12306 1.53956
R16275 VSS.n13362 VSS.n12930 1.53956
R16276 VSS.n13412 VSS.n12898 1.53956
R16277 VSS.n13954 VSS.n13522 1.53956
R16278 VSS.n14004 VSS.n13490 1.53956
R16279 VSS.n14546 VSS.n14114 1.53956
R16280 VSS.n14596 VSS.n14082 1.53956
R16281 VSS.n15138 VSS.n14706 1.53956
R16282 VSS.n15188 VSS.n14674 1.53956
R16283 VSS.n15730 VSS.n15298 1.53956
R16284 VSS.n15780 VSS.n15266 1.53956
R16285 VSS.n15884 VSS.n6842 1.53956
R16286 VSS.n6926 VSS.n6923 1.53956
R16287 VSS.n7442 VSS.n7009 1.53956
R16288 VSS.n7492 VSS.n6977 1.53956
R16289 VSS.n18754 VSS.n107 1.53956
R16290 VSS.n18804 VSS.n75 1.53956
R16291 VSS.n798 VSS.n665 1.53956
R16292 VSS.n757 VSS.n756 1.53956
R16293 VSS.n17912 VSS.n1324 1.53956
R16294 VSS.n1408 VSS.n1405 1.53956
R16295 VSS.n1045 VSS.n1043 1.5005
R16296 VSS.n17553 VSS.n17552 1.5005
R16297 VSS.n18130 VSS.n18129 1.5005
R16298 VSS.n9603 VSS.n9602 1.5005
R16299 VSS.n16452 VSS.n16451 1.5005
R16300 VSS.n1617 VSS.n1616 1.5005
R16301 VSS.n1895 VSS.n1894 1.5005
R16302 VSS.n3094 VSS.n3093 1.5005
R16303 VSS.n3686 VSS.n3685 1.5005
R16304 VSS.n4278 VSS.n4277 1.5005
R16305 VSS.n4870 VSS.n4869 1.5005
R16306 VSS.n2491 VSS.n2490 1.5005
R16307 VSS.n5452 VSS.n5451 1.5005
R16308 VSS.n6025 VSS.n6024 1.5005
R16309 VSS.n7827 VSS.n7826 1.5005
R16310 VSS.n8419 VSS.n8418 1.5005
R16311 VSS.n9011 VSS.n9010 1.5005
R16312 VSS.n10195 VSS.n10194 1.5005
R16313 VSS.n10787 VSS.n10786 1.5005
R16314 VSS.n11379 VSS.n11378 1.5005
R16315 VSS.n11971 VSS.n11970 1.5005
R16316 VSS.n12563 VSS.n12562 1.5005
R16317 VSS.n13155 VSS.n13154 1.5005
R16318 VSS.n13747 VSS.n13746 1.5005
R16319 VSS.n14339 VSS.n14338 1.5005
R16320 VSS.n14931 VSS.n14930 1.5005
R16321 VSS.n15523 VSS.n15522 1.5005
R16322 VSS.n6631 VSS.n6630 1.5005
R16323 VSS.n7141 VSS.n7140 1.5005
R16324 VSS.n312 VSS.n310 1.5005
R16325 VSS.n478 VSS.n476 1.5005
R16326 VSS.n1275 VSS.n1201 1.46336
R16327 VSS.n1141 VSS.n1067 1.46336
R16328 VSS.n16912 VSS.n16904 1.46336
R16329 VSS.n17219 VSS.n16891 1.46336
R16330 VSS.n17085 VSS.n16940 1.46336
R16331 VSS.n17435 VSS.n17429 1.46336
R16332 VSS.n17326 VSS.n17318 1.46336
R16333 VSS.n17811 VSS.n17305 1.46336
R16334 VSS.n17677 VSS.n17354 1.46336
R16335 VSS.n18292 VSS.n18218 1.46336
R16336 VSS.n18380 VSS.n18379 1.46336
R16337 VSS.n18492 VSS.n18386 1.46336
R16338 VSS.n227 VSS.n221 1.46336
R16339 VSS.n9727 VSS.n9404 1.46336
R16340 VSS.n9376 VSS.n9368 1.46336
R16341 VSS.n9861 VSS.n9355 1.46336
R16342 VSS.n9485 VSS.n9479 1.46336
R16343 VSS.n16670 VSS.n16346 1.46336
R16344 VSS.n16318 VSS.n16310 1.46336
R16345 VSS.n16804 VSS.n16297 1.46336
R16346 VSS.n16566 VSS.n16421 1.46336
R16347 VSS.n16077 VSS.n1518 1.46336
R16348 VSS.n1490 VSS.n1482 1.46336
R16349 VSS.n16211 VSS.n1469 1.46336
R16350 VSS.n1731 VSS.n1586 1.46336
R16351 VSS.n2057 VSS.n1983 1.46336
R16352 VSS.n2267 VSS.n2121 1.46336
R16353 VSS.n2186 VSS.n2185 1.46336
R16354 VSS.n1777 VSS.n1771 1.46336
R16355 VSS.n3218 VSS.n2895 1.46336
R16356 VSS.n2867 VSS.n2859 1.46336
R16357 VSS.n3352 VSS.n2846 1.46336
R16358 VSS.n2976 VSS.n2970 1.46336
R16359 VSS.n3810 VSS.n3487 1.46336
R16360 VSS.n3459 VSS.n3451 1.46336
R16361 VSS.n3944 VSS.n3438 1.46336
R16362 VSS.n3568 VSS.n3562 1.46336
R16363 VSS.n4402 VSS.n4079 1.46336
R16364 VSS.n4051 VSS.n4043 1.46336
R16365 VSS.n4536 VSS.n4030 1.46336
R16366 VSS.n4160 VSS.n4154 1.46336
R16367 VSS.n4994 VSS.n4671 1.46336
R16368 VSS.n4643 VSS.n4635 1.46336
R16369 VSS.n5128 VSS.n4622 1.46336
R16370 VSS.n4752 VSS.n4746 1.46336
R16371 VSS.n2653 VSS.n2579 1.46336
R16372 VSS.n5232 VSS.n2717 1.46336
R16373 VSS.n2782 VSS.n2781 1.46336
R16374 VSS.n2373 VSS.n2367 1.46336
R16375 VSS.n5614 VSS.n5540 1.46336
R16376 VSS.n5805 VSS.n5678 1.46336
R16377 VSS.n5756 VSS.n5755 1.46336
R16378 VSS.n5334 VSS.n5328 1.46336
R16379 VSS.n6187 VSS.n6113 1.46336
R16380 VSS.n6397 VSS.n6251 1.46336
R16381 VSS.n6316 VSS.n6315 1.46336
R16382 VSS.n5907 VSS.n5901 1.46336
R16383 VSS.n7951 VSS.n7628 1.46336
R16384 VSS.n7600 VSS.n7592 1.46336
R16385 VSS.n8085 VSS.n7579 1.46336
R16386 VSS.n7709 VSS.n7703 1.46336
R16387 VSS.n8543 VSS.n8220 1.46336
R16388 VSS.n8192 VSS.n8184 1.46336
R16389 VSS.n8677 VSS.n8171 1.46336
R16390 VSS.n8301 VSS.n8295 1.46336
R16391 VSS.n9135 VSS.n8812 1.46336
R16392 VSS.n8784 VSS.n8776 1.46336
R16393 VSS.n9269 VSS.n8763 1.46336
R16394 VSS.n8893 VSS.n8887 1.46336
R16395 VSS.n10319 VSS.n9996 1.46336
R16396 VSS.n9968 VSS.n9960 1.46336
R16397 VSS.n10453 VSS.n9947 1.46336
R16398 VSS.n10077 VSS.n10071 1.46336
R16399 VSS.n10911 VSS.n10588 1.46336
R16400 VSS.n10560 VSS.n10552 1.46336
R16401 VSS.n11045 VSS.n10539 1.46336
R16402 VSS.n10669 VSS.n10663 1.46336
R16403 VSS.n11503 VSS.n11180 1.46336
R16404 VSS.n11152 VSS.n11144 1.46336
R16405 VSS.n11637 VSS.n11131 1.46336
R16406 VSS.n11261 VSS.n11255 1.46336
R16407 VSS.n12095 VSS.n11772 1.46336
R16408 VSS.n11744 VSS.n11736 1.46336
R16409 VSS.n12229 VSS.n11723 1.46336
R16410 VSS.n11853 VSS.n11847 1.46336
R16411 VSS.n12687 VSS.n12364 1.46336
R16412 VSS.n12336 VSS.n12328 1.46336
R16413 VSS.n12821 VSS.n12315 1.46336
R16414 VSS.n12445 VSS.n12439 1.46336
R16415 VSS.n13279 VSS.n12956 1.46336
R16416 VSS.n12928 VSS.n12920 1.46336
R16417 VSS.n13413 VSS.n12907 1.46336
R16418 VSS.n13037 VSS.n13031 1.46336
R16419 VSS.n13871 VSS.n13548 1.46336
R16420 VSS.n13520 VSS.n13512 1.46336
R16421 VSS.n14005 VSS.n13499 1.46336
R16422 VSS.n13629 VSS.n13623 1.46336
R16423 VSS.n14463 VSS.n14140 1.46336
R16424 VSS.n14112 VSS.n14104 1.46336
R16425 VSS.n14597 VSS.n14091 1.46336
R16426 VSS.n14221 VSS.n14215 1.46336
R16427 VSS.n15055 VSS.n14732 1.46336
R16428 VSS.n14704 VSS.n14696 1.46336
R16429 VSS.n15189 VSS.n14683 1.46336
R16430 VSS.n14813 VSS.n14807 1.46336
R16431 VSS.n15647 VSS.n15324 1.46336
R16432 VSS.n15296 VSS.n15288 1.46336
R16433 VSS.n15781 VSS.n15275 1.46336
R16434 VSS.n15405 VSS.n15399 1.46336
R16435 VSS.n6793 VSS.n6719 1.46336
R16436 VSS.n15885 VSS.n6857 1.46336
R16437 VSS.n6922 VSS.n6921 1.46336
R16438 VSS.n6513 VSS.n6507 1.46336
R16439 VSS.n7359 VSS.n7035 1.46336
R16440 VSS.n7007 VSS.n6999 1.46336
R16441 VSS.n7493 VSS.n6986 1.46336
R16442 VSS.n7255 VSS.n7110 1.46336
R16443 VSS.n18671 VSS.n133 1.46336
R16444 VSS.n105 VSS.n97 1.46336
R16445 VSS.n18805 VSS.n84 1.46336
R16446 VSS.n405 VSS.n328 1.46336
R16447 VSS.n616 VSS.n539 1.46336
R16448 VSS.n799 VSS.n680 1.46336
R16449 VSS.n754 VSS.n753 1.46336
R16450 VSS.n960 VSS.n886 1.46336
R16451 VSS.n17913 VSS.n1339 1.46336
R16452 VSS.n1404 VSS.n1403 1.46336
R16453 VSS.n1241 VSS.n1214 1.37193
R16454 VSS.n1251 VSS.n1250 1.37193
R16455 VSS.n1258 VSS.n1257 1.37193
R16456 VSS.n1261 VSS.n1259 1.37193
R16457 VSS.n1106 VSS.n1081 1.37193
R16458 VSS.n1116 VSS.n1115 1.37193
R16459 VSS.n1123 VSS.n1122 1.37193
R16460 VSS.n1126 VSS.n1124 1.37193
R16461 VSS.n17033 VSS.n16976 1.37193
R16462 VSS.n17048 VSS.n16970 1.37193
R16463 VSS.n16971 VSS.n16955 1.37193
R16464 VSS.n17071 VSS.n16956 1.37193
R16465 VSS.n17532 VSS.n17477 1.37193
R16466 VSS.n17478 VSS.n17460 1.37193
R16467 VSS.n17556 VSS.n17448 1.37193
R16468 VSS.n17455 VSS.n17449 1.37193
R16469 VSS.n17625 VSS.n17390 1.37193
R16470 VSS.n17640 VSS.n17384 1.37193
R16471 VSS.n17385 VSS.n17369 1.37193
R16472 VSS.n17663 VSS.n17370 1.37193
R16473 VSS.n18258 VSS.n18231 1.37193
R16474 VSS.n18268 VSS.n18267 1.37193
R16475 VSS.n18275 VSS.n18274 1.37193
R16476 VSS.n18278 VSS.n18276 1.37193
R16477 VSS.n18109 VSS.n269 1.37193
R16478 VSS.n270 VSS.n252 1.37193
R16479 VSS.n18133 VSS.n240 1.37193
R16480 VSS.n247 VSS.n241 1.37193
R16481 VSS.n9675 VSS.n9440 1.37193
R16482 VSS.n9690 VSS.n9434 1.37193
R16483 VSS.n9435 VSS.n9419 1.37193
R16484 VSS.n9713 VSS.n9420 1.37193
R16485 VSS.n9582 VSS.n9527 1.37193
R16486 VSS.n9528 VSS.n9510 1.37193
R16487 VSS.n9606 VSS.n9498 1.37193
R16488 VSS.n9505 VSS.n9499 1.37193
R16489 VSS.n16618 VSS.n16382 1.37193
R16490 VSS.n16633 VSS.n16376 1.37193
R16491 VSS.n16377 VSS.n16361 1.37193
R16492 VSS.n16656 VSS.n16362 1.37193
R16493 VSS.n16513 VSS.n16459 1.37193
R16494 VSS.n16528 VSS.n16453 1.37193
R16495 VSS.n16454 VSS.n16436 1.37193
R16496 VSS.n16551 VSS.n16437 1.37193
R16497 VSS.n16025 VSS.n1554 1.37193
R16498 VSS.n16040 VSS.n1548 1.37193
R16499 VSS.n1549 VSS.n1533 1.37193
R16500 VSS.n16063 VSS.n1534 1.37193
R16501 VSS.n1678 VSS.n1624 1.37193
R16502 VSS.n1693 VSS.n1618 1.37193
R16503 VSS.n1619 VSS.n1601 1.37193
R16504 VSS.n1716 VSS.n1602 1.37193
R16505 VSS.n2023 VSS.n1996 1.37193
R16506 VSS.n2033 VSS.n2032 1.37193
R16507 VSS.n2040 VSS.n2039 1.37193
R16508 VSS.n2043 VSS.n2041 1.37193
R16509 VSS.n1874 VSS.n1819 1.37193
R16510 VSS.n1820 VSS.n1802 1.37193
R16511 VSS.n1898 VSS.n1790 1.37193
R16512 VSS.n1797 VSS.n1791 1.37193
R16513 VSS.n3166 VSS.n2931 1.37193
R16514 VSS.n3181 VSS.n2925 1.37193
R16515 VSS.n2926 VSS.n2910 1.37193
R16516 VSS.n3204 VSS.n2911 1.37193
R16517 VSS.n3073 VSS.n3018 1.37193
R16518 VSS.n3019 VSS.n3001 1.37193
R16519 VSS.n3097 VSS.n2989 1.37193
R16520 VSS.n2996 VSS.n2990 1.37193
R16521 VSS.n3758 VSS.n3523 1.37193
R16522 VSS.n3773 VSS.n3517 1.37193
R16523 VSS.n3518 VSS.n3502 1.37193
R16524 VSS.n3796 VSS.n3503 1.37193
R16525 VSS.n3665 VSS.n3610 1.37193
R16526 VSS.n3611 VSS.n3593 1.37193
R16527 VSS.n3689 VSS.n3581 1.37193
R16528 VSS.n3588 VSS.n3582 1.37193
R16529 VSS.n4350 VSS.n4115 1.37193
R16530 VSS.n4365 VSS.n4109 1.37193
R16531 VSS.n4110 VSS.n4094 1.37193
R16532 VSS.n4388 VSS.n4095 1.37193
R16533 VSS.n4257 VSS.n4202 1.37193
R16534 VSS.n4203 VSS.n4185 1.37193
R16535 VSS.n4281 VSS.n4173 1.37193
R16536 VSS.n4180 VSS.n4174 1.37193
R16537 VSS.n4942 VSS.n4707 1.37193
R16538 VSS.n4957 VSS.n4701 1.37193
R16539 VSS.n4702 VSS.n4686 1.37193
R16540 VSS.n4980 VSS.n4687 1.37193
R16541 VSS.n4849 VSS.n4794 1.37193
R16542 VSS.n4795 VSS.n4777 1.37193
R16543 VSS.n4873 VSS.n4765 1.37193
R16544 VSS.n4772 VSS.n4766 1.37193
R16545 VSS.n2619 VSS.n2592 1.37193
R16546 VSS.n2629 VSS.n2628 1.37193
R16547 VSS.n2636 VSS.n2635 1.37193
R16548 VSS.n2639 VSS.n2637 1.37193
R16549 VSS.n2470 VSS.n2415 1.37193
R16550 VSS.n2416 VSS.n2398 1.37193
R16551 VSS.n2494 VSS.n2386 1.37193
R16552 VSS.n2393 VSS.n2387 1.37193
R16553 VSS.n5580 VSS.n5553 1.37193
R16554 VSS.n5590 VSS.n5589 1.37193
R16555 VSS.n5597 VSS.n5596 1.37193
R16556 VSS.n5600 VSS.n5598 1.37193
R16557 VSS.n5431 VSS.n5376 1.37193
R16558 VSS.n5377 VSS.n5359 1.37193
R16559 VSS.n5455 VSS.n5347 1.37193
R16560 VSS.n5354 VSS.n5348 1.37193
R16561 VSS.n6153 VSS.n6126 1.37193
R16562 VSS.n6163 VSS.n6162 1.37193
R16563 VSS.n6170 VSS.n6169 1.37193
R16564 VSS.n6173 VSS.n6171 1.37193
R16565 VSS.n6004 VSS.n5949 1.37193
R16566 VSS.n5950 VSS.n5932 1.37193
R16567 VSS.n6028 VSS.n5920 1.37193
R16568 VSS.n5927 VSS.n5921 1.37193
R16569 VSS.n7899 VSS.n7664 1.37193
R16570 VSS.n7914 VSS.n7658 1.37193
R16571 VSS.n7659 VSS.n7643 1.37193
R16572 VSS.n7937 VSS.n7644 1.37193
R16573 VSS.n7806 VSS.n7751 1.37193
R16574 VSS.n7752 VSS.n7734 1.37193
R16575 VSS.n7830 VSS.n7722 1.37193
R16576 VSS.n7729 VSS.n7723 1.37193
R16577 VSS.n8491 VSS.n8256 1.37193
R16578 VSS.n8506 VSS.n8250 1.37193
R16579 VSS.n8251 VSS.n8235 1.37193
R16580 VSS.n8529 VSS.n8236 1.37193
R16581 VSS.n8398 VSS.n8343 1.37193
R16582 VSS.n8344 VSS.n8326 1.37193
R16583 VSS.n8422 VSS.n8314 1.37193
R16584 VSS.n8321 VSS.n8315 1.37193
R16585 VSS.n9083 VSS.n8848 1.37193
R16586 VSS.n9098 VSS.n8842 1.37193
R16587 VSS.n8843 VSS.n8827 1.37193
R16588 VSS.n9121 VSS.n8828 1.37193
R16589 VSS.n8990 VSS.n8935 1.37193
R16590 VSS.n8936 VSS.n8918 1.37193
R16591 VSS.n9014 VSS.n8906 1.37193
R16592 VSS.n8913 VSS.n8907 1.37193
R16593 VSS.n10267 VSS.n10032 1.37193
R16594 VSS.n10282 VSS.n10026 1.37193
R16595 VSS.n10027 VSS.n10011 1.37193
R16596 VSS.n10305 VSS.n10012 1.37193
R16597 VSS.n10174 VSS.n10119 1.37193
R16598 VSS.n10120 VSS.n10102 1.37193
R16599 VSS.n10198 VSS.n10090 1.37193
R16600 VSS.n10097 VSS.n10091 1.37193
R16601 VSS.n10859 VSS.n10624 1.37193
R16602 VSS.n10874 VSS.n10618 1.37193
R16603 VSS.n10619 VSS.n10603 1.37193
R16604 VSS.n10897 VSS.n10604 1.37193
R16605 VSS.n10766 VSS.n10711 1.37193
R16606 VSS.n10712 VSS.n10694 1.37193
R16607 VSS.n10790 VSS.n10682 1.37193
R16608 VSS.n10689 VSS.n10683 1.37193
R16609 VSS.n11451 VSS.n11216 1.37193
R16610 VSS.n11466 VSS.n11210 1.37193
R16611 VSS.n11211 VSS.n11195 1.37193
R16612 VSS.n11489 VSS.n11196 1.37193
R16613 VSS.n11358 VSS.n11303 1.37193
R16614 VSS.n11304 VSS.n11286 1.37193
R16615 VSS.n11382 VSS.n11274 1.37193
R16616 VSS.n11281 VSS.n11275 1.37193
R16617 VSS.n12043 VSS.n11808 1.37193
R16618 VSS.n12058 VSS.n11802 1.37193
R16619 VSS.n11803 VSS.n11787 1.37193
R16620 VSS.n12081 VSS.n11788 1.37193
R16621 VSS.n11950 VSS.n11895 1.37193
R16622 VSS.n11896 VSS.n11878 1.37193
R16623 VSS.n11974 VSS.n11866 1.37193
R16624 VSS.n11873 VSS.n11867 1.37193
R16625 VSS.n12635 VSS.n12400 1.37193
R16626 VSS.n12650 VSS.n12394 1.37193
R16627 VSS.n12395 VSS.n12379 1.37193
R16628 VSS.n12673 VSS.n12380 1.37193
R16629 VSS.n12542 VSS.n12487 1.37193
R16630 VSS.n12488 VSS.n12470 1.37193
R16631 VSS.n12566 VSS.n12458 1.37193
R16632 VSS.n12465 VSS.n12459 1.37193
R16633 VSS.n13227 VSS.n12992 1.37193
R16634 VSS.n13242 VSS.n12986 1.37193
R16635 VSS.n12987 VSS.n12971 1.37193
R16636 VSS.n13265 VSS.n12972 1.37193
R16637 VSS.n13134 VSS.n13079 1.37193
R16638 VSS.n13080 VSS.n13062 1.37193
R16639 VSS.n13158 VSS.n13050 1.37193
R16640 VSS.n13057 VSS.n13051 1.37193
R16641 VSS.n13819 VSS.n13584 1.37193
R16642 VSS.n13834 VSS.n13578 1.37193
R16643 VSS.n13579 VSS.n13563 1.37193
R16644 VSS.n13857 VSS.n13564 1.37193
R16645 VSS.n13726 VSS.n13671 1.37193
R16646 VSS.n13672 VSS.n13654 1.37193
R16647 VSS.n13750 VSS.n13642 1.37193
R16648 VSS.n13649 VSS.n13643 1.37193
R16649 VSS.n14411 VSS.n14176 1.37193
R16650 VSS.n14426 VSS.n14170 1.37193
R16651 VSS.n14171 VSS.n14155 1.37193
R16652 VSS.n14449 VSS.n14156 1.37193
R16653 VSS.n14318 VSS.n14263 1.37193
R16654 VSS.n14264 VSS.n14246 1.37193
R16655 VSS.n14342 VSS.n14234 1.37193
R16656 VSS.n14241 VSS.n14235 1.37193
R16657 VSS.n15003 VSS.n14768 1.37193
R16658 VSS.n15018 VSS.n14762 1.37193
R16659 VSS.n14763 VSS.n14747 1.37193
R16660 VSS.n15041 VSS.n14748 1.37193
R16661 VSS.n14910 VSS.n14855 1.37193
R16662 VSS.n14856 VSS.n14838 1.37193
R16663 VSS.n14934 VSS.n14826 1.37193
R16664 VSS.n14833 VSS.n14827 1.37193
R16665 VSS.n15595 VSS.n15360 1.37193
R16666 VSS.n15610 VSS.n15354 1.37193
R16667 VSS.n15355 VSS.n15339 1.37193
R16668 VSS.n15633 VSS.n15340 1.37193
R16669 VSS.n15502 VSS.n15447 1.37193
R16670 VSS.n15448 VSS.n15430 1.37193
R16671 VSS.n15526 VSS.n15418 1.37193
R16672 VSS.n15425 VSS.n15419 1.37193
R16673 VSS.n6759 VSS.n6732 1.37193
R16674 VSS.n6769 VSS.n6768 1.37193
R16675 VSS.n6776 VSS.n6775 1.37193
R16676 VSS.n6779 VSS.n6777 1.37193
R16677 VSS.n6610 VSS.n6555 1.37193
R16678 VSS.n6556 VSS.n6538 1.37193
R16679 VSS.n6634 VSS.n6526 1.37193
R16680 VSS.n6533 VSS.n6527 1.37193
R16681 VSS.n7307 VSS.n7071 1.37193
R16682 VSS.n7322 VSS.n7065 1.37193
R16683 VSS.n7066 VSS.n7050 1.37193
R16684 VSS.n7345 VSS.n7051 1.37193
R16685 VSS.n7202 VSS.n7148 1.37193
R16686 VSS.n7217 VSS.n7142 1.37193
R16687 VSS.n7143 VSS.n7125 1.37193
R16688 VSS.n7240 VSS.n7126 1.37193
R16689 VSS.n18619 VSS.n169 1.37193
R16690 VSS.n18634 VSS.n163 1.37193
R16691 VSS.n164 VSS.n148 1.37193
R16692 VSS.n18657 VSS.n149 1.37193
R16693 VSS.n365 VSS.n342 1.37193
R16694 VSS.n377 VSS.n338 1.37193
R16695 VSS.n380 VSS.n334 1.37193
R16696 VSS.n393 VSS.n332 1.37193
R16697 VSS.n582 VSS.n552 1.37193
R16698 VSS.n592 VSS.n591 1.37193
R16699 VSS.n599 VSS.n598 1.37193
R16700 VSS.n602 VSS.n600 1.37193
R16701 VSS.n925 VSS.n900 1.37193
R16702 VSS.n935 VSS.n934 1.37193
R16703 VSS.n942 VSS.n941 1.37193
R16704 VSS.n945 VSS.n943 1.37193
R16705 VSS.n17162 VSS.n17161 1.2805
R16706 VSS.n17234 VSS.n16879 1.2805
R16707 VSS.n17754 VSS.n17753 1.2805
R16708 VSS.n17826 VSS.n17293 1.2805
R16709 VSS.n18366 VSS.n18343 1.2805
R16710 VSS.n18448 VSS.n18442 1.2805
R16711 VSS.n9804 VSS.n9803 1.2805
R16712 VSS.n9876 VSS.n9343 1.2805
R16713 VSS.n16747 VSS.n16746 1.2805
R16714 VSS.n16819 VSS.n16285 1.2805
R16715 VSS.n16154 VSS.n16153 1.2805
R16716 VSS.n16226 VSS.n1457 1.2805
R16717 VSS.n2277 VSS.n2103 1.2805
R16718 VSS.n2194 VSS.n2158 1.2805
R16719 VSS.n3295 VSS.n3294 1.2805
R16720 VSS.n3367 VSS.n2834 1.2805
R16721 VSS.n3887 VSS.n3886 1.2805
R16722 VSS.n3959 VSS.n3426 1.2805
R16723 VSS.n4479 VSS.n4478 1.2805
R16724 VSS.n4551 VSS.n4018 1.2805
R16725 VSS.n5071 VSS.n5070 1.2805
R16726 VSS.n5143 VSS.n4610 1.2805
R16727 VSS.n5242 VSS.n2699 1.2805
R16728 VSS.n2790 VSS.n2754 1.2805
R16729 VSS.n5815 VSS.n5660 1.2805
R16730 VSS.n5764 VSS.n5715 1.2805
R16731 VSS.n6407 VSS.n6233 1.2805
R16732 VSS.n6324 VSS.n6288 1.2805
R16733 VSS.n8028 VSS.n8027 1.2805
R16734 VSS.n8100 VSS.n7567 1.2805
R16735 VSS.n8620 VSS.n8619 1.2805
R16736 VSS.n8692 VSS.n8159 1.2805
R16737 VSS.n9212 VSS.n9211 1.2805
R16738 VSS.n9284 VSS.n8751 1.2805
R16739 VSS.n10396 VSS.n10395 1.2805
R16740 VSS.n10468 VSS.n9935 1.2805
R16741 VSS.n10988 VSS.n10987 1.2805
R16742 VSS.n11060 VSS.n10527 1.2805
R16743 VSS.n11580 VSS.n11579 1.2805
R16744 VSS.n11652 VSS.n11119 1.2805
R16745 VSS.n12172 VSS.n12171 1.2805
R16746 VSS.n12244 VSS.n11711 1.2805
R16747 VSS.n12764 VSS.n12763 1.2805
R16748 VSS.n12836 VSS.n12303 1.2805
R16749 VSS.n13356 VSS.n13355 1.2805
R16750 VSS.n13428 VSS.n12895 1.2805
R16751 VSS.n13948 VSS.n13947 1.2805
R16752 VSS.n14020 VSS.n13487 1.2805
R16753 VSS.n14540 VSS.n14539 1.2805
R16754 VSS.n14612 VSS.n14079 1.2805
R16755 VSS.n15132 VSS.n15131 1.2805
R16756 VSS.n15204 VSS.n14671 1.2805
R16757 VSS.n15724 VSS.n15723 1.2805
R16758 VSS.n15796 VSS.n15263 1.2805
R16759 VSS.n15895 VSS.n6839 1.2805
R16760 VSS.n6930 VSS.n6894 1.2805
R16761 VSS.n7436 VSS.n7435 1.2805
R16762 VSS.n7508 VSS.n6974 1.2805
R16763 VSS.n18748 VSS.n18747 1.2805
R16764 VSS.n18820 VSS.n72 1.2805
R16765 VSS.n809 VSS.n662 1.2805
R16766 VSS.n743 VSS.n717 1.2805
R16767 VSS.n17923 VSS.n1321 1.2805
R16768 VSS.n1412 VSS.n1376 1.2805
R16769 VSS.n1243 VSS.n1242 1.18907
R16770 VSS.n1273 VSS.n1206 1.18907
R16771 VSS.n1108 VSS.n1107 1.18907
R16772 VSS.n1139 VSS.n1072 1.18907
R16773 VSS.n17032 VSS.n16987 1.18907
R16774 VSS.n17084 VSS.n16951 1.18907
R16775 VSS.n17522 VSS.n17521 1.18907
R16776 VSS.n17456 VSS.n17428 1.18907
R16777 VSS.n17624 VSS.n17401 1.18907
R16778 VSS.n17676 VSS.n17365 1.18907
R16779 VSS.n18260 VSS.n18259 1.18907
R16780 VSS.n18290 VSS.n18223 1.18907
R16781 VSS.n18099 VSS.n18098 1.18907
R16782 VSS.n248 VSS.n220 1.18907
R16783 VSS.n9674 VSS.n9451 1.18907
R16784 VSS.n9726 VSS.n9415 1.18907
R16785 VSS.n9572 VSS.n9571 1.18907
R16786 VSS.n9506 VSS.n9478 1.18907
R16787 VSS.n16617 VSS.n16393 1.18907
R16788 VSS.n16669 VSS.n16357 1.18907
R16789 VSS.n16512 VSS.n16468 1.18907
R16790 VSS.n16565 VSS.n16432 1.18907
R16791 VSS.n16024 VSS.n1565 1.18907
R16792 VSS.n16076 VSS.n1529 1.18907
R16793 VSS.n1677 VSS.n1633 1.18907
R16794 VSS.n1730 VSS.n1597 1.18907
R16795 VSS.n2025 VSS.n2024 1.18907
R16796 VSS.n2055 VSS.n1988 1.18907
R16797 VSS.n1864 VSS.n1863 1.18907
R16798 VSS.n1798 VSS.n1770 1.18907
R16799 VSS.n3165 VSS.n2942 1.18907
R16800 VSS.n3217 VSS.n2906 1.18907
R16801 VSS.n3063 VSS.n3062 1.18907
R16802 VSS.n2997 VSS.n2969 1.18907
R16803 VSS.n3757 VSS.n3534 1.18907
R16804 VSS.n3809 VSS.n3498 1.18907
R16805 VSS.n3655 VSS.n3654 1.18907
R16806 VSS.n3589 VSS.n3561 1.18907
R16807 VSS.n4349 VSS.n4126 1.18907
R16808 VSS.n4401 VSS.n4090 1.18907
R16809 VSS.n4247 VSS.n4246 1.18907
R16810 VSS.n4181 VSS.n4153 1.18907
R16811 VSS.n4941 VSS.n4718 1.18907
R16812 VSS.n4993 VSS.n4682 1.18907
R16813 VSS.n4839 VSS.n4838 1.18907
R16814 VSS.n4773 VSS.n4745 1.18907
R16815 VSS.n2621 VSS.n2620 1.18907
R16816 VSS.n2651 VSS.n2584 1.18907
R16817 VSS.n2460 VSS.n2459 1.18907
R16818 VSS.n2394 VSS.n2366 1.18907
R16819 VSS.n5582 VSS.n5581 1.18907
R16820 VSS.n5612 VSS.n5545 1.18907
R16821 VSS.n5421 VSS.n5420 1.18907
R16822 VSS.n5355 VSS.n5327 1.18907
R16823 VSS.n6155 VSS.n6154 1.18907
R16824 VSS.n6185 VSS.n6118 1.18907
R16825 VSS.n5994 VSS.n5993 1.18907
R16826 VSS.n5928 VSS.n5900 1.18907
R16827 VSS.n7898 VSS.n7675 1.18907
R16828 VSS.n7950 VSS.n7639 1.18907
R16829 VSS.n7796 VSS.n7795 1.18907
R16830 VSS.n7730 VSS.n7702 1.18907
R16831 VSS.n8490 VSS.n8267 1.18907
R16832 VSS.n8542 VSS.n8231 1.18907
R16833 VSS.n8388 VSS.n8387 1.18907
R16834 VSS.n8322 VSS.n8294 1.18907
R16835 VSS.n9082 VSS.n8859 1.18907
R16836 VSS.n9134 VSS.n8823 1.18907
R16837 VSS.n8980 VSS.n8979 1.18907
R16838 VSS.n8914 VSS.n8886 1.18907
R16839 VSS.n10266 VSS.n10043 1.18907
R16840 VSS.n10318 VSS.n10007 1.18907
R16841 VSS.n10164 VSS.n10163 1.18907
R16842 VSS.n10098 VSS.n10070 1.18907
R16843 VSS.n10858 VSS.n10635 1.18907
R16844 VSS.n10910 VSS.n10599 1.18907
R16845 VSS.n10756 VSS.n10755 1.18907
R16846 VSS.n10690 VSS.n10662 1.18907
R16847 VSS.n11450 VSS.n11227 1.18907
R16848 VSS.n11502 VSS.n11191 1.18907
R16849 VSS.n11348 VSS.n11347 1.18907
R16850 VSS.n11282 VSS.n11254 1.18907
R16851 VSS.n12042 VSS.n11819 1.18907
R16852 VSS.n12094 VSS.n11783 1.18907
R16853 VSS.n11940 VSS.n11939 1.18907
R16854 VSS.n11874 VSS.n11846 1.18907
R16855 VSS.n12634 VSS.n12411 1.18907
R16856 VSS.n12686 VSS.n12375 1.18907
R16857 VSS.n12532 VSS.n12531 1.18907
R16858 VSS.n12466 VSS.n12438 1.18907
R16859 VSS.n13226 VSS.n13003 1.18907
R16860 VSS.n13278 VSS.n12967 1.18907
R16861 VSS.n13124 VSS.n13123 1.18907
R16862 VSS.n13058 VSS.n13030 1.18907
R16863 VSS.n13818 VSS.n13595 1.18907
R16864 VSS.n13870 VSS.n13559 1.18907
R16865 VSS.n13716 VSS.n13715 1.18907
R16866 VSS.n13650 VSS.n13622 1.18907
R16867 VSS.n14410 VSS.n14187 1.18907
R16868 VSS.n14462 VSS.n14151 1.18907
R16869 VSS.n14308 VSS.n14307 1.18907
R16870 VSS.n14242 VSS.n14214 1.18907
R16871 VSS.n15002 VSS.n14779 1.18907
R16872 VSS.n15054 VSS.n14743 1.18907
R16873 VSS.n14900 VSS.n14899 1.18907
R16874 VSS.n14834 VSS.n14806 1.18907
R16875 VSS.n15594 VSS.n15371 1.18907
R16876 VSS.n15646 VSS.n15335 1.18907
R16877 VSS.n15492 VSS.n15491 1.18907
R16878 VSS.n15426 VSS.n15398 1.18907
R16879 VSS.n6761 VSS.n6760 1.18907
R16880 VSS.n6791 VSS.n6724 1.18907
R16881 VSS.n6600 VSS.n6599 1.18907
R16882 VSS.n6534 VSS.n6506 1.18907
R16883 VSS.n7306 VSS.n7082 1.18907
R16884 VSS.n7358 VSS.n7046 1.18907
R16885 VSS.n7201 VSS.n7157 1.18907
R16886 VSS.n7254 VSS.n7121 1.18907
R16887 VSS.n18618 VSS.n180 1.18907
R16888 VSS.n18670 VSS.n144 1.18907
R16889 VSS.n364 VSS.n363 1.18907
R16890 VSS.n397 VSS.n394 1.18907
R16891 VSS.n584 VSS.n583 1.18907
R16892 VSS.n614 VSS.n544 1.18907
R16893 VSS.n927 VSS.n926 1.18907
R16894 VSS.n958 VSS.n891 1.18907
R16895 VSS.n18039 VSS.n18038 1.13717
R16896 VSS.n1029 VSS.n1027 1.13717
R16897 VSS.n1038 VSS.n1033 1.13717
R16898 VSS.n1050 VSS.n1048 1.13717
R16899 VSS.n1053 VSS.n1051 1.13717
R16900 VSS.n1059 VSS.n1057 1.13717
R16901 VSS.n17136 VSS.n17135 1.13717
R16902 VSS.n17177 VSS.n17176 1.13717
R16903 VSS.n17194 VSS.n17192 1.13717
R16904 VSS.n16861 VSS.n16860 1.13717
R16905 VSS.n16997 VSS.n16996 1.13717
R16906 VSS.n16995 VSS.n16982 1.13717
R16907 VSS.n17041 VSS.n17040 1.13717
R16908 VSS.n16965 VSS.n16961 1.13717
R16909 VSS.n16945 VSS.n16944 1.13717
R16910 VSS.n16933 VSS.n16932 1.13717
R16911 VSS.n17491 VSS.n17490 1.13717
R16912 VSS.n17489 VSS.n17470 1.13717
R16913 VSS.n17540 VSS.n17539 1.13717
R16914 VSS.n17547 VSS.n17443 1.13717
R16915 VSS.n17440 VSS.n17439 1.13717
R16916 VSS.n17422 VSS.n17421 1.13717
R16917 VSS.n17728 VSS.n17727 1.13717
R16918 VSS.n17769 VSS.n17768 1.13717
R16919 VSS.n17786 VSS.n17784 1.13717
R16920 VSS.n17275 VSS.n17274 1.13717
R16921 VSS.n17411 VSS.n17410 1.13717
R16922 VSS.n17409 VSS.n17396 1.13717
R16923 VSS.n17633 VSS.n17632 1.13717
R16924 VSS.n17379 VSS.n17375 1.13717
R16925 VSS.n17359 VSS.n17358 1.13717
R16926 VSS.n17347 VSS.n17346 1.13717
R16927 VSS.n18579 VSS.n18578 1.13717
R16928 VSS.n18181 VSS.n18179 1.13717
R16929 VSS.n18190 VSS.n18185 1.13717
R16930 VSS.n18201 VSS.n18199 1.13717
R16931 VSS.n18204 VSS.n18202 1.13717
R16932 VSS.n18210 VSS.n18208 1.13717
R16933 VSS.n18330 VSS.n18329 1.13717
R16934 VSS.n18351 VSS.n18346 1.13717
R16935 VSS.n18413 VSS.n18412 1.13717
R16936 VSS.n18468 VSS.n18467 1.13717
R16937 VSS.n283 VSS.n282 1.13717
R16938 VSS.n281 VSS.n262 1.13717
R16939 VSS.n18117 VSS.n18116 1.13717
R16940 VSS.n18124 VSS.n235 1.13717
R16941 VSS.n232 VSS.n231 1.13717
R16942 VSS.n214 VSS.n213 1.13717
R16943 VSS.n9461 VSS.n9460 1.13717
R16944 VSS.n9459 VSS.n9446 1.13717
R16945 VSS.n9683 VSS.n9682 1.13717
R16946 VSS.n9429 VSS.n9425 1.13717
R16947 VSS.n9409 VSS.n9408 1.13717
R16948 VSS.n9397 VSS.n9396 1.13717
R16949 VSS.n9778 VSS.n9777 1.13717
R16950 VSS.n9819 VSS.n9818 1.13717
R16951 VSS.n9836 VSS.n9834 1.13717
R16952 VSS.n9326 VSS.n9325 1.13717
R16953 VSS.n9541 VSS.n9540 1.13717
R16954 VSS.n9539 VSS.n9520 1.13717
R16955 VSS.n9590 VSS.n9589 1.13717
R16956 VSS.n9597 VSS.n9493 1.13717
R16957 VSS.n9490 VSS.n9489 1.13717
R16958 VSS.n9472 VSS.n9471 1.13717
R16959 VSS.n16403 VSS.n16402 1.13717
R16960 VSS.n16401 VSS.n16388 1.13717
R16961 VSS.n16626 VSS.n16625 1.13717
R16962 VSS.n16371 VSS.n16367 1.13717
R16963 VSS.n16351 VSS.n16350 1.13717
R16964 VSS.n16339 VSS.n16338 1.13717
R16965 VSS.n16721 VSS.n16720 1.13717
R16966 VSS.n16762 VSS.n16761 1.13717
R16967 VSS.n16779 VSS.n16777 1.13717
R16968 VSS.n16268 VSS.n16267 1.13717
R16969 VSS.n16478 VSS.n16477 1.13717
R16970 VSS.n16476 VSS.n16465 1.13717
R16971 VSS.n16521 VSS.n16520 1.13717
R16972 VSS.n16446 VSS.n16442 1.13717
R16973 VSS.n16426 VSS.n16425 1.13717
R16974 VSS.n16414 VSS.n16413 1.13717
R16975 VSS.n1575 VSS.n1574 1.13717
R16976 VSS.n1573 VSS.n1560 1.13717
R16977 VSS.n16033 VSS.n16032 1.13717
R16978 VSS.n1543 VSS.n1539 1.13717
R16979 VSS.n1523 VSS.n1522 1.13717
R16980 VSS.n1511 VSS.n1510 1.13717
R16981 VSS.n16128 VSS.n16127 1.13717
R16982 VSS.n16169 VSS.n16168 1.13717
R16983 VSS.n16186 VSS.n16184 1.13717
R16984 VSS.n1440 VSS.n1439 1.13717
R16985 VSS.n1643 VSS.n1642 1.13717
R16986 VSS.n1641 VSS.n1630 1.13717
R16987 VSS.n1686 VSS.n1685 1.13717
R16988 VSS.n1611 VSS.n1607 1.13717
R16989 VSS.n1591 VSS.n1590 1.13717
R16990 VSS.n1579 VSS.n1578 1.13717
R16991 VSS.n2344 VSS.n2343 1.13717
R16992 VSS.n1946 VSS.n1944 1.13717
R16993 VSS.n1955 VSS.n1950 1.13717
R16994 VSS.n1966 VSS.n1964 1.13717
R16995 VSS.n1969 VSS.n1967 1.13717
R16996 VSS.n1975 VSS.n1973 1.13717
R16997 VSS.n2094 VSS.n2093 1.13717
R16998 VSS.n2137 VSS.n2136 1.13717
R16999 VSS.n2165 VSS.n2152 1.13717
R17000 VSS.n2219 VSS.n2202 1.13717
R17001 VSS.n1833 VSS.n1832 1.13717
R17002 VSS.n1831 VSS.n1812 1.13717
R17003 VSS.n1882 VSS.n1881 1.13717
R17004 VSS.n1889 VSS.n1785 1.13717
R17005 VSS.n1782 VSS.n1781 1.13717
R17006 VSS.n1764 VSS.n1763 1.13717
R17007 VSS.n2952 VSS.n2951 1.13717
R17008 VSS.n2950 VSS.n2937 1.13717
R17009 VSS.n3174 VSS.n3173 1.13717
R17010 VSS.n2920 VSS.n2916 1.13717
R17011 VSS.n2900 VSS.n2899 1.13717
R17012 VSS.n2888 VSS.n2887 1.13717
R17013 VSS.n3269 VSS.n3268 1.13717
R17014 VSS.n3310 VSS.n3309 1.13717
R17015 VSS.n3327 VSS.n3325 1.13717
R17016 VSS.n2817 VSS.n2816 1.13717
R17017 VSS.n3032 VSS.n3031 1.13717
R17018 VSS.n3030 VSS.n3011 1.13717
R17019 VSS.n3081 VSS.n3080 1.13717
R17020 VSS.n3088 VSS.n2984 1.13717
R17021 VSS.n2981 VSS.n2980 1.13717
R17022 VSS.n2963 VSS.n2962 1.13717
R17023 VSS.n3544 VSS.n3543 1.13717
R17024 VSS.n3542 VSS.n3529 1.13717
R17025 VSS.n3766 VSS.n3765 1.13717
R17026 VSS.n3512 VSS.n3508 1.13717
R17027 VSS.n3492 VSS.n3491 1.13717
R17028 VSS.n3480 VSS.n3479 1.13717
R17029 VSS.n3861 VSS.n3860 1.13717
R17030 VSS.n3902 VSS.n3901 1.13717
R17031 VSS.n3919 VSS.n3917 1.13717
R17032 VSS.n3409 VSS.n3408 1.13717
R17033 VSS.n3624 VSS.n3623 1.13717
R17034 VSS.n3622 VSS.n3603 1.13717
R17035 VSS.n3673 VSS.n3672 1.13717
R17036 VSS.n3680 VSS.n3576 1.13717
R17037 VSS.n3573 VSS.n3572 1.13717
R17038 VSS.n3555 VSS.n3554 1.13717
R17039 VSS.n4136 VSS.n4135 1.13717
R17040 VSS.n4134 VSS.n4121 1.13717
R17041 VSS.n4358 VSS.n4357 1.13717
R17042 VSS.n4104 VSS.n4100 1.13717
R17043 VSS.n4084 VSS.n4083 1.13717
R17044 VSS.n4072 VSS.n4071 1.13717
R17045 VSS.n4453 VSS.n4452 1.13717
R17046 VSS.n4494 VSS.n4493 1.13717
R17047 VSS.n4511 VSS.n4509 1.13717
R17048 VSS.n4001 VSS.n4000 1.13717
R17049 VSS.n4216 VSS.n4215 1.13717
R17050 VSS.n4214 VSS.n4195 1.13717
R17051 VSS.n4265 VSS.n4264 1.13717
R17052 VSS.n4272 VSS.n4168 1.13717
R17053 VSS.n4165 VSS.n4164 1.13717
R17054 VSS.n4147 VSS.n4146 1.13717
R17055 VSS.n4728 VSS.n4727 1.13717
R17056 VSS.n4726 VSS.n4713 1.13717
R17057 VSS.n4950 VSS.n4949 1.13717
R17058 VSS.n4696 VSS.n4692 1.13717
R17059 VSS.n4676 VSS.n4675 1.13717
R17060 VSS.n4664 VSS.n4663 1.13717
R17061 VSS.n5045 VSS.n5044 1.13717
R17062 VSS.n5086 VSS.n5085 1.13717
R17063 VSS.n5103 VSS.n5101 1.13717
R17064 VSS.n4593 VSS.n4592 1.13717
R17065 VSS.n4808 VSS.n4807 1.13717
R17066 VSS.n4806 VSS.n4787 1.13717
R17067 VSS.n4857 VSS.n4856 1.13717
R17068 VSS.n4864 VSS.n4760 1.13717
R17069 VSS.n4757 VSS.n4756 1.13717
R17070 VSS.n4739 VSS.n4738 1.13717
R17071 VSS.n5309 VSS.n5308 1.13717
R17072 VSS.n2542 VSS.n2540 1.13717
R17073 VSS.n2551 VSS.n2546 1.13717
R17074 VSS.n2562 VSS.n2560 1.13717
R17075 VSS.n2565 VSS.n2563 1.13717
R17076 VSS.n2571 VSS.n2569 1.13717
R17077 VSS.n2690 VSS.n2689 1.13717
R17078 VSS.n2733 VSS.n2732 1.13717
R17079 VSS.n2761 VSS.n2748 1.13717
R17080 VSS.n2815 VSS.n2798 1.13717
R17081 VSS.n2429 VSS.n2428 1.13717
R17082 VSS.n2427 VSS.n2408 1.13717
R17083 VSS.n2478 VSS.n2477 1.13717
R17084 VSS.n2485 VSS.n2381 1.13717
R17085 VSS.n2378 VSS.n2377 1.13717
R17086 VSS.n2360 VSS.n2359 1.13717
R17087 VSS.n5882 VSS.n5881 1.13717
R17088 VSS.n5503 VSS.n5501 1.13717
R17089 VSS.n5512 VSS.n5507 1.13717
R17090 VSS.n5523 VSS.n5521 1.13717
R17091 VSS.n5526 VSS.n5524 1.13717
R17092 VSS.n5532 VSS.n5530 1.13717
R17093 VSS.n5651 VSS.n5650 1.13717
R17094 VSS.n5694 VSS.n5693 1.13717
R17095 VSS.n5722 VSS.n5709 1.13717
R17096 VSS.n2 VSS.n1 1.13717
R17097 VSS.n5390 VSS.n5389 1.13717
R17098 VSS.n5388 VSS.n5369 1.13717
R17099 VSS.n5439 VSS.n5438 1.13717
R17100 VSS.n5446 VSS.n5342 1.13717
R17101 VSS.n5339 VSS.n5338 1.13717
R17102 VSS.n5321 VSS.n5320 1.13717
R17103 VSS.n6474 VSS.n6473 1.13717
R17104 VSS.n6076 VSS.n6074 1.13717
R17105 VSS.n6085 VSS.n6080 1.13717
R17106 VSS.n6096 VSS.n6094 1.13717
R17107 VSS.n6099 VSS.n6097 1.13717
R17108 VSS.n6105 VSS.n6103 1.13717
R17109 VSS.n6224 VSS.n6223 1.13717
R17110 VSS.n6267 VSS.n6266 1.13717
R17111 VSS.n6295 VSS.n6282 1.13717
R17112 VSS.n6349 VSS.n6332 1.13717
R17113 VSS.n5963 VSS.n5962 1.13717
R17114 VSS.n5961 VSS.n5942 1.13717
R17115 VSS.n6012 VSS.n6011 1.13717
R17116 VSS.n6019 VSS.n5915 1.13717
R17117 VSS.n5912 VSS.n5911 1.13717
R17118 VSS.n5894 VSS.n5893 1.13717
R17119 VSS.n7685 VSS.n7684 1.13717
R17120 VSS.n7683 VSS.n7670 1.13717
R17121 VSS.n7907 VSS.n7906 1.13717
R17122 VSS.n7653 VSS.n7649 1.13717
R17123 VSS.n7633 VSS.n7632 1.13717
R17124 VSS.n7621 VSS.n7620 1.13717
R17125 VSS.n8002 VSS.n8001 1.13717
R17126 VSS.n8043 VSS.n8042 1.13717
R17127 VSS.n8060 VSS.n8058 1.13717
R17128 VSS.n7550 VSS.n7549 1.13717
R17129 VSS.n7765 VSS.n7764 1.13717
R17130 VSS.n7763 VSS.n7744 1.13717
R17131 VSS.n7814 VSS.n7813 1.13717
R17132 VSS.n7821 VSS.n7717 1.13717
R17133 VSS.n7714 VSS.n7713 1.13717
R17134 VSS.n7696 VSS.n7695 1.13717
R17135 VSS.n8277 VSS.n8276 1.13717
R17136 VSS.n8275 VSS.n8262 1.13717
R17137 VSS.n8499 VSS.n8498 1.13717
R17138 VSS.n8245 VSS.n8241 1.13717
R17139 VSS.n8225 VSS.n8224 1.13717
R17140 VSS.n8213 VSS.n8212 1.13717
R17141 VSS.n8594 VSS.n8593 1.13717
R17142 VSS.n8635 VSS.n8634 1.13717
R17143 VSS.n8652 VSS.n8650 1.13717
R17144 VSS.n8142 VSS.n8141 1.13717
R17145 VSS.n8357 VSS.n8356 1.13717
R17146 VSS.n8355 VSS.n8336 1.13717
R17147 VSS.n8406 VSS.n8405 1.13717
R17148 VSS.n8413 VSS.n8309 1.13717
R17149 VSS.n8306 VSS.n8305 1.13717
R17150 VSS.n8288 VSS.n8287 1.13717
R17151 VSS.n8869 VSS.n8868 1.13717
R17152 VSS.n8867 VSS.n8854 1.13717
R17153 VSS.n9091 VSS.n9090 1.13717
R17154 VSS.n8837 VSS.n8833 1.13717
R17155 VSS.n8817 VSS.n8816 1.13717
R17156 VSS.n8805 VSS.n8804 1.13717
R17157 VSS.n9186 VSS.n9185 1.13717
R17158 VSS.n9227 VSS.n9226 1.13717
R17159 VSS.n9244 VSS.n9242 1.13717
R17160 VSS.n8734 VSS.n8733 1.13717
R17161 VSS.n8949 VSS.n8948 1.13717
R17162 VSS.n8947 VSS.n8928 1.13717
R17163 VSS.n8998 VSS.n8997 1.13717
R17164 VSS.n9005 VSS.n8901 1.13717
R17165 VSS.n8898 VSS.n8897 1.13717
R17166 VSS.n8880 VSS.n8879 1.13717
R17167 VSS.n10053 VSS.n10052 1.13717
R17168 VSS.n10051 VSS.n10038 1.13717
R17169 VSS.n10275 VSS.n10274 1.13717
R17170 VSS.n10021 VSS.n10017 1.13717
R17171 VSS.n10001 VSS.n10000 1.13717
R17172 VSS.n9989 VSS.n9988 1.13717
R17173 VSS.n10370 VSS.n10369 1.13717
R17174 VSS.n10411 VSS.n10410 1.13717
R17175 VSS.n10428 VSS.n10426 1.13717
R17176 VSS.n9918 VSS.n9917 1.13717
R17177 VSS.n10133 VSS.n10132 1.13717
R17178 VSS.n10131 VSS.n10112 1.13717
R17179 VSS.n10182 VSS.n10181 1.13717
R17180 VSS.n10189 VSS.n10085 1.13717
R17181 VSS.n10082 VSS.n10081 1.13717
R17182 VSS.n10064 VSS.n10063 1.13717
R17183 VSS.n10645 VSS.n10644 1.13717
R17184 VSS.n10643 VSS.n10630 1.13717
R17185 VSS.n10867 VSS.n10866 1.13717
R17186 VSS.n10613 VSS.n10609 1.13717
R17187 VSS.n10593 VSS.n10592 1.13717
R17188 VSS.n10581 VSS.n10580 1.13717
R17189 VSS.n10962 VSS.n10961 1.13717
R17190 VSS.n11003 VSS.n11002 1.13717
R17191 VSS.n11020 VSS.n11018 1.13717
R17192 VSS.n10510 VSS.n10509 1.13717
R17193 VSS.n10725 VSS.n10724 1.13717
R17194 VSS.n10723 VSS.n10704 1.13717
R17195 VSS.n10774 VSS.n10773 1.13717
R17196 VSS.n10781 VSS.n10677 1.13717
R17197 VSS.n10674 VSS.n10673 1.13717
R17198 VSS.n10656 VSS.n10655 1.13717
R17199 VSS.n11237 VSS.n11236 1.13717
R17200 VSS.n11235 VSS.n11222 1.13717
R17201 VSS.n11459 VSS.n11458 1.13717
R17202 VSS.n11205 VSS.n11201 1.13717
R17203 VSS.n11185 VSS.n11184 1.13717
R17204 VSS.n11173 VSS.n11172 1.13717
R17205 VSS.n11554 VSS.n11553 1.13717
R17206 VSS.n11595 VSS.n11594 1.13717
R17207 VSS.n11612 VSS.n11610 1.13717
R17208 VSS.n11102 VSS.n11101 1.13717
R17209 VSS.n11317 VSS.n11316 1.13717
R17210 VSS.n11315 VSS.n11296 1.13717
R17211 VSS.n11366 VSS.n11365 1.13717
R17212 VSS.n11373 VSS.n11269 1.13717
R17213 VSS.n11266 VSS.n11265 1.13717
R17214 VSS.n11248 VSS.n11247 1.13717
R17215 VSS.n11829 VSS.n11828 1.13717
R17216 VSS.n11827 VSS.n11814 1.13717
R17217 VSS.n12051 VSS.n12050 1.13717
R17218 VSS.n11797 VSS.n11793 1.13717
R17219 VSS.n11777 VSS.n11776 1.13717
R17220 VSS.n11765 VSS.n11764 1.13717
R17221 VSS.n12146 VSS.n12145 1.13717
R17222 VSS.n12187 VSS.n12186 1.13717
R17223 VSS.n12204 VSS.n12202 1.13717
R17224 VSS.n11694 VSS.n11693 1.13717
R17225 VSS.n11909 VSS.n11908 1.13717
R17226 VSS.n11907 VSS.n11888 1.13717
R17227 VSS.n11958 VSS.n11957 1.13717
R17228 VSS.n11965 VSS.n11861 1.13717
R17229 VSS.n11858 VSS.n11857 1.13717
R17230 VSS.n11840 VSS.n11839 1.13717
R17231 VSS.n12421 VSS.n12420 1.13717
R17232 VSS.n12419 VSS.n12406 1.13717
R17233 VSS.n12643 VSS.n12642 1.13717
R17234 VSS.n12389 VSS.n12385 1.13717
R17235 VSS.n12369 VSS.n12368 1.13717
R17236 VSS.n12357 VSS.n12356 1.13717
R17237 VSS.n12738 VSS.n12737 1.13717
R17238 VSS.n12779 VSS.n12778 1.13717
R17239 VSS.n12796 VSS.n12794 1.13717
R17240 VSS.n12286 VSS.n12285 1.13717
R17241 VSS.n12501 VSS.n12500 1.13717
R17242 VSS.n12499 VSS.n12480 1.13717
R17243 VSS.n12550 VSS.n12549 1.13717
R17244 VSS.n12557 VSS.n12453 1.13717
R17245 VSS.n12450 VSS.n12449 1.13717
R17246 VSS.n12432 VSS.n12431 1.13717
R17247 VSS.n13013 VSS.n13012 1.13717
R17248 VSS.n13011 VSS.n12998 1.13717
R17249 VSS.n13235 VSS.n13234 1.13717
R17250 VSS.n12981 VSS.n12977 1.13717
R17251 VSS.n12961 VSS.n12960 1.13717
R17252 VSS.n12949 VSS.n12948 1.13717
R17253 VSS.n13330 VSS.n13329 1.13717
R17254 VSS.n13371 VSS.n13370 1.13717
R17255 VSS.n13388 VSS.n13386 1.13717
R17256 VSS.n12878 VSS.n12877 1.13717
R17257 VSS.n13093 VSS.n13092 1.13717
R17258 VSS.n13091 VSS.n13072 1.13717
R17259 VSS.n13142 VSS.n13141 1.13717
R17260 VSS.n13149 VSS.n13045 1.13717
R17261 VSS.n13042 VSS.n13041 1.13717
R17262 VSS.n13024 VSS.n13023 1.13717
R17263 VSS.n13605 VSS.n13604 1.13717
R17264 VSS.n13603 VSS.n13590 1.13717
R17265 VSS.n13827 VSS.n13826 1.13717
R17266 VSS.n13573 VSS.n13569 1.13717
R17267 VSS.n13553 VSS.n13552 1.13717
R17268 VSS.n13541 VSS.n13540 1.13717
R17269 VSS.n13922 VSS.n13921 1.13717
R17270 VSS.n13963 VSS.n13962 1.13717
R17271 VSS.n13980 VSS.n13978 1.13717
R17272 VSS.n13470 VSS.n13469 1.13717
R17273 VSS.n13685 VSS.n13684 1.13717
R17274 VSS.n13683 VSS.n13664 1.13717
R17275 VSS.n13734 VSS.n13733 1.13717
R17276 VSS.n13741 VSS.n13637 1.13717
R17277 VSS.n13634 VSS.n13633 1.13717
R17278 VSS.n13616 VSS.n13615 1.13717
R17279 VSS.n14197 VSS.n14196 1.13717
R17280 VSS.n14195 VSS.n14182 1.13717
R17281 VSS.n14419 VSS.n14418 1.13717
R17282 VSS.n14165 VSS.n14161 1.13717
R17283 VSS.n14145 VSS.n14144 1.13717
R17284 VSS.n14133 VSS.n14132 1.13717
R17285 VSS.n14514 VSS.n14513 1.13717
R17286 VSS.n14555 VSS.n14554 1.13717
R17287 VSS.n14572 VSS.n14570 1.13717
R17288 VSS.n14062 VSS.n14061 1.13717
R17289 VSS.n14277 VSS.n14276 1.13717
R17290 VSS.n14275 VSS.n14256 1.13717
R17291 VSS.n14326 VSS.n14325 1.13717
R17292 VSS.n14333 VSS.n14229 1.13717
R17293 VSS.n14226 VSS.n14225 1.13717
R17294 VSS.n14208 VSS.n14207 1.13717
R17295 VSS.n14789 VSS.n14788 1.13717
R17296 VSS.n14787 VSS.n14774 1.13717
R17297 VSS.n15011 VSS.n15010 1.13717
R17298 VSS.n14757 VSS.n14753 1.13717
R17299 VSS.n14737 VSS.n14736 1.13717
R17300 VSS.n14725 VSS.n14724 1.13717
R17301 VSS.n15106 VSS.n15105 1.13717
R17302 VSS.n15147 VSS.n15146 1.13717
R17303 VSS.n15164 VSS.n15162 1.13717
R17304 VSS.n14654 VSS.n14653 1.13717
R17305 VSS.n14869 VSS.n14868 1.13717
R17306 VSS.n14867 VSS.n14848 1.13717
R17307 VSS.n14918 VSS.n14917 1.13717
R17308 VSS.n14925 VSS.n14821 1.13717
R17309 VSS.n14818 VSS.n14817 1.13717
R17310 VSS.n14800 VSS.n14799 1.13717
R17311 VSS.n15381 VSS.n15380 1.13717
R17312 VSS.n15379 VSS.n15366 1.13717
R17313 VSS.n15603 VSS.n15602 1.13717
R17314 VSS.n15349 VSS.n15345 1.13717
R17315 VSS.n15329 VSS.n15328 1.13717
R17316 VSS.n15317 VSS.n15316 1.13717
R17317 VSS.n15698 VSS.n15697 1.13717
R17318 VSS.n15739 VSS.n15738 1.13717
R17319 VSS.n15756 VSS.n15754 1.13717
R17320 VSS.n15246 VSS.n15245 1.13717
R17321 VSS.n15461 VSS.n15460 1.13717
R17322 VSS.n15459 VSS.n15440 1.13717
R17323 VSS.n15510 VSS.n15509 1.13717
R17324 VSS.n15517 VSS.n15413 1.13717
R17325 VSS.n15410 VSS.n15409 1.13717
R17326 VSS.n15392 VSS.n15391 1.13717
R17327 VSS.n15962 VSS.n15961 1.13717
R17328 VSS.n6682 VSS.n6680 1.13717
R17329 VSS.n6691 VSS.n6686 1.13717
R17330 VSS.n6702 VSS.n6700 1.13717
R17331 VSS.n6705 VSS.n6703 1.13717
R17332 VSS.n6711 VSS.n6709 1.13717
R17333 VSS.n6830 VSS.n6829 1.13717
R17334 VSS.n6873 VSS.n6872 1.13717
R17335 VSS.n6901 VSS.n6888 1.13717
R17336 VSS.n6955 VSS.n6938 1.13717
R17337 VSS.n6569 VSS.n6568 1.13717
R17338 VSS.n6567 VSS.n6548 1.13717
R17339 VSS.n6618 VSS.n6617 1.13717
R17340 VSS.n6625 VSS.n6521 1.13717
R17341 VSS.n6518 VSS.n6517 1.13717
R17342 VSS.n6500 VSS.n6499 1.13717
R17343 VSS.n7092 VSS.n7091 1.13717
R17344 VSS.n7090 VSS.n7077 1.13717
R17345 VSS.n7315 VSS.n7314 1.13717
R17346 VSS.n7060 VSS.n7056 1.13717
R17347 VSS.n7040 VSS.n7039 1.13717
R17348 VSS.n7028 VSS.n7027 1.13717
R17349 VSS.n7410 VSS.n7409 1.13717
R17350 VSS.n7451 VSS.n7450 1.13717
R17351 VSS.n7468 VSS.n7466 1.13717
R17352 VSS.n6957 VSS.n6956 1.13717
R17353 VSS.n7167 VSS.n7166 1.13717
R17354 VSS.n7165 VSS.n7154 1.13717
R17355 VSS.n7210 VSS.n7209 1.13717
R17356 VSS.n7135 VSS.n7131 1.13717
R17357 VSS.n7115 VSS.n7114 1.13717
R17358 VSS.n7103 VSS.n7102 1.13717
R17359 VSS.n190 VSS.n189 1.13717
R17360 VSS.n188 VSS.n175 1.13717
R17361 VSS.n18627 VSS.n18626 1.13717
R17362 VSS.n158 VSS.n154 1.13717
R17363 VSS.n138 VSS.n137 1.13717
R17364 VSS.n126 VSS.n125 1.13717
R17365 VSS.n18722 VSS.n18721 1.13717
R17366 VSS.n18763 VSS.n18762 1.13717
R17367 VSS.n18780 VSS.n18778 1.13717
R17368 VSS.n55 VSS.n54 1.13717
R17369 VSS.n448 VSS.n447 1.13717
R17370 VSS.n296 VSS.n294 1.13717
R17371 VSS.n305 VSS.n300 1.13717
R17372 VSS.n317 VSS.n315 1.13717
R17373 VSS.n320 VSS.n318 1.13717
R17374 VSS.n194 VSS.n193 1.13717
R17375 VSS.n52 VSS.n51 1.13717
R17376 VSS.n496 VSS.n495 1.13717
R17377 VSS.n502 VSS.n500 1.13717
R17378 VSS.n511 VSS.n506 1.13717
R17379 VSS.n522 VSS.n520 1.13717
R17380 VSS.n525 VSS.n523 1.13717
R17381 VSS.n531 VSS.n529 1.13717
R17382 VSS.n653 VSS.n652 1.13717
R17383 VSS.n696 VSS.n695 1.13717
R17384 VSS.n724 VSS.n711 1.13717
R17385 VSS.n1013 VSS.n1012 1.13717
R17386 VSS.n462 VSS.n460 1.13717
R17387 VSS.n471 VSS.n466 1.13717
R17388 VSS.n483 VSS.n481 1.13717
R17389 VSS.n486 VSS.n484 1.13717
R17390 VSS.n492 VSS.n490 1.13717
R17391 VSS.n17990 VSS.n17989 1.13717
R17392 VSS.n1164 VSS.n1162 1.13717
R17393 VSS.n1173 VSS.n1168 1.13717
R17394 VSS.n1184 VSS.n1182 1.13717
R17395 VSS.n1187 VSS.n1185 1.13717
R17396 VSS.n1193 VSS.n1191 1.13717
R17397 VSS.n1312 VSS.n1311 1.13717
R17398 VSS.n1355 VSS.n1354 1.13717
R17399 VSS.n1383 VSS.n1370 1.13717
R17400 VSS.n1437 VSS.n1420 1.13717
R17401 VSS.n1179 VSS.n1175 1.1255
R17402 VSS.n17056 VSS.n16968 1.1255
R17403 VSS.n17648 VSS.n17382 1.1255
R17404 VSS.n18196 VSS.n18192 1.1255
R17405 VSS.n9698 VSS.n9432 1.1255
R17406 VSS.n16641 VSS.n16374 1.1255
R17407 VSS.n16048 VSS.n1546 1.1255
R17408 VSS.n1961 VSS.n1957 1.1255
R17409 VSS.n3189 VSS.n2923 1.1255
R17410 VSS.n3781 VSS.n3515 1.1255
R17411 VSS.n4373 VSS.n4107 1.1255
R17412 VSS.n4965 VSS.n4699 1.1255
R17413 VSS.n2557 VSS.n2553 1.1255
R17414 VSS.n5518 VSS.n5514 1.1255
R17415 VSS.n6091 VSS.n6087 1.1255
R17416 VSS.n7922 VSS.n7656 1.1255
R17417 VSS.n8514 VSS.n8248 1.1255
R17418 VSS.n9106 VSS.n8840 1.1255
R17419 VSS.n10290 VSS.n10024 1.1255
R17420 VSS.n10882 VSS.n10616 1.1255
R17421 VSS.n11474 VSS.n11208 1.1255
R17422 VSS.n12066 VSS.n11800 1.1255
R17423 VSS.n12658 VSS.n12392 1.1255
R17424 VSS.n13250 VSS.n12984 1.1255
R17425 VSS.n13842 VSS.n13576 1.1255
R17426 VSS.n14434 VSS.n14168 1.1255
R17427 VSS.n15026 VSS.n14760 1.1255
R17428 VSS.n15618 VSS.n15352 1.1255
R17429 VSS.n6697 VSS.n6693 1.1255
R17430 VSS.n7330 VSS.n7063 1.1255
R17431 VSS.n18642 VSS.n161 1.1255
R17432 VSS.n517 VSS.n513 1.1255
R17433 VSS.n17116 VSS.n16922 1.09764
R17434 VSS.n17259 VSS.n17257 1.09764
R17435 VSS.n17708 VSS.n17336 1.09764
R17436 VSS.n17851 VSS.n17849 1.09764
R17437 VSS.n18528 VSS.n18527 1.09764
R17438 VSS.n18455 VSS.n18421 1.09764
R17439 VSS.n9758 VSS.n9386 1.09764
R17440 VSS.n9902 VSS.n9900 1.09764
R17441 VSS.n16701 VSS.n16328 1.09764
R17442 VSS.n16845 VSS.n16843 1.09764
R17443 VSS.n16108 VSS.n1500 1.09764
R17444 VSS.n16252 VSS.n16250 1.09764
R17445 VSS.n2293 VSS.n2292 1.09764
R17446 VSS.n2232 VSS.n2174 1.09764
R17447 VSS.n3249 VSS.n2877 1.09764
R17448 VSS.n3393 VSS.n3391 1.09764
R17449 VSS.n3841 VSS.n3469 1.09764
R17450 VSS.n3985 VSS.n3983 1.09764
R17451 VSS.n4433 VSS.n4061 1.09764
R17452 VSS.n4577 VSS.n4575 1.09764
R17453 VSS.n5025 VSS.n4653 1.09764
R17454 VSS.n5169 VSS.n5167 1.09764
R17455 VSS.n5258 VSS.n5257 1.09764
R17456 VSS.n5197 VSS.n2770 1.09764
R17457 VSS.n5831 VSS.n5830 1.09764
R17458 VSS.n5770 VSS.n5744 1.09764
R17459 VSS.n6423 VSS.n6422 1.09764
R17460 VSS.n6362 VSS.n6304 1.09764
R17461 VSS.n7982 VSS.n7610 1.09764
R17462 VSS.n8126 VSS.n8124 1.09764
R17463 VSS.n8574 VSS.n8202 1.09764
R17464 VSS.n8718 VSS.n8716 1.09764
R17465 VSS.n9166 VSS.n8794 1.09764
R17466 VSS.n9310 VSS.n9308 1.09764
R17467 VSS.n10350 VSS.n9978 1.09764
R17468 VSS.n10494 VSS.n10492 1.09764
R17469 VSS.n10942 VSS.n10570 1.09764
R17470 VSS.n11086 VSS.n11084 1.09764
R17471 VSS.n11534 VSS.n11162 1.09764
R17472 VSS.n11678 VSS.n11676 1.09764
R17473 VSS.n12126 VSS.n11754 1.09764
R17474 VSS.n12270 VSS.n12268 1.09764
R17475 VSS.n12718 VSS.n12346 1.09764
R17476 VSS.n12862 VSS.n12860 1.09764
R17477 VSS.n13310 VSS.n12938 1.09764
R17478 VSS.n13454 VSS.n13452 1.09764
R17479 VSS.n13902 VSS.n13530 1.09764
R17480 VSS.n14046 VSS.n14044 1.09764
R17481 VSS.n14494 VSS.n14122 1.09764
R17482 VSS.n14638 VSS.n14636 1.09764
R17483 VSS.n15086 VSS.n14714 1.09764
R17484 VSS.n15230 VSS.n15228 1.09764
R17485 VSS.n15678 VSS.n15306 1.09764
R17486 VSS.n15822 VSS.n15820 1.09764
R17487 VSS.n15911 VSS.n15910 1.09764
R17488 VSS.n15850 VSS.n6910 1.09764
R17489 VSS.n7390 VSS.n7017 1.09764
R17490 VSS.n7534 VSS.n7532 1.09764
R17491 VSS.n18702 VSS.n115 1.09764
R17492 VSS.n18846 VSS.n18844 1.09764
R17493 VSS.n825 VSS.n824 1.09764
R17494 VSS.n18868 VSS.n48 1.09764
R17495 VSS.n17939 VSS.n17938 1.09764
R17496 VSS.n17878 VSS.n1392 1.09764
R17497 VSS.n16899 VSS.n16897 1.04225
R17498 VSS.n17313 VSS.n17311 1.04225
R17499 VSS.n18356 VSS.n18354 1.04225
R17500 VSS.n9363 VSS.n9361 1.04225
R17501 VSS.n16305 VSS.n16303 1.04225
R17502 VSS.n1477 VSS.n1475 1.04225
R17503 VSS.n2129 VSS.n2127 1.04225
R17504 VSS.n2854 VSS.n2852 1.04225
R17505 VSS.n3446 VSS.n3444 1.04225
R17506 VSS.n4038 VSS.n4036 1.04225
R17507 VSS.n4630 VSS.n4628 1.04225
R17508 VSS.n2725 VSS.n2723 1.04225
R17509 VSS.n5686 VSS.n5684 1.04225
R17510 VSS.n6259 VSS.n6257 1.04225
R17511 VSS.n7587 VSS.n7585 1.04225
R17512 VSS.n8179 VSS.n8177 1.04225
R17513 VSS.n8771 VSS.n8769 1.04225
R17514 VSS.n9955 VSS.n9953 1.04225
R17515 VSS.n10547 VSS.n10545 1.04225
R17516 VSS.n11139 VSS.n11137 1.04225
R17517 VSS.n11731 VSS.n11729 1.04225
R17518 VSS.n12323 VSS.n12321 1.04225
R17519 VSS.n12915 VSS.n12913 1.04225
R17520 VSS.n13507 VSS.n13505 1.04225
R17521 VSS.n14099 VSS.n14097 1.04225
R17522 VSS.n14691 VSS.n14689 1.04225
R17523 VSS.n15283 VSS.n15281 1.04225
R17524 VSS.n6865 VSS.n6863 1.04225
R17525 VSS.n6994 VSS.n6992 1.04225
R17526 VSS.n92 VSS.n90 1.04225
R17527 VSS.n688 VSS.n686 1.04225
R17528 VSS.n1347 VSS.n1345 1.04225
R17529 VSS.n1221 VSS.n1158 1.00621
R17530 VSS.n1284 VSS.n1197 1.00621
R17531 VSS.n1088 VSS.n1023 1.00621
R17532 VSS.n1150 VSS.n1063 1.00621
R17533 VSS.n17150 VSS.n16922 1.00621
R17534 VSS.n17152 VSS.n17151 1.00621
R17535 VSS.n17200 VSS.n17199 1.00621
R17536 VSS.n17005 VSS.n17000 1.00621
R17537 VSS.n17101 VSS.n16936 1.00621
R17538 VSS.n17500 VSS.n17494 1.00621
R17539 VSS.n17436 VSS.n17425 1.00621
R17540 VSS.n17742 VSS.n17336 1.00621
R17541 VSS.n17744 VSS.n17743 1.00621
R17542 VSS.n17792 VSS.n17791 1.00621
R17543 VSS.n17419 VSS.n17414 1.00621
R17544 VSS.n17693 VSS.n17350 1.00621
R17545 VSS.n18238 VSS.n211 1.00621
R17546 VSS.n18301 VSS.n18214 1.00621
R17547 VSS.n18527 VSS.n18313 1.00621
R17548 VSS.n18365 VSS.n18364 1.00621
R17549 VSS.n18405 VSS.n18404 1.00621
R17550 VSS.n18077 VSS.n286 1.00621
R17551 VSS.n228 VSS.n217 1.00621
R17552 VSS.n9469 VSS.n9464 1.00621
R17553 VSS.n9743 VSS.n9400 1.00621
R17554 VSS.n9792 VSS.n9386 1.00621
R17555 VSS.n9794 VSS.n9793 1.00621
R17556 VSS.n9842 VSS.n9841 1.00621
R17557 VSS.n9550 VSS.n9544 1.00621
R17558 VSS.n9486 VSS.n9475 1.00621
R17559 VSS.n16411 VSS.n16406 1.00621
R17560 VSS.n16686 VSS.n16342 1.00621
R17561 VSS.n16735 VSS.n16328 1.00621
R17562 VSS.n16737 VSS.n16736 1.00621
R17563 VSS.n16785 VSS.n16784 1.00621
R17564 VSS.n16486 VSS.n16481 1.00621
R17565 VSS.n16582 VSS.n16417 1.00621
R17566 VSS.n1754 VSS.n1753 1.00621
R17567 VSS.n16093 VSS.n1514 1.00621
R17568 VSS.n16142 VSS.n1500 1.00621
R17569 VSS.n16144 VSS.n16143 1.00621
R17570 VSS.n16192 VSS.n16191 1.00621
R17571 VSS.n1651 VSS.n1646 1.00621
R17572 VSS.n1747 VSS.n1582 1.00621
R17573 VSS.n2003 VSS.n1761 1.00621
R17574 VSS.n2066 VSS.n1979 1.00621
R17575 VSS.n2292 VSS.n2078 1.00621
R17576 VSS.n2285 VSS.n2284 1.00621
R17577 VSS.n2179 VSS.n2178 1.00621
R17578 VSS.n1842 VSS.n1836 1.00621
R17579 VSS.n1778 VSS.n1767 1.00621
R17580 VSS.n2960 VSS.n2955 1.00621
R17581 VSS.n3234 VSS.n2891 1.00621
R17582 VSS.n3283 VSS.n2877 1.00621
R17583 VSS.n3285 VSS.n3284 1.00621
R17584 VSS.n3333 VSS.n3332 1.00621
R17585 VSS.n3041 VSS.n3035 1.00621
R17586 VSS.n2977 VSS.n2966 1.00621
R17587 VSS.n3552 VSS.n3547 1.00621
R17588 VSS.n3826 VSS.n3483 1.00621
R17589 VSS.n3875 VSS.n3469 1.00621
R17590 VSS.n3877 VSS.n3876 1.00621
R17591 VSS.n3925 VSS.n3924 1.00621
R17592 VSS.n3633 VSS.n3627 1.00621
R17593 VSS.n3569 VSS.n3558 1.00621
R17594 VSS.n4144 VSS.n4139 1.00621
R17595 VSS.n4418 VSS.n4075 1.00621
R17596 VSS.n4467 VSS.n4061 1.00621
R17597 VSS.n4469 VSS.n4468 1.00621
R17598 VSS.n4517 VSS.n4516 1.00621
R17599 VSS.n4225 VSS.n4219 1.00621
R17600 VSS.n4161 VSS.n4150 1.00621
R17601 VSS.n4736 VSS.n4731 1.00621
R17602 VSS.n5010 VSS.n4667 1.00621
R17603 VSS.n5059 VSS.n4653 1.00621
R17604 VSS.n5061 VSS.n5060 1.00621
R17605 VSS.n5109 VSS.n5108 1.00621
R17606 VSS.n4817 VSS.n4811 1.00621
R17607 VSS.n4753 VSS.n4742 1.00621
R17608 VSS.n2599 VSS.n2357 1.00621
R17609 VSS.n2662 VSS.n2575 1.00621
R17610 VSS.n5257 VSS.n2674 1.00621
R17611 VSS.n5250 VSS.n5249 1.00621
R17612 VSS.n2775 VSS.n2774 1.00621
R17613 VSS.n2438 VSS.n2432 1.00621
R17614 VSS.n2374 VSS.n2363 1.00621
R17615 VSS.n5560 VSS.n5318 1.00621
R17616 VSS.n5623 VSS.n5536 1.00621
R17617 VSS.n5830 VSS.n5635 1.00621
R17618 VSS.n5823 VSS.n5822 1.00621
R17619 VSS.n5749 VSS.n5748 1.00621
R17620 VSS.n5399 VSS.n5393 1.00621
R17621 VSS.n5335 VSS.n5324 1.00621
R17622 VSS.n6133 VSS.n5891 1.00621
R17623 VSS.n6196 VSS.n6109 1.00621
R17624 VSS.n6422 VSS.n6208 1.00621
R17625 VSS.n6415 VSS.n6414 1.00621
R17626 VSS.n6309 VSS.n6308 1.00621
R17627 VSS.n5972 VSS.n5966 1.00621
R17628 VSS.n5908 VSS.n5897 1.00621
R17629 VSS.n7693 VSS.n7688 1.00621
R17630 VSS.n7967 VSS.n7624 1.00621
R17631 VSS.n8016 VSS.n7610 1.00621
R17632 VSS.n8018 VSS.n8017 1.00621
R17633 VSS.n8066 VSS.n8065 1.00621
R17634 VSS.n7774 VSS.n7768 1.00621
R17635 VSS.n7710 VSS.n7699 1.00621
R17636 VSS.n8285 VSS.n8280 1.00621
R17637 VSS.n8559 VSS.n8216 1.00621
R17638 VSS.n8608 VSS.n8202 1.00621
R17639 VSS.n8610 VSS.n8609 1.00621
R17640 VSS.n8658 VSS.n8657 1.00621
R17641 VSS.n8366 VSS.n8360 1.00621
R17642 VSS.n8302 VSS.n8291 1.00621
R17643 VSS.n8877 VSS.n8872 1.00621
R17644 VSS.n9151 VSS.n8808 1.00621
R17645 VSS.n9200 VSS.n8794 1.00621
R17646 VSS.n9202 VSS.n9201 1.00621
R17647 VSS.n9250 VSS.n9249 1.00621
R17648 VSS.n8958 VSS.n8952 1.00621
R17649 VSS.n8894 VSS.n8883 1.00621
R17650 VSS.n10061 VSS.n10056 1.00621
R17651 VSS.n10335 VSS.n9992 1.00621
R17652 VSS.n10384 VSS.n9978 1.00621
R17653 VSS.n10386 VSS.n10385 1.00621
R17654 VSS.n10434 VSS.n10433 1.00621
R17655 VSS.n10142 VSS.n10136 1.00621
R17656 VSS.n10078 VSS.n10067 1.00621
R17657 VSS.n10653 VSS.n10648 1.00621
R17658 VSS.n10927 VSS.n10584 1.00621
R17659 VSS.n10976 VSS.n10570 1.00621
R17660 VSS.n10978 VSS.n10977 1.00621
R17661 VSS.n11026 VSS.n11025 1.00621
R17662 VSS.n10734 VSS.n10728 1.00621
R17663 VSS.n10670 VSS.n10659 1.00621
R17664 VSS.n11245 VSS.n11240 1.00621
R17665 VSS.n11519 VSS.n11176 1.00621
R17666 VSS.n11568 VSS.n11162 1.00621
R17667 VSS.n11570 VSS.n11569 1.00621
R17668 VSS.n11618 VSS.n11617 1.00621
R17669 VSS.n11326 VSS.n11320 1.00621
R17670 VSS.n11262 VSS.n11251 1.00621
R17671 VSS.n11837 VSS.n11832 1.00621
R17672 VSS.n12111 VSS.n11768 1.00621
R17673 VSS.n12160 VSS.n11754 1.00621
R17674 VSS.n12162 VSS.n12161 1.00621
R17675 VSS.n12210 VSS.n12209 1.00621
R17676 VSS.n11918 VSS.n11912 1.00621
R17677 VSS.n11854 VSS.n11843 1.00621
R17678 VSS.n12429 VSS.n12424 1.00621
R17679 VSS.n12703 VSS.n12360 1.00621
R17680 VSS.n12752 VSS.n12346 1.00621
R17681 VSS.n12754 VSS.n12753 1.00621
R17682 VSS.n12802 VSS.n12801 1.00621
R17683 VSS.n12510 VSS.n12504 1.00621
R17684 VSS.n12446 VSS.n12435 1.00621
R17685 VSS.n13021 VSS.n13016 1.00621
R17686 VSS.n13295 VSS.n12952 1.00621
R17687 VSS.n13344 VSS.n12938 1.00621
R17688 VSS.n13346 VSS.n13345 1.00621
R17689 VSS.n13394 VSS.n13393 1.00621
R17690 VSS.n13102 VSS.n13096 1.00621
R17691 VSS.n13038 VSS.n13027 1.00621
R17692 VSS.n13613 VSS.n13608 1.00621
R17693 VSS.n13887 VSS.n13544 1.00621
R17694 VSS.n13936 VSS.n13530 1.00621
R17695 VSS.n13938 VSS.n13937 1.00621
R17696 VSS.n13986 VSS.n13985 1.00621
R17697 VSS.n13694 VSS.n13688 1.00621
R17698 VSS.n13630 VSS.n13619 1.00621
R17699 VSS.n14205 VSS.n14200 1.00621
R17700 VSS.n14479 VSS.n14136 1.00621
R17701 VSS.n14528 VSS.n14122 1.00621
R17702 VSS.n14530 VSS.n14529 1.00621
R17703 VSS.n14578 VSS.n14577 1.00621
R17704 VSS.n14286 VSS.n14280 1.00621
R17705 VSS.n14222 VSS.n14211 1.00621
R17706 VSS.n14797 VSS.n14792 1.00621
R17707 VSS.n15071 VSS.n14728 1.00621
R17708 VSS.n15120 VSS.n14714 1.00621
R17709 VSS.n15122 VSS.n15121 1.00621
R17710 VSS.n15170 VSS.n15169 1.00621
R17711 VSS.n14878 VSS.n14872 1.00621
R17712 VSS.n14814 VSS.n14803 1.00621
R17713 VSS.n15389 VSS.n15384 1.00621
R17714 VSS.n15663 VSS.n15320 1.00621
R17715 VSS.n15712 VSS.n15306 1.00621
R17716 VSS.n15714 VSS.n15713 1.00621
R17717 VSS.n15762 VSS.n15761 1.00621
R17718 VSS.n15470 VSS.n15464 1.00621
R17719 VSS.n15406 VSS.n15395 1.00621
R17720 VSS.n6739 VSS.n6497 1.00621
R17721 VSS.n6802 VSS.n6715 1.00621
R17722 VSS.n15910 VSS.n6814 1.00621
R17723 VSS.n15903 VSS.n15902 1.00621
R17724 VSS.n6915 VSS.n6914 1.00621
R17725 VSS.n6578 VSS.n6572 1.00621
R17726 VSS.n6514 VSS.n6503 1.00621
R17727 VSS.n7100 VSS.n7095 1.00621
R17728 VSS.n7375 VSS.n7031 1.00621
R17729 VSS.n7424 VSS.n7017 1.00621
R17730 VSS.n7426 VSS.n7425 1.00621
R17731 VSS.n7474 VSS.n7473 1.00621
R17732 VSS.n7175 VSS.n7170 1.00621
R17733 VSS.n7271 VSS.n7106 1.00621
R17734 VSS.n203 VSS.n202 1.00621
R17735 VSS.n18687 VSS.n129 1.00621
R17736 VSS.n18736 VSS.n115 1.00621
R17737 VSS.n18738 VSS.n18737 1.00621
R17738 VSS.n18786 VSS.n18785 1.00621
R17739 VSS.n357 VSS.n290 1.00621
R17740 VSS.n403 VSS.n197 1.00621
R17741 VSS.n564 VSS.n557 1.00621
R17742 VSS.n625 VSS.n535 1.00621
R17743 VSS.n824 VSS.n637 1.00621
R17744 VSS.n817 VSS.n816 1.00621
R17745 VSS.n747 VSS.n746 1.00621
R17746 VSS.n907 VSS.n456 1.00621
R17747 VSS.n969 VSS.n882 1.00621
R17748 VSS.n17938 VSS.n1296 1.00621
R17749 VSS.n17931 VSS.n17930 1.00621
R17750 VSS.n1397 VSS.n1396 1.00621
R17751 VSS.n17122 VSS.n17107 0.914786
R17752 VSS.n17184 VSS.n17183 0.914786
R17753 VSS.n17185 VSS.n16895 0.914786
R17754 VSS.n17241 VSS.n17240 0.914786
R17755 VSS.n17257 VSS.n16870 0.914786
R17756 VSS.n17267 VSS.n17266 0.914786
R17757 VSS.n17714 VSS.n17699 0.914786
R17758 VSS.n17776 VSS.n17775 0.914786
R17759 VSS.n17777 VSS.n17309 0.914786
R17760 VSS.n17833 VSS.n17832 0.914786
R17761 VSS.n17849 VSS.n17284 0.914786
R17762 VSS.n17859 VSS.n17858 0.914786
R17763 VSS.n18534 VSS.n18307 0.914786
R17764 VSS.n18375 VSS.n18374 0.914786
R17765 VSS.n18499 VSS.n18357 0.914786
R17766 VSS.n18481 VSS.n18480 0.914786
R17767 VSS.n18479 VSS.n18421 0.914786
R17768 VSS.n18463 VSS.n18462 0.914786
R17769 VSS.n9764 VSS.n9749 0.914786
R17770 VSS.n9826 VSS.n9825 0.914786
R17771 VSS.n9827 VSS.n9359 0.914786
R17772 VSS.n9883 VSS.n9882 0.914786
R17773 VSS.n9900 VSS.n9335 0.914786
R17774 VSS.n9910 VSS.n9909 0.914786
R17775 VSS.n16707 VSS.n16692 0.914786
R17776 VSS.n16769 VSS.n16768 0.914786
R17777 VSS.n16770 VSS.n16301 0.914786
R17778 VSS.n16826 VSS.n16825 0.914786
R17779 VSS.n16843 VSS.n16277 0.914786
R17780 VSS.n16853 VSS.n16852 0.914786
R17781 VSS.n16114 VSS.n16099 0.914786
R17782 VSS.n16176 VSS.n16175 0.914786
R17783 VSS.n16177 VSS.n1473 0.914786
R17784 VSS.n16233 VSS.n16232 0.914786
R17785 VSS.n16250 VSS.n1449 0.914786
R17786 VSS.n16260 VSS.n16259 0.914786
R17787 VSS.n2299 VSS.n2072 0.914786
R17788 VSS.n2144 VSS.n2143 0.914786
R17789 VSS.n2145 VSS.n2125 0.914786
R17790 VSS.n2192 VSS.n2173 0.914786
R17791 VSS.n2233 VSS.n2232 0.914786
R17792 VSS.n2206 VSS.n2199 0.914786
R17793 VSS.n3255 VSS.n3240 0.914786
R17794 VSS.n3317 VSS.n3316 0.914786
R17795 VSS.n3318 VSS.n2850 0.914786
R17796 VSS.n3374 VSS.n3373 0.914786
R17797 VSS.n3391 VSS.n2826 0.914786
R17798 VSS.n3401 VSS.n3400 0.914786
R17799 VSS.n3847 VSS.n3832 0.914786
R17800 VSS.n3909 VSS.n3908 0.914786
R17801 VSS.n3910 VSS.n3442 0.914786
R17802 VSS.n3966 VSS.n3965 0.914786
R17803 VSS.n3983 VSS.n3418 0.914786
R17804 VSS.n3993 VSS.n3992 0.914786
R17805 VSS.n4439 VSS.n4424 0.914786
R17806 VSS.n4501 VSS.n4500 0.914786
R17807 VSS.n4502 VSS.n4034 0.914786
R17808 VSS.n4558 VSS.n4557 0.914786
R17809 VSS.n4575 VSS.n4010 0.914786
R17810 VSS.n4585 VSS.n4584 0.914786
R17811 VSS.n5031 VSS.n5016 0.914786
R17812 VSS.n5093 VSS.n5092 0.914786
R17813 VSS.n5094 VSS.n4626 0.914786
R17814 VSS.n5150 VSS.n5149 0.914786
R17815 VSS.n5167 VSS.n4602 0.914786
R17816 VSS.n5177 VSS.n5176 0.914786
R17817 VSS.n5264 VSS.n2668 0.914786
R17818 VSS.n2740 VSS.n2739 0.914786
R17819 VSS.n2741 VSS.n2721 0.914786
R17820 VSS.n2788 VSS.n2769 0.914786
R17821 VSS.n5198 VSS.n5197 0.914786
R17822 VSS.n2802 VSS.n2795 0.914786
R17823 VSS.n5837 VSS.n5629 0.914786
R17824 VSS.n5701 VSS.n5700 0.914786
R17825 VSS.n5702 VSS.n5682 0.914786
R17826 VSS.n5762 VSS.n5742 0.914786
R17827 VSS.n5771 VSS.n5770 0.914786
R17828 VSS.n18883 VSS.n18882 0.914786
R17829 VSS.n6429 VSS.n6202 0.914786
R17830 VSS.n6274 VSS.n6273 0.914786
R17831 VSS.n6275 VSS.n6255 0.914786
R17832 VSS.n6322 VSS.n6303 0.914786
R17833 VSS.n6363 VSS.n6362 0.914786
R17834 VSS.n6336 VSS.n6329 0.914786
R17835 VSS.n7988 VSS.n7973 0.914786
R17836 VSS.n8050 VSS.n8049 0.914786
R17837 VSS.n8051 VSS.n7583 0.914786
R17838 VSS.n8107 VSS.n8106 0.914786
R17839 VSS.n8124 VSS.n7559 0.914786
R17840 VSS.n8134 VSS.n8133 0.914786
R17841 VSS.n8580 VSS.n8565 0.914786
R17842 VSS.n8642 VSS.n8641 0.914786
R17843 VSS.n8643 VSS.n8175 0.914786
R17844 VSS.n8699 VSS.n8698 0.914786
R17845 VSS.n8716 VSS.n8151 0.914786
R17846 VSS.n8726 VSS.n8725 0.914786
R17847 VSS.n9172 VSS.n9157 0.914786
R17848 VSS.n9234 VSS.n9233 0.914786
R17849 VSS.n9235 VSS.n8767 0.914786
R17850 VSS.n9291 VSS.n9290 0.914786
R17851 VSS.n9308 VSS.n8743 0.914786
R17852 VSS.n9318 VSS.n9317 0.914786
R17853 VSS.n10356 VSS.n10341 0.914786
R17854 VSS.n10418 VSS.n10417 0.914786
R17855 VSS.n10419 VSS.n9951 0.914786
R17856 VSS.n10475 VSS.n10474 0.914786
R17857 VSS.n10492 VSS.n9927 0.914786
R17858 VSS.n10502 VSS.n10501 0.914786
R17859 VSS.n10948 VSS.n10933 0.914786
R17860 VSS.n11010 VSS.n11009 0.914786
R17861 VSS.n11011 VSS.n10543 0.914786
R17862 VSS.n11067 VSS.n11066 0.914786
R17863 VSS.n11084 VSS.n10519 0.914786
R17864 VSS.n11094 VSS.n11093 0.914786
R17865 VSS.n11540 VSS.n11525 0.914786
R17866 VSS.n11602 VSS.n11601 0.914786
R17867 VSS.n11603 VSS.n11135 0.914786
R17868 VSS.n11659 VSS.n11658 0.914786
R17869 VSS.n11676 VSS.n11111 0.914786
R17870 VSS.n11686 VSS.n11685 0.914786
R17871 VSS.n12132 VSS.n12117 0.914786
R17872 VSS.n12194 VSS.n12193 0.914786
R17873 VSS.n12195 VSS.n11727 0.914786
R17874 VSS.n12251 VSS.n12250 0.914786
R17875 VSS.n12268 VSS.n11703 0.914786
R17876 VSS.n12278 VSS.n12277 0.914786
R17877 VSS.n12724 VSS.n12709 0.914786
R17878 VSS.n12786 VSS.n12785 0.914786
R17879 VSS.n12787 VSS.n12319 0.914786
R17880 VSS.n12843 VSS.n12842 0.914786
R17881 VSS.n12860 VSS.n12295 0.914786
R17882 VSS.n12870 VSS.n12869 0.914786
R17883 VSS.n13316 VSS.n13301 0.914786
R17884 VSS.n13378 VSS.n13377 0.914786
R17885 VSS.n13379 VSS.n12911 0.914786
R17886 VSS.n13435 VSS.n13434 0.914786
R17887 VSS.n13452 VSS.n12887 0.914786
R17888 VSS.n13462 VSS.n13461 0.914786
R17889 VSS.n13908 VSS.n13893 0.914786
R17890 VSS.n13970 VSS.n13969 0.914786
R17891 VSS.n13971 VSS.n13503 0.914786
R17892 VSS.n14027 VSS.n14026 0.914786
R17893 VSS.n14044 VSS.n13479 0.914786
R17894 VSS.n14054 VSS.n14053 0.914786
R17895 VSS.n14500 VSS.n14485 0.914786
R17896 VSS.n14562 VSS.n14561 0.914786
R17897 VSS.n14563 VSS.n14095 0.914786
R17898 VSS.n14619 VSS.n14618 0.914786
R17899 VSS.n14636 VSS.n14071 0.914786
R17900 VSS.n14646 VSS.n14645 0.914786
R17901 VSS.n15092 VSS.n15077 0.914786
R17902 VSS.n15154 VSS.n15153 0.914786
R17903 VSS.n15155 VSS.n14687 0.914786
R17904 VSS.n15211 VSS.n15210 0.914786
R17905 VSS.n15228 VSS.n14663 0.914786
R17906 VSS.n15238 VSS.n15237 0.914786
R17907 VSS.n15684 VSS.n15669 0.914786
R17908 VSS.n15746 VSS.n15745 0.914786
R17909 VSS.n15747 VSS.n15279 0.914786
R17910 VSS.n15803 VSS.n15802 0.914786
R17911 VSS.n15820 VSS.n15255 0.914786
R17912 VSS.n15830 VSS.n15829 0.914786
R17913 VSS.n15917 VSS.n6808 0.914786
R17914 VSS.n6880 VSS.n6879 0.914786
R17915 VSS.n6881 VSS.n6861 0.914786
R17916 VSS.n6928 VSS.n6909 0.914786
R17917 VSS.n15851 VSS.n15850 0.914786
R17918 VSS.n6942 VSS.n6935 0.914786
R17919 VSS.n7396 VSS.n7381 0.914786
R17920 VSS.n7458 VSS.n7457 0.914786
R17921 VSS.n7459 VSS.n6990 0.914786
R17922 VSS.n7515 VSS.n7514 0.914786
R17923 VSS.n7532 VSS.n6966 0.914786
R17924 VSS.n7542 VSS.n7541 0.914786
R17925 VSS.n18708 VSS.n18693 0.914786
R17926 VSS.n18770 VSS.n18769 0.914786
R17927 VSS.n18771 VSS.n88 0.914786
R17928 VSS.n18827 VSS.n18826 0.914786
R17929 VSS.n18844 VSS.n64 0.914786
R17930 VSS.n18854 VSS.n18853 0.914786
R17931 VSS.n831 VSS.n631 0.914786
R17932 VSS.n703 VSS.n702 0.914786
R17933 VSS.n704 VSS.n684 0.914786
R17934 VSS.n764 VSS.n763 0.914786
R17935 VSS.n765 VSS.n48 0.914786
R17936 VSS.n18874 VSS.n43 0.914786
R17937 VSS.n17945 VSS.n1290 0.914786
R17938 VSS.n1362 VSS.n1361 0.914786
R17939 VSS.n1363 VSS.n1343 0.914786
R17940 VSS.n1410 VSS.n1391 0.914786
R17941 VSS.n17879 VSS.n17878 0.914786
R17942 VSS.n1424 VSS.n1417 0.914786
R17943 VSS.n17270 VSS.n16862 0.908949
R17944 VSS.n17862 VSS.n17276 0.908949
R17945 VSS.n18466 VSS.n18432 0.908949
R17946 VSS.n9913 VSS.n9327 0.908949
R17947 VSS.n16856 VSS.n16269 0.908949
R17948 VSS.n16263 VSS.n1441 0.908949
R17949 VSS.n2222 VSS.n2207 0.908949
R17950 VSS.n3404 VSS.n2818 0.908949
R17951 VSS.n3996 VSS.n3410 0.908949
R17952 VSS.n4588 VSS.n4002 0.908949
R17953 VSS.n5180 VSS.n4594 0.908949
R17954 VSS.n5187 VSS.n2803 0.908949
R17955 VSS.n18886 VSS.n3 0.908949
R17956 VSS.n6352 VSS.n6337 0.908949
R17957 VSS.n8137 VSS.n7551 0.908949
R17958 VSS.n8729 VSS.n8143 0.908949
R17959 VSS.n9321 VSS.n8735 0.908949
R17960 VSS.n10505 VSS.n9919 0.908949
R17961 VSS.n11097 VSS.n10511 0.908949
R17962 VSS.n11689 VSS.n11103 0.908949
R17963 VSS.n12281 VSS.n11695 0.908949
R17964 VSS.n12873 VSS.n12287 0.908949
R17965 VSS.n13465 VSS.n12879 0.908949
R17966 VSS.n14057 VSS.n13471 0.908949
R17967 VSS.n14649 VSS.n14063 0.908949
R17968 VSS.n15241 VSS.n14655 0.908949
R17969 VSS.n15833 VSS.n15247 0.908949
R17970 VSS.n15840 VSS.n6943 0.908949
R17971 VSS.n7545 VSS.n6958 0.908949
R17972 VSS.n18857 VSS.n56 0.908949
R17973 VSS.n18863 VSS.n44 0.908949
R17974 VSS.n17868 VSS.n1425 0.908949
R17975 VSS.n17110 VSS.n16931 0.908879
R17976 VSS.n17702 VSS.n17345 0.908879
R17977 VSS.n18326 VSS.n18308 0.908879
R17978 VSS.n9752 VSS.n9395 0.908879
R17979 VSS.n16695 VSS.n16337 0.908879
R17980 VSS.n16102 VSS.n1509 0.908879
R17981 VSS.n2090 VSS.n2073 0.908879
R17982 VSS.n3243 VSS.n2886 0.908879
R17983 VSS.n3835 VSS.n3478 0.908879
R17984 VSS.n4427 VSS.n4070 0.908879
R17985 VSS.n5019 VSS.n4662 0.908879
R17986 VSS.n2686 VSS.n2669 0.908879
R17987 VSS.n5647 VSS.n5630 0.908879
R17988 VSS.n6220 VSS.n6203 0.908879
R17989 VSS.n7976 VSS.n7619 0.908879
R17990 VSS.n8568 VSS.n8211 0.908879
R17991 VSS.n9160 VSS.n8803 0.908879
R17992 VSS.n10344 VSS.n9987 0.908879
R17993 VSS.n10936 VSS.n10579 0.908879
R17994 VSS.n11528 VSS.n11171 0.908879
R17995 VSS.n12120 VSS.n11763 0.908879
R17996 VSS.n12712 VSS.n12355 0.908879
R17997 VSS.n13304 VSS.n12947 0.908879
R17998 VSS.n13896 VSS.n13539 0.908879
R17999 VSS.n14488 VSS.n14131 0.908879
R18000 VSS.n15080 VSS.n14723 0.908879
R18001 VSS.n15672 VSS.n15315 0.908879
R18002 VSS.n6826 VSS.n6809 0.908879
R18003 VSS.n7384 VSS.n7026 0.908879
R18004 VSS.n18696 VSS.n124 0.908879
R18005 VSS.n649 VSS.n632 0.908879
R18006 VSS.n1308 VSS.n1291 0.908879
R18007 VSS.n17145 VSS.n16926 0.853
R18008 VSS.n17191 VSS.n16899 0.853
R18009 VSS.n16876 VSS.n16875 0.853
R18010 VSS.n17737 VSS.n17340 0.853
R18011 VSS.n17783 VSS.n17313 0.853
R18012 VSS.n17290 VSS.n17289 0.853
R18013 VSS.n18521 VSS.n18317 0.853
R18014 VSS.n18354 VSS.n18352 0.853
R18015 VSS.n18417 VSS.n18415 0.853
R18016 VSS.n9787 VSS.n9390 0.853
R18017 VSS.n9833 VSS.n9363 0.853
R18018 VSS.n9341 VSS.n9340 0.853
R18019 VSS.n16730 VSS.n16332 0.853
R18020 VSS.n16776 VSS.n16305 0.853
R18021 VSS.n16283 VSS.n16282 0.853
R18022 VSS.n16137 VSS.n1504 0.853
R18023 VSS.n16183 VSS.n1477 0.853
R18024 VSS.n1455 VSS.n1454 0.853
R18025 VSS.n2112 VSS.n2082 0.853
R18026 VSS.n2151 VSS.n2129 0.853
R18027 VSS.n2238 VSS.n2164 0.853
R18028 VSS.n3278 VSS.n2881 0.853
R18029 VSS.n3324 VSS.n2854 0.853
R18030 VSS.n2832 VSS.n2831 0.853
R18031 VSS.n3870 VSS.n3473 0.853
R18032 VSS.n3916 VSS.n3446 0.853
R18033 VSS.n3424 VSS.n3423 0.853
R18034 VSS.n4462 VSS.n4065 0.853
R18035 VSS.n4508 VSS.n4038 0.853
R18036 VSS.n4016 VSS.n4015 0.853
R18037 VSS.n5054 VSS.n4657 0.853
R18038 VSS.n5100 VSS.n4630 0.853
R18039 VSS.n4608 VSS.n4607 0.853
R18040 VSS.n2708 VSS.n2678 0.853
R18041 VSS.n2747 VSS.n2725 0.853
R18042 VSS.n5203 VSS.n2760 0.853
R18043 VSS.n5669 VSS.n5639 0.853
R18044 VSS.n5708 VSS.n5686 0.853
R18045 VSS.n5776 VSS.n5721 0.853
R18046 VSS.n6242 VSS.n6212 0.853
R18047 VSS.n6281 VSS.n6259 0.853
R18048 VSS.n6368 VSS.n6294 0.853
R18049 VSS.n8011 VSS.n7614 0.853
R18050 VSS.n8057 VSS.n7587 0.853
R18051 VSS.n7565 VSS.n7564 0.853
R18052 VSS.n8603 VSS.n8206 0.853
R18053 VSS.n8649 VSS.n8179 0.853
R18054 VSS.n8157 VSS.n8156 0.853
R18055 VSS.n9195 VSS.n8798 0.853
R18056 VSS.n9241 VSS.n8771 0.853
R18057 VSS.n8749 VSS.n8748 0.853
R18058 VSS.n10379 VSS.n9982 0.853
R18059 VSS.n10425 VSS.n9955 0.853
R18060 VSS.n9933 VSS.n9932 0.853
R18061 VSS.n10971 VSS.n10574 0.853
R18062 VSS.n11017 VSS.n10547 0.853
R18063 VSS.n10525 VSS.n10524 0.853
R18064 VSS.n11563 VSS.n11166 0.853
R18065 VSS.n11609 VSS.n11139 0.853
R18066 VSS.n11117 VSS.n11116 0.853
R18067 VSS.n12155 VSS.n11758 0.853
R18068 VSS.n12201 VSS.n11731 0.853
R18069 VSS.n11709 VSS.n11708 0.853
R18070 VSS.n12747 VSS.n12350 0.853
R18071 VSS.n12793 VSS.n12323 0.853
R18072 VSS.n12301 VSS.n12300 0.853
R18073 VSS.n13339 VSS.n12942 0.853
R18074 VSS.n13385 VSS.n12915 0.853
R18075 VSS.n12893 VSS.n12892 0.853
R18076 VSS.n13931 VSS.n13534 0.853
R18077 VSS.n13977 VSS.n13507 0.853
R18078 VSS.n13485 VSS.n13484 0.853
R18079 VSS.n14523 VSS.n14126 0.853
R18080 VSS.n14569 VSS.n14099 0.853
R18081 VSS.n14077 VSS.n14076 0.853
R18082 VSS.n15115 VSS.n14718 0.853
R18083 VSS.n15161 VSS.n14691 0.853
R18084 VSS.n14669 VSS.n14668 0.853
R18085 VSS.n15707 VSS.n15310 0.853
R18086 VSS.n15753 VSS.n15283 0.853
R18087 VSS.n15261 VSS.n15260 0.853
R18088 VSS.n6848 VSS.n6818 0.853
R18089 VSS.n6887 VSS.n6865 0.853
R18090 VSS.n15856 VSS.n6900 0.853
R18091 VSS.n7419 VSS.n7021 0.853
R18092 VSS.n7465 VSS.n6994 0.853
R18093 VSS.n6972 VSS.n6971 0.853
R18094 VSS.n18731 VSS.n119 0.853
R18095 VSS.n18777 VSS.n92 0.853
R18096 VSS.n70 VSS.n69 0.853
R18097 VSS.n671 VSS.n641 0.853
R18098 VSS.n710 VSS.n688 0.853
R18099 VSS.n770 VSS.n723 0.853
R18100 VSS.n1330 VSS.n1300 0.853
R18101 VSS.n1369 VSS.n1347 0.853
R18102 VSS.n17884 VSS.n1382 0.853
R18103 VSS.n17161 VSS.n16918 0.823357
R18104 VSS.n17170 VSS.n16910 0.823357
R18105 VSS.n17212 VSS.n16896 0.823357
R18106 VSS.n17222 VSS.n16883 0.823357
R18107 VSS.n17753 VSS.n17332 0.823357
R18108 VSS.n17762 VSS.n17324 0.823357
R18109 VSS.n17804 VSS.n17310 0.823357
R18110 VSS.n17814 VSS.n17297 0.823357
R18111 VSS.n18511 VSS.n18343 0.823357
R18112 VSS.n18510 VSS.n18509 0.823357
R18113 VSS.n18396 VSS.n18358 0.823357
R18114 VSS.n18441 VSS.n18387 0.823357
R18115 VSS.n9803 VSS.n9382 0.823357
R18116 VSS.n9812 VSS.n9374 0.823357
R18117 VSS.n9854 VSS.n9360 0.823357
R18118 VSS.n9864 VSS.n9347 0.823357
R18119 VSS.n16746 VSS.n16324 0.823357
R18120 VSS.n16755 VSS.n16316 0.823357
R18121 VSS.n16797 VSS.n16302 0.823357
R18122 VSS.n16807 VSS.n16289 0.823357
R18123 VSS.n16153 VSS.n1496 0.823357
R18124 VSS.n16162 VSS.n1488 0.823357
R18125 VSS.n16204 VSS.n1474 0.823357
R18126 VSS.n16214 VSS.n1461 0.823357
R18127 VSS.n2277 VSS.n2107 0.823357
R18128 VSS.n2269 VSS.n2119 0.823357
R18129 VSS.n2260 VSS.n2126 0.823357
R18130 VSS.n2249 VSS.n2248 0.823357
R18131 VSS.n3294 VSS.n2873 0.823357
R18132 VSS.n3303 VSS.n2865 0.823357
R18133 VSS.n3345 VSS.n2851 0.823357
R18134 VSS.n3355 VSS.n2838 0.823357
R18135 VSS.n3886 VSS.n3465 0.823357
R18136 VSS.n3895 VSS.n3457 0.823357
R18137 VSS.n3937 VSS.n3443 0.823357
R18138 VSS.n3947 VSS.n3430 0.823357
R18139 VSS.n4478 VSS.n4057 0.823357
R18140 VSS.n4487 VSS.n4049 0.823357
R18141 VSS.n4529 VSS.n4035 0.823357
R18142 VSS.n4539 VSS.n4022 0.823357
R18143 VSS.n5070 VSS.n4649 0.823357
R18144 VSS.n5079 VSS.n4641 0.823357
R18145 VSS.n5121 VSS.n4627 0.823357
R18146 VSS.n5131 VSS.n4614 0.823357
R18147 VSS.n5242 VSS.n2703 0.823357
R18148 VSS.n5234 VSS.n2715 0.823357
R18149 VSS.n5225 VSS.n2722 0.823357
R18150 VSS.n5214 VSS.n5213 0.823357
R18151 VSS.n5815 VSS.n5664 0.823357
R18152 VSS.n5807 VSS.n5676 0.823357
R18153 VSS.n5798 VSS.n5683 0.823357
R18154 VSS.n5787 VSS.n5786 0.823357
R18155 VSS.n6407 VSS.n6237 0.823357
R18156 VSS.n6399 VSS.n6249 0.823357
R18157 VSS.n6390 VSS.n6256 0.823357
R18158 VSS.n6379 VSS.n6378 0.823357
R18159 VSS.n8027 VSS.n7606 0.823357
R18160 VSS.n8036 VSS.n7598 0.823357
R18161 VSS.n8078 VSS.n7584 0.823357
R18162 VSS.n8088 VSS.n7571 0.823357
R18163 VSS.n8619 VSS.n8198 0.823357
R18164 VSS.n8628 VSS.n8190 0.823357
R18165 VSS.n8670 VSS.n8176 0.823357
R18166 VSS.n8680 VSS.n8163 0.823357
R18167 VSS.n9211 VSS.n8790 0.823357
R18168 VSS.n9220 VSS.n8782 0.823357
R18169 VSS.n9262 VSS.n8768 0.823357
R18170 VSS.n9272 VSS.n8755 0.823357
R18171 VSS.n10395 VSS.n9974 0.823357
R18172 VSS.n10404 VSS.n9966 0.823357
R18173 VSS.n10446 VSS.n9952 0.823357
R18174 VSS.n10456 VSS.n9939 0.823357
R18175 VSS.n10987 VSS.n10566 0.823357
R18176 VSS.n10996 VSS.n10558 0.823357
R18177 VSS.n11038 VSS.n10544 0.823357
R18178 VSS.n11048 VSS.n10531 0.823357
R18179 VSS.n11579 VSS.n11158 0.823357
R18180 VSS.n11588 VSS.n11150 0.823357
R18181 VSS.n11630 VSS.n11136 0.823357
R18182 VSS.n11640 VSS.n11123 0.823357
R18183 VSS.n12171 VSS.n11750 0.823357
R18184 VSS.n12180 VSS.n11742 0.823357
R18185 VSS.n12222 VSS.n11728 0.823357
R18186 VSS.n12232 VSS.n11715 0.823357
R18187 VSS.n12763 VSS.n12342 0.823357
R18188 VSS.n12772 VSS.n12334 0.823357
R18189 VSS.n12814 VSS.n12320 0.823357
R18190 VSS.n12824 VSS.n12307 0.823357
R18191 VSS.n13355 VSS.n12934 0.823357
R18192 VSS.n13364 VSS.n12926 0.823357
R18193 VSS.n13406 VSS.n12912 0.823357
R18194 VSS.n13416 VSS.n12899 0.823357
R18195 VSS.n13947 VSS.n13526 0.823357
R18196 VSS.n13956 VSS.n13518 0.823357
R18197 VSS.n13998 VSS.n13504 0.823357
R18198 VSS.n14008 VSS.n13491 0.823357
R18199 VSS.n14539 VSS.n14118 0.823357
R18200 VSS.n14548 VSS.n14110 0.823357
R18201 VSS.n14590 VSS.n14096 0.823357
R18202 VSS.n14600 VSS.n14083 0.823357
R18203 VSS.n15131 VSS.n14710 0.823357
R18204 VSS.n15140 VSS.n14702 0.823357
R18205 VSS.n15182 VSS.n14688 0.823357
R18206 VSS.n15192 VSS.n14675 0.823357
R18207 VSS.n15723 VSS.n15302 0.823357
R18208 VSS.n15732 VSS.n15294 0.823357
R18209 VSS.n15774 VSS.n15280 0.823357
R18210 VSS.n15784 VSS.n15267 0.823357
R18211 VSS.n15895 VSS.n6843 0.823357
R18212 VSS.n15887 VSS.n6855 0.823357
R18213 VSS.n15878 VSS.n6862 0.823357
R18214 VSS.n15867 VSS.n15866 0.823357
R18215 VSS.n7435 VSS.n7013 0.823357
R18216 VSS.n7444 VSS.n7005 0.823357
R18217 VSS.n7486 VSS.n6991 0.823357
R18218 VSS.n7496 VSS.n6978 0.823357
R18219 VSS.n18747 VSS.n111 0.823357
R18220 VSS.n18756 VSS.n103 0.823357
R18221 VSS.n18798 VSS.n89 0.823357
R18222 VSS.n18808 VSS.n76 0.823357
R18223 VSS.n809 VSS.n666 0.823357
R18224 VSS.n801 VSS.n678 0.823357
R18225 VSS.n792 VSS.n685 0.823357
R18226 VSS.n781 VSS.n780 0.823357
R18227 VSS.n17923 VSS.n1325 0.823357
R18228 VSS.n17915 VSS.n1337 0.823357
R18229 VSS.n17906 VSS.n1344 0.823357
R18230 VSS.n17895 VSS.n17894 0.823357
R18231 VSS.n16918 VSS.n16910 0.731929
R18232 VSS.n17222 VSS.n17221 0.731929
R18233 VSS.n17234 VSS.n16883 0.731929
R18234 VSS.n17332 VSS.n17324 0.731929
R18235 VSS.n17814 VSS.n17813 0.731929
R18236 VSS.n17826 VSS.n17297 0.731929
R18237 VSS.n18511 VSS.n18510 0.731929
R18238 VSS.n18490 VSS.n18387 0.731929
R18239 VSS.n18448 VSS.n18441 0.731929
R18240 VSS.n9382 VSS.n9374 0.731929
R18241 VSS.n9864 VSS.n9863 0.731929
R18242 VSS.n9876 VSS.n9347 0.731929
R18243 VSS.n16324 VSS.n16316 0.731929
R18244 VSS.n16807 VSS.n16806 0.731929
R18245 VSS.n16819 VSS.n16289 0.731929
R18246 VSS.n1496 VSS.n1488 0.731929
R18247 VSS.n16214 VSS.n16213 0.731929
R18248 VSS.n16226 VSS.n1461 0.731929
R18249 VSS.n2119 VSS.n2107 0.731929
R18250 VSS.n2250 VSS.n2249 0.731929
R18251 VSS.n2248 VSS.n2158 0.731929
R18252 VSS.n2873 VSS.n2865 0.731929
R18253 VSS.n3355 VSS.n3354 0.731929
R18254 VSS.n3367 VSS.n2838 0.731929
R18255 VSS.n3465 VSS.n3457 0.731929
R18256 VSS.n3947 VSS.n3946 0.731929
R18257 VSS.n3959 VSS.n3430 0.731929
R18258 VSS.n4057 VSS.n4049 0.731929
R18259 VSS.n4539 VSS.n4538 0.731929
R18260 VSS.n4551 VSS.n4022 0.731929
R18261 VSS.n4649 VSS.n4641 0.731929
R18262 VSS.n5131 VSS.n5130 0.731929
R18263 VSS.n5143 VSS.n4614 0.731929
R18264 VSS.n2715 VSS.n2703 0.731929
R18265 VSS.n5215 VSS.n5214 0.731929
R18266 VSS.n5213 VSS.n2754 0.731929
R18267 VSS.n5676 VSS.n5664 0.731929
R18268 VSS.n5788 VSS.n5787 0.731929
R18269 VSS.n5786 VSS.n5715 0.731929
R18270 VSS.n6249 VSS.n6237 0.731929
R18271 VSS.n6380 VSS.n6379 0.731929
R18272 VSS.n6378 VSS.n6288 0.731929
R18273 VSS.n7606 VSS.n7598 0.731929
R18274 VSS.n8088 VSS.n8087 0.731929
R18275 VSS.n8100 VSS.n7571 0.731929
R18276 VSS.n8198 VSS.n8190 0.731929
R18277 VSS.n8680 VSS.n8679 0.731929
R18278 VSS.n8692 VSS.n8163 0.731929
R18279 VSS.n8790 VSS.n8782 0.731929
R18280 VSS.n9272 VSS.n9271 0.731929
R18281 VSS.n9284 VSS.n8755 0.731929
R18282 VSS.n9974 VSS.n9966 0.731929
R18283 VSS.n10456 VSS.n10455 0.731929
R18284 VSS.n10468 VSS.n9939 0.731929
R18285 VSS.n10566 VSS.n10558 0.731929
R18286 VSS.n11048 VSS.n11047 0.731929
R18287 VSS.n11060 VSS.n10531 0.731929
R18288 VSS.n11158 VSS.n11150 0.731929
R18289 VSS.n11640 VSS.n11639 0.731929
R18290 VSS.n11652 VSS.n11123 0.731929
R18291 VSS.n11750 VSS.n11742 0.731929
R18292 VSS.n12232 VSS.n12231 0.731929
R18293 VSS.n12244 VSS.n11715 0.731929
R18294 VSS.n12342 VSS.n12334 0.731929
R18295 VSS.n12824 VSS.n12823 0.731929
R18296 VSS.n12836 VSS.n12307 0.731929
R18297 VSS.n12934 VSS.n12926 0.731929
R18298 VSS.n13416 VSS.n13415 0.731929
R18299 VSS.n13428 VSS.n12899 0.731929
R18300 VSS.n13526 VSS.n13518 0.731929
R18301 VSS.n14008 VSS.n14007 0.731929
R18302 VSS.n14020 VSS.n13491 0.731929
R18303 VSS.n14118 VSS.n14110 0.731929
R18304 VSS.n14600 VSS.n14599 0.731929
R18305 VSS.n14612 VSS.n14083 0.731929
R18306 VSS.n14710 VSS.n14702 0.731929
R18307 VSS.n15192 VSS.n15191 0.731929
R18308 VSS.n15204 VSS.n14675 0.731929
R18309 VSS.n15302 VSS.n15294 0.731929
R18310 VSS.n15784 VSS.n15783 0.731929
R18311 VSS.n15796 VSS.n15267 0.731929
R18312 VSS.n6855 VSS.n6843 0.731929
R18313 VSS.n15868 VSS.n15867 0.731929
R18314 VSS.n15866 VSS.n6894 0.731929
R18315 VSS.n7013 VSS.n7005 0.731929
R18316 VSS.n7496 VSS.n7495 0.731929
R18317 VSS.n7508 VSS.n6978 0.731929
R18318 VSS.n111 VSS.n103 0.731929
R18319 VSS.n18808 VSS.n18807 0.731929
R18320 VSS.n18820 VSS.n76 0.731929
R18321 VSS.n678 VSS.n666 0.731929
R18322 VSS.n782 VSS.n781 0.731929
R18323 VSS.n780 VSS.n717 0.731929
R18324 VSS.n1337 VSS.n1325 0.731929
R18325 VSS.n17896 VSS.n17895 0.731929
R18326 VSS.n17894 VSS.n1376 0.731929
R18327 VSS VSS.n7548 0.680647
R18328 VSS.n12284 VSS 0.680647
R18329 VSS VSS.n0 0.680647
R18330 VSS VSS.n16266 0.680647
R18331 VSS.n17114 VSS.n17107 0.6405
R18332 VSS.n17183 VSS.n16904 0.6405
R18333 VSS.n17241 VSS.n16870 0.6405
R18334 VSS.n17267 VSS.n16864 0.6405
R18335 VSS.n17706 VSS.n17699 0.6405
R18336 VSS.n17775 VSS.n17318 0.6405
R18337 VSS.n17833 VSS.n17284 0.6405
R18338 VSS.n17859 VSS.n17278 0.6405
R18339 VSS.n18322 VSS.n18307 0.6405
R18340 VSS.n18379 VSS.n18374 0.6405
R18341 VSS.n18480 VSS.n18479 0.6405
R18342 VSS.n18463 VSS.n18435 0.6405
R18343 VSS.n9756 VSS.n9749 0.6405
R18344 VSS.n9825 VSS.n9368 0.6405
R18345 VSS.n9883 VSS.n9335 0.6405
R18346 VSS.n9910 VSS.n9329 0.6405
R18347 VSS.n16699 VSS.n16692 0.6405
R18348 VSS.n16768 VSS.n16310 0.6405
R18349 VSS.n16826 VSS.n16277 0.6405
R18350 VSS.n16853 VSS.n16271 0.6405
R18351 VSS.n16106 VSS.n16099 0.6405
R18352 VSS.n16175 VSS.n1482 0.6405
R18353 VSS.n16233 VSS.n1449 0.6405
R18354 VSS.n16260 VSS.n1443 0.6405
R18355 VSS.n2086 VSS.n2072 0.6405
R18356 VSS.n2143 VSS.n2121 0.6405
R18357 VSS.n2233 VSS.n2173 0.6405
R18358 VSS.n2225 VSS.n2199 0.6405
R18359 VSS.n3247 VSS.n3240 0.6405
R18360 VSS.n3316 VSS.n2859 0.6405
R18361 VSS.n3374 VSS.n2826 0.6405
R18362 VSS.n3401 VSS.n2820 0.6405
R18363 VSS.n3839 VSS.n3832 0.6405
R18364 VSS.n3908 VSS.n3451 0.6405
R18365 VSS.n3966 VSS.n3418 0.6405
R18366 VSS.n3993 VSS.n3412 0.6405
R18367 VSS.n4431 VSS.n4424 0.6405
R18368 VSS.n4500 VSS.n4043 0.6405
R18369 VSS.n4558 VSS.n4010 0.6405
R18370 VSS.n4585 VSS.n4004 0.6405
R18371 VSS.n5023 VSS.n5016 0.6405
R18372 VSS.n5092 VSS.n4635 0.6405
R18373 VSS.n5150 VSS.n4602 0.6405
R18374 VSS.n5177 VSS.n4596 0.6405
R18375 VSS.n2682 VSS.n2668 0.6405
R18376 VSS.n2739 VSS.n2717 0.6405
R18377 VSS.n5198 VSS.n2769 0.6405
R18378 VSS.n5190 VSS.n2795 0.6405
R18379 VSS.n5643 VSS.n5629 0.6405
R18380 VSS.n5700 VSS.n5678 0.6405
R18381 VSS.n5771 VSS.n5742 0.6405
R18382 VSS.n18883 VSS.n5 0.6405
R18383 VSS.n6216 VSS.n6202 0.6405
R18384 VSS.n6273 VSS.n6251 0.6405
R18385 VSS.n6363 VSS.n6303 0.6405
R18386 VSS.n6355 VSS.n6329 0.6405
R18387 VSS.n7980 VSS.n7973 0.6405
R18388 VSS.n8049 VSS.n7592 0.6405
R18389 VSS.n8107 VSS.n7559 0.6405
R18390 VSS.n8134 VSS.n7553 0.6405
R18391 VSS.n8572 VSS.n8565 0.6405
R18392 VSS.n8641 VSS.n8184 0.6405
R18393 VSS.n8699 VSS.n8151 0.6405
R18394 VSS.n8726 VSS.n8145 0.6405
R18395 VSS.n9164 VSS.n9157 0.6405
R18396 VSS.n9233 VSS.n8776 0.6405
R18397 VSS.n9291 VSS.n8743 0.6405
R18398 VSS.n9318 VSS.n8737 0.6405
R18399 VSS.n10348 VSS.n10341 0.6405
R18400 VSS.n10417 VSS.n9960 0.6405
R18401 VSS.n10475 VSS.n9927 0.6405
R18402 VSS.n10502 VSS.n9921 0.6405
R18403 VSS.n10940 VSS.n10933 0.6405
R18404 VSS.n11009 VSS.n10552 0.6405
R18405 VSS.n11067 VSS.n10519 0.6405
R18406 VSS.n11094 VSS.n10513 0.6405
R18407 VSS.n11532 VSS.n11525 0.6405
R18408 VSS.n11601 VSS.n11144 0.6405
R18409 VSS.n11659 VSS.n11111 0.6405
R18410 VSS.n11686 VSS.n11105 0.6405
R18411 VSS.n12124 VSS.n12117 0.6405
R18412 VSS.n12193 VSS.n11736 0.6405
R18413 VSS.n12251 VSS.n11703 0.6405
R18414 VSS.n12278 VSS.n11697 0.6405
R18415 VSS.n12716 VSS.n12709 0.6405
R18416 VSS.n12785 VSS.n12328 0.6405
R18417 VSS.n12843 VSS.n12295 0.6405
R18418 VSS.n12870 VSS.n12289 0.6405
R18419 VSS.n13308 VSS.n13301 0.6405
R18420 VSS.n13377 VSS.n12920 0.6405
R18421 VSS.n13435 VSS.n12887 0.6405
R18422 VSS.n13462 VSS.n12881 0.6405
R18423 VSS.n13900 VSS.n13893 0.6405
R18424 VSS.n13969 VSS.n13512 0.6405
R18425 VSS.n14027 VSS.n13479 0.6405
R18426 VSS.n14054 VSS.n13473 0.6405
R18427 VSS.n14492 VSS.n14485 0.6405
R18428 VSS.n14561 VSS.n14104 0.6405
R18429 VSS.n14619 VSS.n14071 0.6405
R18430 VSS.n14646 VSS.n14065 0.6405
R18431 VSS.n15084 VSS.n15077 0.6405
R18432 VSS.n15153 VSS.n14696 0.6405
R18433 VSS.n15211 VSS.n14663 0.6405
R18434 VSS.n15238 VSS.n14657 0.6405
R18435 VSS.n15676 VSS.n15669 0.6405
R18436 VSS.n15745 VSS.n15288 0.6405
R18437 VSS.n15803 VSS.n15255 0.6405
R18438 VSS.n15830 VSS.n15249 0.6405
R18439 VSS.n6822 VSS.n6808 0.6405
R18440 VSS.n6879 VSS.n6857 0.6405
R18441 VSS.n15851 VSS.n6909 0.6405
R18442 VSS.n15843 VSS.n6935 0.6405
R18443 VSS.n7388 VSS.n7381 0.6405
R18444 VSS.n7457 VSS.n6999 0.6405
R18445 VSS.n7515 VSS.n6966 0.6405
R18446 VSS.n7542 VSS.n6960 0.6405
R18447 VSS.n18700 VSS.n18693 0.6405
R18448 VSS.n18769 VSS.n97 0.6405
R18449 VSS.n18827 VSS.n64 0.6405
R18450 VSS.n18854 VSS.n58 0.6405
R18451 VSS.n645 VSS.n631 0.6405
R18452 VSS.n702 VSS.n680 0.6405
R18453 VSS.n765 VSS.n764 0.6405
R18454 VSS.n18866 VSS.n43 0.6405
R18455 VSS.n1304 VSS.n1290 0.6405
R18456 VSS.n1361 VSS.n1339 0.6405
R18457 VSS.n17879 VSS.n1391 0.6405
R18458 VSS.n17871 VSS.n1417 0.6405
R18459 VSS.n17151 VSS.n17150 0.549071
R18460 VSS.n17200 VSS.n16891 0.549071
R18461 VSS.n17743 VSS.n17742 0.549071
R18462 VSS.n17792 VSS.n17305 0.549071
R18463 VSS.n18364 VSS.n18313 0.549071
R18464 VSS.n18405 VSS.n18386 0.549071
R18465 VSS.n9793 VSS.n9792 0.549071
R18466 VSS.n9842 VSS.n9355 0.549071
R18467 VSS.n16736 VSS.n16735 0.549071
R18468 VSS.n16785 VSS.n16297 0.549071
R18469 VSS.n16143 VSS.n16142 0.549071
R18470 VSS.n16192 VSS.n1469 0.549071
R18471 VSS.n2285 VSS.n2078 0.549071
R18472 VSS.n2185 VSS.n2178 0.549071
R18473 VSS.n3284 VSS.n3283 0.549071
R18474 VSS.n3333 VSS.n2846 0.549071
R18475 VSS.n3876 VSS.n3875 0.549071
R18476 VSS.n3925 VSS.n3438 0.549071
R18477 VSS.n4468 VSS.n4467 0.549071
R18478 VSS.n4517 VSS.n4030 0.549071
R18479 VSS.n5060 VSS.n5059 0.549071
R18480 VSS.n5109 VSS.n4622 0.549071
R18481 VSS.n5250 VSS.n2674 0.549071
R18482 VSS.n2781 VSS.n2774 0.549071
R18483 VSS.n5823 VSS.n5635 0.549071
R18484 VSS.n5755 VSS.n5748 0.549071
R18485 VSS.n6415 VSS.n6208 0.549071
R18486 VSS.n6315 VSS.n6308 0.549071
R18487 VSS.n8017 VSS.n8016 0.549071
R18488 VSS.n8066 VSS.n7579 0.549071
R18489 VSS.n8609 VSS.n8608 0.549071
R18490 VSS.n8658 VSS.n8171 0.549071
R18491 VSS.n9201 VSS.n9200 0.549071
R18492 VSS.n9250 VSS.n8763 0.549071
R18493 VSS.n10385 VSS.n10384 0.549071
R18494 VSS.n10434 VSS.n9947 0.549071
R18495 VSS.n10977 VSS.n10976 0.549071
R18496 VSS.n11026 VSS.n10539 0.549071
R18497 VSS.n11569 VSS.n11568 0.549071
R18498 VSS.n11618 VSS.n11131 0.549071
R18499 VSS.n12161 VSS.n12160 0.549071
R18500 VSS.n12210 VSS.n11723 0.549071
R18501 VSS.n12753 VSS.n12752 0.549071
R18502 VSS.n12802 VSS.n12315 0.549071
R18503 VSS.n13345 VSS.n13344 0.549071
R18504 VSS.n13394 VSS.n12907 0.549071
R18505 VSS.n13937 VSS.n13936 0.549071
R18506 VSS.n13986 VSS.n13499 0.549071
R18507 VSS.n14529 VSS.n14528 0.549071
R18508 VSS.n14578 VSS.n14091 0.549071
R18509 VSS.n15121 VSS.n15120 0.549071
R18510 VSS.n15170 VSS.n14683 0.549071
R18511 VSS.n15713 VSS.n15712 0.549071
R18512 VSS.n15762 VSS.n15275 0.549071
R18513 VSS.n15903 VSS.n6814 0.549071
R18514 VSS.n6921 VSS.n6914 0.549071
R18515 VSS.n7425 VSS.n7424 0.549071
R18516 VSS.n7474 VSS.n6986 0.549071
R18517 VSS.n18737 VSS.n18736 0.549071
R18518 VSS.n18786 VSS.n84 0.549071
R18519 VSS.n817 VSS.n637 0.549071
R18520 VSS.n753 VSS.n746 0.549071
R18521 VSS.n17931 VSS.n1296 0.549071
R18522 VSS.n1403 VSS.n1396 0.549071
R18523 VSS.n9916 VSS 0.533588
R18524 VSS.n17134 VSS 0.517836
R18525 VSS.n17726 VSS 0.517836
R18526 VSS.n18328 VSS 0.517836
R18527 VSS.n9776 VSS 0.517836
R18528 VSS.n16719 VSS 0.517836
R18529 VSS.n16126 VSS 0.517836
R18530 VSS.n2092 VSS 0.517836
R18531 VSS.n3267 VSS 0.517836
R18532 VSS.n3859 VSS 0.517836
R18533 VSS.n4451 VSS 0.517836
R18534 VSS.n5043 VSS 0.517836
R18535 VSS.n2688 VSS 0.517836
R18536 VSS.n5649 VSS 0.517836
R18537 VSS.n6222 VSS 0.517836
R18538 VSS.n8000 VSS 0.517836
R18539 VSS.n8592 VSS 0.517836
R18540 VSS.n9184 VSS 0.517836
R18541 VSS.n10368 VSS 0.517836
R18542 VSS.n10960 VSS 0.517836
R18543 VSS.n11552 VSS 0.517836
R18544 VSS.n12144 VSS 0.517836
R18545 VSS.n12736 VSS 0.517836
R18546 VSS.n13328 VSS 0.517836
R18547 VSS.n13920 VSS 0.517836
R18548 VSS.n14512 VSS 0.517836
R18549 VSS.n15104 VSS 0.517836
R18550 VSS.n15696 VSS 0.517836
R18551 VSS.n6828 VSS 0.517836
R18552 VSS.n7408 VSS 0.517836
R18553 VSS.n18720 VSS 0.517836
R18554 VSS.n651 VSS 0.517836
R18555 VSS.n1310 VSS 0.517836
R18556 VSS.n17993 VSS.n1158 0.465127
R18557 VSS.n18042 VSS.n1023 0.465127
R18558 VSS.n17006 VSS.n17005 0.465127
R18559 VSS.n17501 VSS.n17500 0.465127
R18560 VSS.n17420 VSS.n17419 0.465127
R18561 VSS.n18582 VSS.n211 0.465127
R18562 VSS.n18078 VSS.n18077 0.465127
R18563 VSS.n9470 VSS.n9469 0.465127
R18564 VSS.n9551 VSS.n9550 0.465127
R18565 VSS.n16412 VSS.n16411 0.465127
R18566 VSS.n16487 VSS.n16486 0.465127
R18567 VSS.n1754 VSS.n1577 0.465127
R18568 VSS.n1652 VSS.n1651 0.465127
R18569 VSS.n2347 VSS.n1761 0.465127
R18570 VSS.n1843 VSS.n1842 0.465127
R18571 VSS.n2961 VSS.n2960 0.465127
R18572 VSS.n3042 VSS.n3041 0.465127
R18573 VSS.n3553 VSS.n3552 0.465127
R18574 VSS.n3634 VSS.n3633 0.465127
R18575 VSS.n4145 VSS.n4144 0.465127
R18576 VSS.n4226 VSS.n4225 0.465127
R18577 VSS.n4737 VSS.n4736 0.465127
R18578 VSS.n4818 VSS.n4817 0.465127
R18579 VSS.n5312 VSS.n2357 0.465127
R18580 VSS.n2439 VSS.n2438 0.465127
R18581 VSS.n5885 VSS.n5318 0.465127
R18582 VSS.n5400 VSS.n5399 0.465127
R18583 VSS.n6477 VSS.n5891 0.465127
R18584 VSS.n5973 VSS.n5972 0.465127
R18585 VSS.n7694 VSS.n7693 0.465127
R18586 VSS.n7775 VSS.n7774 0.465127
R18587 VSS.n8286 VSS.n8285 0.465127
R18588 VSS.n8367 VSS.n8366 0.465127
R18589 VSS.n8878 VSS.n8877 0.465127
R18590 VSS.n8959 VSS.n8958 0.465127
R18591 VSS.n10062 VSS.n10061 0.465127
R18592 VSS.n10143 VSS.n10142 0.465127
R18593 VSS.n10654 VSS.n10653 0.465127
R18594 VSS.n10735 VSS.n10734 0.465127
R18595 VSS.n11246 VSS.n11245 0.465127
R18596 VSS.n11327 VSS.n11326 0.465127
R18597 VSS.n11838 VSS.n11837 0.465127
R18598 VSS.n11919 VSS.n11918 0.465127
R18599 VSS.n12430 VSS.n12429 0.465127
R18600 VSS.n12511 VSS.n12510 0.465127
R18601 VSS.n13022 VSS.n13021 0.465127
R18602 VSS.n13103 VSS.n13102 0.465127
R18603 VSS.n13614 VSS.n13613 0.465127
R18604 VSS.n13695 VSS.n13694 0.465127
R18605 VSS.n14206 VSS.n14205 0.465127
R18606 VSS.n14287 VSS.n14286 0.465127
R18607 VSS.n14798 VSS.n14797 0.465127
R18608 VSS.n14879 VSS.n14878 0.465127
R18609 VSS.n15390 VSS.n15389 0.465127
R18610 VSS.n15471 VSS.n15470 0.465127
R18611 VSS.n15965 VSS.n6497 0.465127
R18612 VSS.n6579 VSS.n6578 0.465127
R18613 VSS.n7101 VSS.n7100 0.465127
R18614 VSS.n7176 VSS.n7175 0.465127
R18615 VSS.n203 VSS.n192 0.465127
R18616 VSS.n451 VSS.n290 0.465127
R18617 VSS.n557 VSS.n497 0.465127
R18618 VSS.n1016 VSS.n456 0.465127
R18619 VSS.n17953 VSS.n1197 0.457643
R18620 VSS.n18002 VSS.n1063 0.457643
R18621 VSS.n17116 VSS.n17115 0.457643
R18622 VSS.n17259 VSS.n17258 0.457643
R18623 VSS.n17130 VSS.n16936 0.457643
R18624 VSS.n17596 VSS.n17425 0.457643
R18625 VSS.n17708 VSS.n17707 0.457643
R18626 VSS.n17851 VSS.n17850 0.457643
R18627 VSS.n17722 VSS.n17350 0.457643
R18628 VSS.n18542 VSS.n18214 0.457643
R18629 VSS.n18528 VSS.n18312 0.457643
R18630 VSS.n18455 VSS.n18454 0.457643
R18631 VSS.n18173 VSS.n217 0.457643
R18632 VSS.n9772 VSS.n9400 0.457643
R18633 VSS.n9758 VSS.n9757 0.457643
R18634 VSS.n9902 VSS.n9901 0.457643
R18635 VSS.n9646 VSS.n9475 0.457643
R18636 VSS.n16715 VSS.n16342 0.457643
R18637 VSS.n16701 VSS.n16700 0.457643
R18638 VSS.n16845 VSS.n16844 0.457643
R18639 VSS.n16589 VSS.n16417 0.457643
R18640 VSS.n16122 VSS.n1514 0.457643
R18641 VSS.n16108 VSS.n16107 0.457643
R18642 VSS.n16252 VSS.n16251 0.457643
R18643 VSS.n15996 VSS.n1582 0.457643
R18644 VSS.n2307 VSS.n1979 0.457643
R18645 VSS.n2293 VSS.n2077 0.457643
R18646 VSS.n2226 VSS.n2174 0.457643
R18647 VSS.n1938 VSS.n1767 0.457643
R18648 VSS.n3263 VSS.n2891 0.457643
R18649 VSS.n3249 VSS.n3248 0.457643
R18650 VSS.n3393 VSS.n3392 0.457643
R18651 VSS.n3137 VSS.n2966 0.457643
R18652 VSS.n3855 VSS.n3483 0.457643
R18653 VSS.n3841 VSS.n3840 0.457643
R18654 VSS.n3985 VSS.n3984 0.457643
R18655 VSS.n3729 VSS.n3558 0.457643
R18656 VSS.n4447 VSS.n4075 0.457643
R18657 VSS.n4433 VSS.n4432 0.457643
R18658 VSS.n4577 VSS.n4576 0.457643
R18659 VSS.n4321 VSS.n4150 0.457643
R18660 VSS.n5039 VSS.n4667 0.457643
R18661 VSS.n5025 VSS.n5024 0.457643
R18662 VSS.n5169 VSS.n5168 0.457643
R18663 VSS.n4913 VSS.n4742 0.457643
R18664 VSS.n5272 VSS.n2575 0.457643
R18665 VSS.n5258 VSS.n2673 0.457643
R18666 VSS.n5191 VSS.n2770 0.457643
R18667 VSS.n2534 VSS.n2363 0.457643
R18668 VSS.n5845 VSS.n5536 0.457643
R18669 VSS.n5831 VSS.n5634 0.457643
R18670 VSS.n5744 VSS.n5743 0.457643
R18671 VSS.n5495 VSS.n5324 0.457643
R18672 VSS.n6437 VSS.n6109 0.457643
R18673 VSS.n6423 VSS.n6207 0.457643
R18674 VSS.n6356 VSS.n6304 0.457643
R18675 VSS.n6068 VSS.n5897 0.457643
R18676 VSS.n7996 VSS.n7624 0.457643
R18677 VSS.n7982 VSS.n7981 0.457643
R18678 VSS.n8126 VSS.n8125 0.457643
R18679 VSS.n7870 VSS.n7699 0.457643
R18680 VSS.n8588 VSS.n8216 0.457643
R18681 VSS.n8574 VSS.n8573 0.457643
R18682 VSS.n8718 VSS.n8717 0.457643
R18683 VSS.n8462 VSS.n8291 0.457643
R18684 VSS.n9180 VSS.n8808 0.457643
R18685 VSS.n9166 VSS.n9165 0.457643
R18686 VSS.n9310 VSS.n9309 0.457643
R18687 VSS.n9054 VSS.n8883 0.457643
R18688 VSS.n10364 VSS.n9992 0.457643
R18689 VSS.n10350 VSS.n10349 0.457643
R18690 VSS.n10494 VSS.n10493 0.457643
R18691 VSS.n10238 VSS.n10067 0.457643
R18692 VSS.n10956 VSS.n10584 0.457643
R18693 VSS.n10942 VSS.n10941 0.457643
R18694 VSS.n11086 VSS.n11085 0.457643
R18695 VSS.n10830 VSS.n10659 0.457643
R18696 VSS.n11548 VSS.n11176 0.457643
R18697 VSS.n11534 VSS.n11533 0.457643
R18698 VSS.n11678 VSS.n11677 0.457643
R18699 VSS.n11422 VSS.n11251 0.457643
R18700 VSS.n12140 VSS.n11768 0.457643
R18701 VSS.n12126 VSS.n12125 0.457643
R18702 VSS.n12270 VSS.n12269 0.457643
R18703 VSS.n12014 VSS.n11843 0.457643
R18704 VSS.n12732 VSS.n12360 0.457643
R18705 VSS.n12718 VSS.n12717 0.457643
R18706 VSS.n12862 VSS.n12861 0.457643
R18707 VSS.n12606 VSS.n12435 0.457643
R18708 VSS.n13324 VSS.n12952 0.457643
R18709 VSS.n13310 VSS.n13309 0.457643
R18710 VSS.n13454 VSS.n13453 0.457643
R18711 VSS.n13198 VSS.n13027 0.457643
R18712 VSS.n13916 VSS.n13544 0.457643
R18713 VSS.n13902 VSS.n13901 0.457643
R18714 VSS.n14046 VSS.n14045 0.457643
R18715 VSS.n13790 VSS.n13619 0.457643
R18716 VSS.n14508 VSS.n14136 0.457643
R18717 VSS.n14494 VSS.n14493 0.457643
R18718 VSS.n14638 VSS.n14637 0.457643
R18719 VSS.n14382 VSS.n14211 0.457643
R18720 VSS.n15100 VSS.n14728 0.457643
R18721 VSS.n15086 VSS.n15085 0.457643
R18722 VSS.n15230 VSS.n15229 0.457643
R18723 VSS.n14974 VSS.n14803 0.457643
R18724 VSS.n15692 VSS.n15320 0.457643
R18725 VSS.n15678 VSS.n15677 0.457643
R18726 VSS.n15822 VSS.n15821 0.457643
R18727 VSS.n15566 VSS.n15395 0.457643
R18728 VSS.n15925 VSS.n6715 0.457643
R18729 VSS.n15911 VSS.n6813 0.457643
R18730 VSS.n15844 VSS.n6910 0.457643
R18731 VSS.n6674 VSS.n6503 0.457643
R18732 VSS.n7404 VSS.n7031 0.457643
R18733 VSS.n7390 VSS.n7389 0.457643
R18734 VSS.n7534 VSS.n7533 0.457643
R18735 VSS.n7278 VSS.n7106 0.457643
R18736 VSS.n18716 VSS.n129 0.457643
R18737 VSS.n18702 VSS.n18701 0.457643
R18738 VSS.n18846 VSS.n18845 0.457643
R18739 VSS.n18590 VSS.n197 0.457643
R18740 VSS.n839 VSS.n535 0.457643
R18741 VSS.n825 VSS.n636 0.457643
R18742 VSS.n18868 VSS.n18867 0.457643
R18743 VSS.n976 VSS.n882 0.457643
R18744 VSS.n17939 VSS.n1295 0.457643
R18745 VSS.n17872 VSS.n1392 0.457643
R18746 VSS.n18861 VSS 0.415989
R18747 VSS.n15837 VSS 0.415941
R18748 VSS.n14060 VSS 0.415941
R18749 VSS.n11692 VSS 0.415941
R18750 VSS.n9324 VSS 0.415941
R18751 VSS.n18889 VSS 0.415941
R18752 VSS.n3999 VSS 0.415941
R18753 VSS VSS.n16859 0.415941
R18754 VSS.n14652 VSS 0.382853
R18755 VSS.n4591 VSS 0.382853
R18756 VSS.n1243 VSS.n1234 0.366214
R18757 VSS.n1274 VSS.n1273 0.366214
R18758 VSS.n1108 VSS.n1101 0.366214
R18759 VSS.n1140 VSS.n1139 0.366214
R18760 VSS.n17026 VSS.n16987 0.366214
R18761 VSS.n17086 VSS.n17084 0.366214
R18762 VSS.n17522 VSS.n17520 0.366214
R18763 VSS.n17588 VSS.n17428 0.366214
R18764 VSS.n17618 VSS.n17401 0.366214
R18765 VSS.n17678 VSS.n17676 0.366214
R18766 VSS.n18260 VSS.n18251 0.366214
R18767 VSS.n18291 VSS.n18290 0.366214
R18768 VSS.n18099 VSS.n18097 0.366214
R18769 VSS.n18165 VSS.n220 0.366214
R18770 VSS.n9668 VSS.n9451 0.366214
R18771 VSS.n9728 VSS.n9726 0.366214
R18772 VSS.n9572 VSS.n9570 0.366214
R18773 VSS.n9638 VSS.n9478 0.366214
R18774 VSS.n16611 VSS.n16393 0.366214
R18775 VSS.n16671 VSS.n16669 0.366214
R18776 VSS.n16506 VSS.n16468 0.366214
R18777 VSS.n16567 VSS.n16565 0.366214
R18778 VSS.n16018 VSS.n1565 0.366214
R18779 VSS.n16078 VSS.n16076 0.366214
R18780 VSS.n1671 VSS.n1633 0.366214
R18781 VSS.n1732 VSS.n1730 0.366214
R18782 VSS.n2025 VSS.n2016 0.366214
R18783 VSS.n2056 VSS.n2055 0.366214
R18784 VSS.n1864 VSS.n1862 0.366214
R18785 VSS.n1930 VSS.n1770 0.366214
R18786 VSS.n3159 VSS.n2942 0.366214
R18787 VSS.n3219 VSS.n3217 0.366214
R18788 VSS.n3063 VSS.n3061 0.366214
R18789 VSS.n3129 VSS.n2969 0.366214
R18790 VSS.n3751 VSS.n3534 0.366214
R18791 VSS.n3811 VSS.n3809 0.366214
R18792 VSS.n3655 VSS.n3653 0.366214
R18793 VSS.n3721 VSS.n3561 0.366214
R18794 VSS.n4343 VSS.n4126 0.366214
R18795 VSS.n4403 VSS.n4401 0.366214
R18796 VSS.n4247 VSS.n4245 0.366214
R18797 VSS.n4313 VSS.n4153 0.366214
R18798 VSS.n4935 VSS.n4718 0.366214
R18799 VSS.n4995 VSS.n4993 0.366214
R18800 VSS.n4839 VSS.n4837 0.366214
R18801 VSS.n4905 VSS.n4745 0.366214
R18802 VSS.n2621 VSS.n2612 0.366214
R18803 VSS.n2652 VSS.n2651 0.366214
R18804 VSS.n2460 VSS.n2458 0.366214
R18805 VSS.n2526 VSS.n2366 0.366214
R18806 VSS.n5582 VSS.n5573 0.366214
R18807 VSS.n5613 VSS.n5612 0.366214
R18808 VSS.n5421 VSS.n5419 0.366214
R18809 VSS.n5487 VSS.n5327 0.366214
R18810 VSS.n6155 VSS.n6146 0.366214
R18811 VSS.n6186 VSS.n6185 0.366214
R18812 VSS.n5994 VSS.n5992 0.366214
R18813 VSS.n6060 VSS.n5900 0.366214
R18814 VSS.n7892 VSS.n7675 0.366214
R18815 VSS.n7952 VSS.n7950 0.366214
R18816 VSS.n7796 VSS.n7794 0.366214
R18817 VSS.n7862 VSS.n7702 0.366214
R18818 VSS.n8484 VSS.n8267 0.366214
R18819 VSS.n8544 VSS.n8542 0.366214
R18820 VSS.n8388 VSS.n8386 0.366214
R18821 VSS.n8454 VSS.n8294 0.366214
R18822 VSS.n9076 VSS.n8859 0.366214
R18823 VSS.n9136 VSS.n9134 0.366214
R18824 VSS.n8980 VSS.n8978 0.366214
R18825 VSS.n9046 VSS.n8886 0.366214
R18826 VSS.n10260 VSS.n10043 0.366214
R18827 VSS.n10320 VSS.n10318 0.366214
R18828 VSS.n10164 VSS.n10162 0.366214
R18829 VSS.n10230 VSS.n10070 0.366214
R18830 VSS.n10852 VSS.n10635 0.366214
R18831 VSS.n10912 VSS.n10910 0.366214
R18832 VSS.n10756 VSS.n10754 0.366214
R18833 VSS.n10822 VSS.n10662 0.366214
R18834 VSS.n11444 VSS.n11227 0.366214
R18835 VSS.n11504 VSS.n11502 0.366214
R18836 VSS.n11348 VSS.n11346 0.366214
R18837 VSS.n11414 VSS.n11254 0.366214
R18838 VSS.n12036 VSS.n11819 0.366214
R18839 VSS.n12096 VSS.n12094 0.366214
R18840 VSS.n11940 VSS.n11938 0.366214
R18841 VSS.n12006 VSS.n11846 0.366214
R18842 VSS.n12628 VSS.n12411 0.366214
R18843 VSS.n12688 VSS.n12686 0.366214
R18844 VSS.n12532 VSS.n12530 0.366214
R18845 VSS.n12598 VSS.n12438 0.366214
R18846 VSS.n13220 VSS.n13003 0.366214
R18847 VSS.n13280 VSS.n13278 0.366214
R18848 VSS.n13124 VSS.n13122 0.366214
R18849 VSS.n13190 VSS.n13030 0.366214
R18850 VSS.n13812 VSS.n13595 0.366214
R18851 VSS.n13872 VSS.n13870 0.366214
R18852 VSS.n13716 VSS.n13714 0.366214
R18853 VSS.n13782 VSS.n13622 0.366214
R18854 VSS.n14404 VSS.n14187 0.366214
R18855 VSS.n14464 VSS.n14462 0.366214
R18856 VSS.n14308 VSS.n14306 0.366214
R18857 VSS.n14374 VSS.n14214 0.366214
R18858 VSS.n14996 VSS.n14779 0.366214
R18859 VSS.n15056 VSS.n15054 0.366214
R18860 VSS.n14900 VSS.n14898 0.366214
R18861 VSS.n14966 VSS.n14806 0.366214
R18862 VSS.n15588 VSS.n15371 0.366214
R18863 VSS.n15648 VSS.n15646 0.366214
R18864 VSS.n15492 VSS.n15490 0.366214
R18865 VSS.n15558 VSS.n15398 0.366214
R18866 VSS.n6761 VSS.n6752 0.366214
R18867 VSS.n6792 VSS.n6791 0.366214
R18868 VSS.n6600 VSS.n6598 0.366214
R18869 VSS.n6666 VSS.n6506 0.366214
R18870 VSS.n7300 VSS.n7082 0.366214
R18871 VSS.n7360 VSS.n7358 0.366214
R18872 VSS.n7195 VSS.n7157 0.366214
R18873 VSS.n7256 VSS.n7254 0.366214
R18874 VSS.n18612 VSS.n180 0.366214
R18875 VSS.n18672 VSS.n18670 0.366214
R18876 VSS.n363 VSS.n343 0.366214
R18877 VSS.n397 VSS.n396 0.366214
R18878 VSS.n584 VSS.n575 0.366214
R18879 VSS.n615 VSS.n614 0.366214
R18880 VSS.n927 VSS.n920 0.366214
R18881 VSS.n959 VSS.n958 0.366214
R18882 VSS.n1025 VSS 0.301636
R18883 VSS.n17502 VSS 0.301636
R18884 VSS.n18079 VSS 0.301636
R18885 VSS.n16488 VSS 0.301636
R18886 VSS.n1653 VSS 0.301636
R18887 VSS.n1844 VSS 0.301636
R18888 VSS.n3043 VSS 0.301636
R18889 VSS.n3635 VSS 0.301636
R18890 VSS.n4227 VSS 0.301636
R18891 VSS.n4819 VSS 0.301636
R18892 VSS.n2440 VSS 0.301636
R18893 VSS.n5401 VSS 0.301636
R18894 VSS.n5974 VSS 0.301636
R18895 VSS.n7776 VSS 0.301636
R18896 VSS.n8368 VSS 0.301636
R18897 VSS.n8960 VSS 0.301636
R18898 VSS.n10144 VSS 0.301636
R18899 VSS.n10736 VSS 0.301636
R18900 VSS.n11328 VSS 0.301636
R18901 VSS.n11920 VSS 0.301636
R18902 VSS.n12512 VSS 0.301636
R18903 VSS.n13104 VSS 0.301636
R18904 VSS.n13696 VSS 0.301636
R18905 VSS.n14288 VSS 0.301636
R18906 VSS.n14880 VSS 0.301636
R18907 VSS.n15472 VSS 0.301636
R18908 VSS.n6580 VSS 0.301636
R18909 VSS.n7177 VSS 0.301636
R18910 VSS.n292 VSS 0.301636
R18911 VSS.n458 VSS 0.301636
R18912 VSS.n1160 VSS 0.301636
R18913 VSS VSS.n17271 0.300964
R18914 VSS VSS.n17863 0.300964
R18915 VSS.n18430 VSS 0.300964
R18916 VSS VSS.n9914 0.300964
R18917 VSS VSS.n16857 0.300964
R18918 VSS VSS.n16264 0.300964
R18919 VSS.n2221 VSS 0.300964
R18920 VSS VSS.n3405 0.300964
R18921 VSS VSS.n3997 0.300964
R18922 VSS VSS.n4589 0.300964
R18923 VSS VSS.n5181 0.300964
R18924 VSS.n5186 VSS 0.300964
R18925 VSS VSS.n18887 0.300964
R18926 VSS.n6351 VSS 0.300964
R18927 VSS VSS.n8138 0.300964
R18928 VSS VSS.n8730 0.300964
R18929 VSS VSS.n9322 0.300964
R18930 VSS VSS.n10506 0.300964
R18931 VSS VSS.n11098 0.300964
R18932 VSS VSS.n11690 0.300964
R18933 VSS VSS.n12282 0.300964
R18934 VSS VSS.n12874 0.300964
R18935 VSS VSS.n13466 0.300964
R18936 VSS VSS.n14058 0.300964
R18937 VSS VSS.n14650 0.300964
R18938 VSS VSS.n15242 0.300964
R18939 VSS VSS.n15834 0.300964
R18940 VSS.n15839 VSS 0.300964
R18941 VSS VSS.n7546 0.300964
R18942 VSS VSS.n18858 0.300964
R18943 VSS.n18862 VSS 0.300964
R18944 VSS.n17867 VSS 0.300964
R18945 VSS.n9552 VSS 0.2995
R18946 VSS.n17008 VSS 0.29425
R18947 VSS.n17600 VSS 0.29425
R18948 VSS.n18177 VSS 0.29425
R18949 VSS.n9650 VSS 0.29425
R18950 VSS.n16593 VSS 0.29425
R18951 VSS.n16000 VSS 0.29425
R18952 VSS.n1942 VSS 0.29425
R18953 VSS.n3141 VSS 0.29425
R18954 VSS.n3733 VSS 0.29425
R18955 VSS.n4325 VSS 0.29425
R18956 VSS.n4917 VSS 0.29425
R18957 VSS.n2538 VSS 0.29425
R18958 VSS.n5499 VSS 0.29425
R18959 VSS.n6072 VSS 0.29425
R18960 VSS.n7874 VSS 0.29425
R18961 VSS.n8466 VSS 0.29425
R18962 VSS.n9058 VSS 0.29425
R18963 VSS.n10242 VSS 0.29425
R18964 VSS.n10834 VSS 0.29425
R18965 VSS.n11426 VSS 0.29425
R18966 VSS.n12018 VSS 0.29425
R18967 VSS.n12610 VSS 0.29425
R18968 VSS.n13202 VSS 0.29425
R18969 VSS.n13794 VSS 0.29425
R18970 VSS.n14386 VSS 0.29425
R18971 VSS.n14978 VSS 0.29425
R18972 VSS.n15570 VSS 0.29425
R18973 VSS.n6678 VSS 0.29425
R18974 VSS.n7282 VSS 0.29425
R18975 VSS.n18594 VSS 0.29425
R18976 VSS VSS.n879 0.29425
R18977 VSS.n17162 VSS.n16917 0.274786
R18978 VSS.n17185 VSS.n17184 0.274786
R18979 VSS.n17199 VSS.n16896 0.274786
R18980 VSS.n17239 VSS.n16879 0.274786
R18981 VSS.n17754 VSS.n17331 0.274786
R18982 VSS.n17777 VSS.n17776 0.274786
R18983 VSS.n17791 VSS.n17310 0.274786
R18984 VSS.n17831 VSS.n17293 0.274786
R18985 VSS.n18367 VSS.n18366 0.274786
R18986 VSS.n18375 VSS.n18357 0.274786
R18987 VSS.n18404 VSS.n18396 0.274786
R18988 VSS.n18442 VSS.n18420 0.274786
R18989 VSS.n9804 VSS.n9381 0.274786
R18990 VSS.n9827 VSS.n9826 0.274786
R18991 VSS.n9841 VSS.n9360 0.274786
R18992 VSS.n9881 VSS.n9343 0.274786
R18993 VSS.n16747 VSS.n16323 0.274786
R18994 VSS.n16770 VSS.n16769 0.274786
R18995 VSS.n16784 VSS.n16302 0.274786
R18996 VSS.n16824 VSS.n16285 0.274786
R18997 VSS.n16154 VSS.n1495 0.274786
R18998 VSS.n16177 VSS.n16176 0.274786
R18999 VSS.n16191 VSS.n1474 0.274786
R19000 VSS.n16231 VSS.n1457 0.274786
R19001 VSS.n2283 VSS.n2103 0.274786
R19002 VSS.n2145 VSS.n2144 0.274786
R19003 VSS.n2179 VSS.n2126 0.274786
R19004 VSS.n2194 VSS.n2193 0.274786
R19005 VSS.n3295 VSS.n2872 0.274786
R19006 VSS.n3318 VSS.n3317 0.274786
R19007 VSS.n3332 VSS.n2851 0.274786
R19008 VSS.n3372 VSS.n2834 0.274786
R19009 VSS.n3887 VSS.n3464 0.274786
R19010 VSS.n3910 VSS.n3909 0.274786
R19011 VSS.n3924 VSS.n3443 0.274786
R19012 VSS.n3964 VSS.n3426 0.274786
R19013 VSS.n4479 VSS.n4056 0.274786
R19014 VSS.n4502 VSS.n4501 0.274786
R19015 VSS.n4516 VSS.n4035 0.274786
R19016 VSS.n4556 VSS.n4018 0.274786
R19017 VSS.n5071 VSS.n4648 0.274786
R19018 VSS.n5094 VSS.n5093 0.274786
R19019 VSS.n5108 VSS.n4627 0.274786
R19020 VSS.n5148 VSS.n4610 0.274786
R19021 VSS.n5248 VSS.n2699 0.274786
R19022 VSS.n2741 VSS.n2740 0.274786
R19023 VSS.n2775 VSS.n2722 0.274786
R19024 VSS.n2790 VSS.n2789 0.274786
R19025 VSS.n5821 VSS.n5660 0.274786
R19026 VSS.n5702 VSS.n5701 0.274786
R19027 VSS.n5749 VSS.n5683 0.274786
R19028 VSS.n5764 VSS.n5763 0.274786
R19029 VSS.n6413 VSS.n6233 0.274786
R19030 VSS.n6275 VSS.n6274 0.274786
R19031 VSS.n6309 VSS.n6256 0.274786
R19032 VSS.n6324 VSS.n6323 0.274786
R19033 VSS.n8028 VSS.n7605 0.274786
R19034 VSS.n8051 VSS.n8050 0.274786
R19035 VSS.n8065 VSS.n7584 0.274786
R19036 VSS.n8105 VSS.n7567 0.274786
R19037 VSS.n8620 VSS.n8197 0.274786
R19038 VSS.n8643 VSS.n8642 0.274786
R19039 VSS.n8657 VSS.n8176 0.274786
R19040 VSS.n8697 VSS.n8159 0.274786
R19041 VSS.n9212 VSS.n8789 0.274786
R19042 VSS.n9235 VSS.n9234 0.274786
R19043 VSS.n9249 VSS.n8768 0.274786
R19044 VSS.n9289 VSS.n8751 0.274786
R19045 VSS.n10396 VSS.n9973 0.274786
R19046 VSS.n10419 VSS.n10418 0.274786
R19047 VSS.n10433 VSS.n9952 0.274786
R19048 VSS.n10473 VSS.n9935 0.274786
R19049 VSS.n10988 VSS.n10565 0.274786
R19050 VSS.n11011 VSS.n11010 0.274786
R19051 VSS.n11025 VSS.n10544 0.274786
R19052 VSS.n11065 VSS.n10527 0.274786
R19053 VSS.n11580 VSS.n11157 0.274786
R19054 VSS.n11603 VSS.n11602 0.274786
R19055 VSS.n11617 VSS.n11136 0.274786
R19056 VSS.n11657 VSS.n11119 0.274786
R19057 VSS.n12172 VSS.n11749 0.274786
R19058 VSS.n12195 VSS.n12194 0.274786
R19059 VSS.n12209 VSS.n11728 0.274786
R19060 VSS.n12249 VSS.n11711 0.274786
R19061 VSS.n12764 VSS.n12341 0.274786
R19062 VSS.n12787 VSS.n12786 0.274786
R19063 VSS.n12801 VSS.n12320 0.274786
R19064 VSS.n12841 VSS.n12303 0.274786
R19065 VSS.n13356 VSS.n12933 0.274786
R19066 VSS.n13379 VSS.n13378 0.274786
R19067 VSS.n13393 VSS.n12912 0.274786
R19068 VSS.n13433 VSS.n12895 0.274786
R19069 VSS.n13948 VSS.n13525 0.274786
R19070 VSS.n13971 VSS.n13970 0.274786
R19071 VSS.n13985 VSS.n13504 0.274786
R19072 VSS.n14025 VSS.n13487 0.274786
R19073 VSS.n14540 VSS.n14117 0.274786
R19074 VSS.n14563 VSS.n14562 0.274786
R19075 VSS.n14577 VSS.n14096 0.274786
R19076 VSS.n14617 VSS.n14079 0.274786
R19077 VSS.n15132 VSS.n14709 0.274786
R19078 VSS.n15155 VSS.n15154 0.274786
R19079 VSS.n15169 VSS.n14688 0.274786
R19080 VSS.n15209 VSS.n14671 0.274786
R19081 VSS.n15724 VSS.n15301 0.274786
R19082 VSS.n15747 VSS.n15746 0.274786
R19083 VSS.n15761 VSS.n15280 0.274786
R19084 VSS.n15801 VSS.n15263 0.274786
R19085 VSS.n15901 VSS.n6839 0.274786
R19086 VSS.n6881 VSS.n6880 0.274786
R19087 VSS.n6915 VSS.n6862 0.274786
R19088 VSS.n6930 VSS.n6929 0.274786
R19089 VSS.n7436 VSS.n7012 0.274786
R19090 VSS.n7459 VSS.n7458 0.274786
R19091 VSS.n7473 VSS.n6991 0.274786
R19092 VSS.n7513 VSS.n6974 0.274786
R19093 VSS.n18748 VSS.n110 0.274786
R19094 VSS.n18771 VSS.n18770 0.274786
R19095 VSS.n18785 VSS.n89 0.274786
R19096 VSS.n18825 VSS.n72 0.274786
R19097 VSS.n815 VSS.n662 0.274786
R19098 VSS.n704 VSS.n703 0.274786
R19099 VSS.n747 VSS.n685 0.274786
R19100 VSS.n762 VSS.n743 0.274786
R19101 VSS.n17929 VSS.n1321 0.274786
R19102 VSS.n1363 VSS.n1362 0.274786
R19103 VSS.n1397 VSS.n1344 0.274786
R19104 VSS.n1412 VSS.n1411 0.274786
R19105 VSS VSS.n17007 0.206964
R19106 VSS VSS.n17599 0.206964
R19107 VSS VSS.n18176 0.206964
R19108 VSS VSS.n16592 0.206964
R19109 VSS VSS.n15999 0.206964
R19110 VSS VSS.n1941 0.206964
R19111 VSS VSS.n3140 0.206964
R19112 VSS VSS.n3732 0.206964
R19113 VSS VSS.n4324 0.206964
R19114 VSS VSS.n4916 0.206964
R19115 VSS VSS.n2537 0.206964
R19116 VSS VSS.n5498 0.206964
R19117 VSS VSS.n6071 0.206964
R19118 VSS VSS.n7873 0.206964
R19119 VSS VSS.n8465 0.206964
R19120 VSS VSS.n9057 0.206964
R19121 VSS VSS.n10241 0.206964
R19122 VSS VSS.n10833 0.206964
R19123 VSS VSS.n11425 0.206964
R19124 VSS VSS.n12017 0.206964
R19125 VSS VSS.n12609 0.206964
R19126 VSS VSS.n13201 0.206964
R19127 VSS VSS.n13793 0.206964
R19128 VSS VSS.n14385 0.206964
R19129 VSS VSS.n14977 0.206964
R19130 VSS VSS.n15569 0.206964
R19131 VSS VSS.n6677 0.206964
R19132 VSS VSS.n7281 0.206964
R19133 VSS VSS.n18593 0.206964
R19134 VSS.n880 VSS 0.206964
R19135 VSS VSS.n9649 0.2055
R19136 VSS.n1249 VSS.n1214 0.183357
R19137 VSS.n1250 VSS.n1249 0.183357
R19138 VSS.n1268 VSS.n1258 0.183357
R19139 VSS.n1268 VSS.n1259 0.183357
R19140 VSS.n1114 VSS.n1081 0.183357
R19141 VSS.n1115 VSS.n1114 0.183357
R19142 VSS.n1133 VSS.n1123 0.183357
R19143 VSS.n1133 VSS.n1124 0.183357
R19144 VSS.n17047 VSS.n16976 0.183357
R19145 VSS.n17048 VSS.n17047 0.183357
R19146 VSS.n17079 VSS.n16955 0.183357
R19147 VSS.n17079 VSS.n16956 0.183357
R19148 VSS.n17532 VSS.n17531 0.183357
R19149 VSS.n17531 VSS.n17478 0.183357
R19150 VSS.n17564 VSS.n17448 0.183357
R19151 VSS.n17564 VSS.n17449 0.183357
R19152 VSS.n17639 VSS.n17390 0.183357
R19153 VSS.n17640 VSS.n17639 0.183357
R19154 VSS.n17671 VSS.n17369 0.183357
R19155 VSS.n17671 VSS.n17370 0.183357
R19156 VSS.n18266 VSS.n18231 0.183357
R19157 VSS.n18267 VSS.n18266 0.183357
R19158 VSS.n18285 VSS.n18275 0.183357
R19159 VSS.n18285 VSS.n18276 0.183357
R19160 VSS.n18109 VSS.n18108 0.183357
R19161 VSS.n18108 VSS.n270 0.183357
R19162 VSS.n18141 VSS.n240 0.183357
R19163 VSS.n18141 VSS.n241 0.183357
R19164 VSS.n9689 VSS.n9440 0.183357
R19165 VSS.n9690 VSS.n9689 0.183357
R19166 VSS.n9721 VSS.n9419 0.183357
R19167 VSS.n9721 VSS.n9420 0.183357
R19168 VSS.n9582 VSS.n9581 0.183357
R19169 VSS.n9581 VSS.n9528 0.183357
R19170 VSS.n9614 VSS.n9498 0.183357
R19171 VSS.n9614 VSS.n9499 0.183357
R19172 VSS.n16632 VSS.n16382 0.183357
R19173 VSS.n16633 VSS.n16632 0.183357
R19174 VSS.n16664 VSS.n16361 0.183357
R19175 VSS.n16664 VSS.n16362 0.183357
R19176 VSS.n16527 VSS.n16459 0.183357
R19177 VSS.n16528 VSS.n16527 0.183357
R19178 VSS.n16559 VSS.n16436 0.183357
R19179 VSS.n16559 VSS.n16437 0.183357
R19180 VSS.n16039 VSS.n1554 0.183357
R19181 VSS.n16040 VSS.n16039 0.183357
R19182 VSS.n16071 VSS.n1533 0.183357
R19183 VSS.n16071 VSS.n1534 0.183357
R19184 VSS.n1692 VSS.n1624 0.183357
R19185 VSS.n1693 VSS.n1692 0.183357
R19186 VSS.n1724 VSS.n1601 0.183357
R19187 VSS.n1724 VSS.n1602 0.183357
R19188 VSS.n2031 VSS.n1996 0.183357
R19189 VSS.n2032 VSS.n2031 0.183357
R19190 VSS.n2050 VSS.n2040 0.183357
R19191 VSS.n2050 VSS.n2041 0.183357
R19192 VSS.n1874 VSS.n1873 0.183357
R19193 VSS.n1873 VSS.n1820 0.183357
R19194 VSS.n1906 VSS.n1790 0.183357
R19195 VSS.n1906 VSS.n1791 0.183357
R19196 VSS.n3180 VSS.n2931 0.183357
R19197 VSS.n3181 VSS.n3180 0.183357
R19198 VSS.n3212 VSS.n2910 0.183357
R19199 VSS.n3212 VSS.n2911 0.183357
R19200 VSS.n3073 VSS.n3072 0.183357
R19201 VSS.n3072 VSS.n3019 0.183357
R19202 VSS.n3105 VSS.n2989 0.183357
R19203 VSS.n3105 VSS.n2990 0.183357
R19204 VSS.n3772 VSS.n3523 0.183357
R19205 VSS.n3773 VSS.n3772 0.183357
R19206 VSS.n3804 VSS.n3502 0.183357
R19207 VSS.n3804 VSS.n3503 0.183357
R19208 VSS.n3665 VSS.n3664 0.183357
R19209 VSS.n3664 VSS.n3611 0.183357
R19210 VSS.n3697 VSS.n3581 0.183357
R19211 VSS.n3697 VSS.n3582 0.183357
R19212 VSS.n4364 VSS.n4115 0.183357
R19213 VSS.n4365 VSS.n4364 0.183357
R19214 VSS.n4396 VSS.n4094 0.183357
R19215 VSS.n4396 VSS.n4095 0.183357
R19216 VSS.n4257 VSS.n4256 0.183357
R19217 VSS.n4256 VSS.n4203 0.183357
R19218 VSS.n4289 VSS.n4173 0.183357
R19219 VSS.n4289 VSS.n4174 0.183357
R19220 VSS.n4956 VSS.n4707 0.183357
R19221 VSS.n4957 VSS.n4956 0.183357
R19222 VSS.n4988 VSS.n4686 0.183357
R19223 VSS.n4988 VSS.n4687 0.183357
R19224 VSS.n4849 VSS.n4848 0.183357
R19225 VSS.n4848 VSS.n4795 0.183357
R19226 VSS.n4881 VSS.n4765 0.183357
R19227 VSS.n4881 VSS.n4766 0.183357
R19228 VSS.n2627 VSS.n2592 0.183357
R19229 VSS.n2628 VSS.n2627 0.183357
R19230 VSS.n2646 VSS.n2636 0.183357
R19231 VSS.n2646 VSS.n2637 0.183357
R19232 VSS.n2470 VSS.n2469 0.183357
R19233 VSS.n2469 VSS.n2416 0.183357
R19234 VSS.n2502 VSS.n2386 0.183357
R19235 VSS.n2502 VSS.n2387 0.183357
R19236 VSS.n5588 VSS.n5553 0.183357
R19237 VSS.n5589 VSS.n5588 0.183357
R19238 VSS.n5607 VSS.n5597 0.183357
R19239 VSS.n5607 VSS.n5598 0.183357
R19240 VSS.n5431 VSS.n5430 0.183357
R19241 VSS.n5430 VSS.n5377 0.183357
R19242 VSS.n5463 VSS.n5347 0.183357
R19243 VSS.n5463 VSS.n5348 0.183357
R19244 VSS.n6161 VSS.n6126 0.183357
R19245 VSS.n6162 VSS.n6161 0.183357
R19246 VSS.n6180 VSS.n6170 0.183357
R19247 VSS.n6180 VSS.n6171 0.183357
R19248 VSS.n6004 VSS.n6003 0.183357
R19249 VSS.n6003 VSS.n5950 0.183357
R19250 VSS.n6036 VSS.n5920 0.183357
R19251 VSS.n6036 VSS.n5921 0.183357
R19252 VSS.n7913 VSS.n7664 0.183357
R19253 VSS.n7914 VSS.n7913 0.183357
R19254 VSS.n7945 VSS.n7643 0.183357
R19255 VSS.n7945 VSS.n7644 0.183357
R19256 VSS.n7806 VSS.n7805 0.183357
R19257 VSS.n7805 VSS.n7752 0.183357
R19258 VSS.n7838 VSS.n7722 0.183357
R19259 VSS.n7838 VSS.n7723 0.183357
R19260 VSS.n8505 VSS.n8256 0.183357
R19261 VSS.n8506 VSS.n8505 0.183357
R19262 VSS.n8537 VSS.n8235 0.183357
R19263 VSS.n8537 VSS.n8236 0.183357
R19264 VSS.n8398 VSS.n8397 0.183357
R19265 VSS.n8397 VSS.n8344 0.183357
R19266 VSS.n8430 VSS.n8314 0.183357
R19267 VSS.n8430 VSS.n8315 0.183357
R19268 VSS.n9097 VSS.n8848 0.183357
R19269 VSS.n9098 VSS.n9097 0.183357
R19270 VSS.n9129 VSS.n8827 0.183357
R19271 VSS.n9129 VSS.n8828 0.183357
R19272 VSS.n8990 VSS.n8989 0.183357
R19273 VSS.n8989 VSS.n8936 0.183357
R19274 VSS.n9022 VSS.n8906 0.183357
R19275 VSS.n9022 VSS.n8907 0.183357
R19276 VSS.n10281 VSS.n10032 0.183357
R19277 VSS.n10282 VSS.n10281 0.183357
R19278 VSS.n10313 VSS.n10011 0.183357
R19279 VSS.n10313 VSS.n10012 0.183357
R19280 VSS.n10174 VSS.n10173 0.183357
R19281 VSS.n10173 VSS.n10120 0.183357
R19282 VSS.n10206 VSS.n10090 0.183357
R19283 VSS.n10206 VSS.n10091 0.183357
R19284 VSS.n10873 VSS.n10624 0.183357
R19285 VSS.n10874 VSS.n10873 0.183357
R19286 VSS.n10905 VSS.n10603 0.183357
R19287 VSS.n10905 VSS.n10604 0.183357
R19288 VSS.n10766 VSS.n10765 0.183357
R19289 VSS.n10765 VSS.n10712 0.183357
R19290 VSS.n10798 VSS.n10682 0.183357
R19291 VSS.n10798 VSS.n10683 0.183357
R19292 VSS.n11465 VSS.n11216 0.183357
R19293 VSS.n11466 VSS.n11465 0.183357
R19294 VSS.n11497 VSS.n11195 0.183357
R19295 VSS.n11497 VSS.n11196 0.183357
R19296 VSS.n11358 VSS.n11357 0.183357
R19297 VSS.n11357 VSS.n11304 0.183357
R19298 VSS.n11390 VSS.n11274 0.183357
R19299 VSS.n11390 VSS.n11275 0.183357
R19300 VSS.n12057 VSS.n11808 0.183357
R19301 VSS.n12058 VSS.n12057 0.183357
R19302 VSS.n12089 VSS.n11787 0.183357
R19303 VSS.n12089 VSS.n11788 0.183357
R19304 VSS.n11950 VSS.n11949 0.183357
R19305 VSS.n11949 VSS.n11896 0.183357
R19306 VSS.n11982 VSS.n11866 0.183357
R19307 VSS.n11982 VSS.n11867 0.183357
R19308 VSS.n12649 VSS.n12400 0.183357
R19309 VSS.n12650 VSS.n12649 0.183357
R19310 VSS.n12681 VSS.n12379 0.183357
R19311 VSS.n12681 VSS.n12380 0.183357
R19312 VSS.n12542 VSS.n12541 0.183357
R19313 VSS.n12541 VSS.n12488 0.183357
R19314 VSS.n12574 VSS.n12458 0.183357
R19315 VSS.n12574 VSS.n12459 0.183357
R19316 VSS.n13241 VSS.n12992 0.183357
R19317 VSS.n13242 VSS.n13241 0.183357
R19318 VSS.n13273 VSS.n12971 0.183357
R19319 VSS.n13273 VSS.n12972 0.183357
R19320 VSS.n13134 VSS.n13133 0.183357
R19321 VSS.n13133 VSS.n13080 0.183357
R19322 VSS.n13166 VSS.n13050 0.183357
R19323 VSS.n13166 VSS.n13051 0.183357
R19324 VSS.n13833 VSS.n13584 0.183357
R19325 VSS.n13834 VSS.n13833 0.183357
R19326 VSS.n13865 VSS.n13563 0.183357
R19327 VSS.n13865 VSS.n13564 0.183357
R19328 VSS.n13726 VSS.n13725 0.183357
R19329 VSS.n13725 VSS.n13672 0.183357
R19330 VSS.n13758 VSS.n13642 0.183357
R19331 VSS.n13758 VSS.n13643 0.183357
R19332 VSS.n14425 VSS.n14176 0.183357
R19333 VSS.n14426 VSS.n14425 0.183357
R19334 VSS.n14457 VSS.n14155 0.183357
R19335 VSS.n14457 VSS.n14156 0.183357
R19336 VSS.n14318 VSS.n14317 0.183357
R19337 VSS.n14317 VSS.n14264 0.183357
R19338 VSS.n14350 VSS.n14234 0.183357
R19339 VSS.n14350 VSS.n14235 0.183357
R19340 VSS.n15017 VSS.n14768 0.183357
R19341 VSS.n15018 VSS.n15017 0.183357
R19342 VSS.n15049 VSS.n14747 0.183357
R19343 VSS.n15049 VSS.n14748 0.183357
R19344 VSS.n14910 VSS.n14909 0.183357
R19345 VSS.n14909 VSS.n14856 0.183357
R19346 VSS.n14942 VSS.n14826 0.183357
R19347 VSS.n14942 VSS.n14827 0.183357
R19348 VSS.n15609 VSS.n15360 0.183357
R19349 VSS.n15610 VSS.n15609 0.183357
R19350 VSS.n15641 VSS.n15339 0.183357
R19351 VSS.n15641 VSS.n15340 0.183357
R19352 VSS.n15502 VSS.n15501 0.183357
R19353 VSS.n15501 VSS.n15448 0.183357
R19354 VSS.n15534 VSS.n15418 0.183357
R19355 VSS.n15534 VSS.n15419 0.183357
R19356 VSS.n6767 VSS.n6732 0.183357
R19357 VSS.n6768 VSS.n6767 0.183357
R19358 VSS.n6786 VSS.n6776 0.183357
R19359 VSS.n6786 VSS.n6777 0.183357
R19360 VSS.n6610 VSS.n6609 0.183357
R19361 VSS.n6609 VSS.n6556 0.183357
R19362 VSS.n6642 VSS.n6526 0.183357
R19363 VSS.n6642 VSS.n6527 0.183357
R19364 VSS.n7321 VSS.n7071 0.183357
R19365 VSS.n7322 VSS.n7321 0.183357
R19366 VSS.n7353 VSS.n7050 0.183357
R19367 VSS.n7353 VSS.n7051 0.183357
R19368 VSS.n7216 VSS.n7148 0.183357
R19369 VSS.n7217 VSS.n7216 0.183357
R19370 VSS.n7248 VSS.n7125 0.183357
R19371 VSS.n7248 VSS.n7126 0.183357
R19372 VSS.n18633 VSS.n169 0.183357
R19373 VSS.n18634 VSS.n18633 0.183357
R19374 VSS.n18665 VSS.n148 0.183357
R19375 VSS.n18665 VSS.n149 0.183357
R19376 VSS.n371 VSS.n342 0.183357
R19377 VSS.n371 VSS.n338 0.183357
R19378 VSS.n386 VSS.n334 0.183357
R19379 VSS.n386 VSS.n332 0.183357
R19380 VSS.n590 VSS.n552 0.183357
R19381 VSS.n591 VSS.n590 0.183357
R19382 VSS.n609 VSS.n599 0.183357
R19383 VSS.n609 VSS.n600 0.183357
R19384 VSS.n933 VSS.n900 0.183357
R19385 VSS.n934 VSS.n933 0.183357
R19386 VSS.n952 VSS.n942 0.183357
R19387 VSS.n952 VSS.n943 0.183357
R19388 VSS.n17272 VSS 0.107929
R19389 VSS.n17864 VSS 0.107929
R19390 VSS VSS.n18429 0.107929
R19391 VSS.n9915 VSS 0.107929
R19392 VSS.n16858 VSS 0.107929
R19393 VSS.n16265 VSS 0.107929
R19394 VSS VSS.n2220 0.107929
R19395 VSS.n3406 VSS 0.107929
R19396 VSS.n3998 VSS 0.107929
R19397 VSS.n4590 VSS 0.107929
R19398 VSS.n5182 VSS 0.107929
R19399 VSS VSS.n5185 0.107929
R19400 VSS.n18888 VSS 0.107929
R19401 VSS VSS.n6350 0.107929
R19402 VSS.n8139 VSS 0.107929
R19403 VSS.n8731 VSS 0.107929
R19404 VSS.n9323 VSS 0.107929
R19405 VSS.n10507 VSS 0.107929
R19406 VSS.n11099 VSS 0.107929
R19407 VSS.n11691 VSS 0.107929
R19408 VSS.n12283 VSS 0.107929
R19409 VSS.n12875 VSS 0.107929
R19410 VSS.n13467 VSS 0.107929
R19411 VSS.n14059 VSS 0.107929
R19412 VSS.n14651 VSS 0.107929
R19413 VSS.n15243 VSS 0.107929
R19414 VSS.n15835 VSS 0.107929
R19415 VSS VSS.n15838 0.107929
R19416 VSS.n7547 VSS 0.107929
R19417 VSS.n18859 VSS 0.107929
R19418 VSS VSS.n18861 0.107929
R19419 VSS VSS.n17866 0.107929
R19420 VSS VSS.n17133 0.107593
R19421 VSS VSS.n17725 0.107593
R19422 VSS VSS.n18327 0.107593
R19423 VSS VSS.n9775 0.107593
R19424 VSS VSS.n16718 0.107593
R19425 VSS VSS.n16125 0.107593
R19426 VSS VSS.n2091 0.107593
R19427 VSS VSS.n3266 0.107593
R19428 VSS VSS.n3858 0.107593
R19429 VSS VSS.n4450 0.107593
R19430 VSS VSS.n5042 0.107593
R19431 VSS VSS.n2687 0.107593
R19432 VSS VSS.n5648 0.107593
R19433 VSS VSS.n6221 0.107593
R19434 VSS VSS.n7999 0.107593
R19435 VSS VSS.n8591 0.107593
R19436 VSS VSS.n9183 0.107593
R19437 VSS VSS.n10367 0.107593
R19438 VSS VSS.n10959 0.107593
R19439 VSS VSS.n11551 0.107593
R19440 VSS VSS.n12143 0.107593
R19441 VSS VSS.n12735 0.107593
R19442 VSS VSS.n13327 0.107593
R19443 VSS VSS.n13919 0.107593
R19444 VSS VSS.n14511 0.107593
R19445 VSS VSS.n15103 0.107593
R19446 VSS VSS.n15695 0.107593
R19447 VSS VSS.n6827 0.107593
R19448 VSS VSS.n7407 0.107593
R19449 VSS VSS.n18719 0.107593
R19450 VSS VSS.n650 0.107593
R19451 VSS VSS.n1309 0.107593
R19452 VSS.n1275 VSS.n1274 0.0919286
R19453 VSS.n1283 VSS.n1201 0.0919286
R19454 VSS.n17953 VSS.n17952 0.0919286
R19455 VSS.n1141 VSS.n1140 0.0919286
R19456 VSS.n1149 VSS.n1067 0.0919286
R19457 VSS.n18002 VSS.n18001 0.0919286
R19458 VSS.n17169 VSS.n16912 0.0919286
R19459 VSS.n17220 VSS.n17219 0.0919286
R19460 VSS.n17086 VSS.n17085 0.0919286
R19461 VSS.n17100 VSS.n16940 0.0919286
R19462 VSS.n17130 VSS.n17129 0.0919286
R19463 VSS.n17588 VSS.n17429 0.0919286
R19464 VSS.n17437 VSS.n17435 0.0919286
R19465 VSS.n17596 VSS.n17595 0.0919286
R19466 VSS.n17761 VSS.n17326 0.0919286
R19467 VSS.n17812 VSS.n17811 0.0919286
R19468 VSS.n17678 VSS.n17677 0.0919286
R19469 VSS.n17692 VSS.n17354 0.0919286
R19470 VSS.n17722 VSS.n17721 0.0919286
R19471 VSS.n18292 VSS.n18291 0.0919286
R19472 VSS.n18300 VSS.n18218 0.0919286
R19473 VSS.n18542 VSS.n18541 0.0919286
R19474 VSS.n18380 VSS.n18344 0.0919286
R19475 VSS.n18492 VSS.n18491 0.0919286
R19476 VSS.n18165 VSS.n221 0.0919286
R19477 VSS.n229 VSS.n227 0.0919286
R19478 VSS.n18173 VSS.n18172 0.0919286
R19479 VSS.n9728 VSS.n9727 0.0919286
R19480 VSS.n9742 VSS.n9404 0.0919286
R19481 VSS.n9772 VSS.n9771 0.0919286
R19482 VSS.n9811 VSS.n9376 0.0919286
R19483 VSS.n9862 VSS.n9861 0.0919286
R19484 VSS.n9638 VSS.n9479 0.0919286
R19485 VSS.n9487 VSS.n9485 0.0919286
R19486 VSS.n9646 VSS.n9645 0.0919286
R19487 VSS.n16671 VSS.n16670 0.0919286
R19488 VSS.n16685 VSS.n16346 0.0919286
R19489 VSS.n16715 VSS.n16714 0.0919286
R19490 VSS.n16754 VSS.n16318 0.0919286
R19491 VSS.n16805 VSS.n16804 0.0919286
R19492 VSS.n16567 VSS.n16566 0.0919286
R19493 VSS.n16581 VSS.n16421 0.0919286
R19494 VSS.n16589 VSS.n16588 0.0919286
R19495 VSS.n16078 VSS.n16077 0.0919286
R19496 VSS.n16092 VSS.n1518 0.0919286
R19497 VSS.n16122 VSS.n16121 0.0919286
R19498 VSS.n16161 VSS.n1490 0.0919286
R19499 VSS.n16212 VSS.n16211 0.0919286
R19500 VSS.n1732 VSS.n1731 0.0919286
R19501 VSS.n1746 VSS.n1586 0.0919286
R19502 VSS.n15996 VSS.n15995 0.0919286
R19503 VSS.n2057 VSS.n2056 0.0919286
R19504 VSS.n2065 VSS.n1983 0.0919286
R19505 VSS.n2307 VSS.n2306 0.0919286
R19506 VSS.n2268 VSS.n2267 0.0919286
R19507 VSS.n2186 VSS.n2157 0.0919286
R19508 VSS.n1930 VSS.n1771 0.0919286
R19509 VSS.n1779 VSS.n1777 0.0919286
R19510 VSS.n1938 VSS.n1937 0.0919286
R19511 VSS.n3219 VSS.n3218 0.0919286
R19512 VSS.n3233 VSS.n2895 0.0919286
R19513 VSS.n3263 VSS.n3262 0.0919286
R19514 VSS.n3302 VSS.n2867 0.0919286
R19515 VSS.n3353 VSS.n3352 0.0919286
R19516 VSS.n3129 VSS.n2970 0.0919286
R19517 VSS.n2978 VSS.n2976 0.0919286
R19518 VSS.n3137 VSS.n3136 0.0919286
R19519 VSS.n3811 VSS.n3810 0.0919286
R19520 VSS.n3825 VSS.n3487 0.0919286
R19521 VSS.n3855 VSS.n3854 0.0919286
R19522 VSS.n3894 VSS.n3459 0.0919286
R19523 VSS.n3945 VSS.n3944 0.0919286
R19524 VSS.n3721 VSS.n3562 0.0919286
R19525 VSS.n3570 VSS.n3568 0.0919286
R19526 VSS.n3729 VSS.n3728 0.0919286
R19527 VSS.n4403 VSS.n4402 0.0919286
R19528 VSS.n4417 VSS.n4079 0.0919286
R19529 VSS.n4447 VSS.n4446 0.0919286
R19530 VSS.n4486 VSS.n4051 0.0919286
R19531 VSS.n4537 VSS.n4536 0.0919286
R19532 VSS.n4313 VSS.n4154 0.0919286
R19533 VSS.n4162 VSS.n4160 0.0919286
R19534 VSS.n4321 VSS.n4320 0.0919286
R19535 VSS.n4995 VSS.n4994 0.0919286
R19536 VSS.n5009 VSS.n4671 0.0919286
R19537 VSS.n5039 VSS.n5038 0.0919286
R19538 VSS.n5078 VSS.n4643 0.0919286
R19539 VSS.n5129 VSS.n5128 0.0919286
R19540 VSS.n4905 VSS.n4746 0.0919286
R19541 VSS.n4754 VSS.n4752 0.0919286
R19542 VSS.n4913 VSS.n4912 0.0919286
R19543 VSS.n2653 VSS.n2652 0.0919286
R19544 VSS.n2661 VSS.n2579 0.0919286
R19545 VSS.n5272 VSS.n5271 0.0919286
R19546 VSS.n5233 VSS.n5232 0.0919286
R19547 VSS.n2782 VSS.n2753 0.0919286
R19548 VSS.n2526 VSS.n2367 0.0919286
R19549 VSS.n2375 VSS.n2373 0.0919286
R19550 VSS.n2534 VSS.n2533 0.0919286
R19551 VSS.n5614 VSS.n5613 0.0919286
R19552 VSS.n5622 VSS.n5540 0.0919286
R19553 VSS.n5845 VSS.n5844 0.0919286
R19554 VSS.n5806 VSS.n5805 0.0919286
R19555 VSS.n5756 VSS.n5714 0.0919286
R19556 VSS.n5487 VSS.n5328 0.0919286
R19557 VSS.n5336 VSS.n5334 0.0919286
R19558 VSS.n5495 VSS.n5494 0.0919286
R19559 VSS.n6187 VSS.n6186 0.0919286
R19560 VSS.n6195 VSS.n6113 0.0919286
R19561 VSS.n6437 VSS.n6436 0.0919286
R19562 VSS.n6398 VSS.n6397 0.0919286
R19563 VSS.n6316 VSS.n6287 0.0919286
R19564 VSS.n6060 VSS.n5901 0.0919286
R19565 VSS.n5909 VSS.n5907 0.0919286
R19566 VSS.n6068 VSS.n6067 0.0919286
R19567 VSS.n7952 VSS.n7951 0.0919286
R19568 VSS.n7966 VSS.n7628 0.0919286
R19569 VSS.n7996 VSS.n7995 0.0919286
R19570 VSS.n8035 VSS.n7600 0.0919286
R19571 VSS.n8086 VSS.n8085 0.0919286
R19572 VSS.n7862 VSS.n7703 0.0919286
R19573 VSS.n7711 VSS.n7709 0.0919286
R19574 VSS.n7870 VSS.n7869 0.0919286
R19575 VSS.n8544 VSS.n8543 0.0919286
R19576 VSS.n8558 VSS.n8220 0.0919286
R19577 VSS.n8588 VSS.n8587 0.0919286
R19578 VSS.n8627 VSS.n8192 0.0919286
R19579 VSS.n8678 VSS.n8677 0.0919286
R19580 VSS.n8454 VSS.n8295 0.0919286
R19581 VSS.n8303 VSS.n8301 0.0919286
R19582 VSS.n8462 VSS.n8461 0.0919286
R19583 VSS.n9136 VSS.n9135 0.0919286
R19584 VSS.n9150 VSS.n8812 0.0919286
R19585 VSS.n9180 VSS.n9179 0.0919286
R19586 VSS.n9219 VSS.n8784 0.0919286
R19587 VSS.n9270 VSS.n9269 0.0919286
R19588 VSS.n9046 VSS.n8887 0.0919286
R19589 VSS.n8895 VSS.n8893 0.0919286
R19590 VSS.n9054 VSS.n9053 0.0919286
R19591 VSS.n10320 VSS.n10319 0.0919286
R19592 VSS.n10334 VSS.n9996 0.0919286
R19593 VSS.n10364 VSS.n10363 0.0919286
R19594 VSS.n10403 VSS.n9968 0.0919286
R19595 VSS.n10454 VSS.n10453 0.0919286
R19596 VSS.n10230 VSS.n10071 0.0919286
R19597 VSS.n10079 VSS.n10077 0.0919286
R19598 VSS.n10238 VSS.n10237 0.0919286
R19599 VSS.n10912 VSS.n10911 0.0919286
R19600 VSS.n10926 VSS.n10588 0.0919286
R19601 VSS.n10956 VSS.n10955 0.0919286
R19602 VSS.n10995 VSS.n10560 0.0919286
R19603 VSS.n11046 VSS.n11045 0.0919286
R19604 VSS.n10822 VSS.n10663 0.0919286
R19605 VSS.n10671 VSS.n10669 0.0919286
R19606 VSS.n10830 VSS.n10829 0.0919286
R19607 VSS.n11504 VSS.n11503 0.0919286
R19608 VSS.n11518 VSS.n11180 0.0919286
R19609 VSS.n11548 VSS.n11547 0.0919286
R19610 VSS.n11587 VSS.n11152 0.0919286
R19611 VSS.n11638 VSS.n11637 0.0919286
R19612 VSS.n11414 VSS.n11255 0.0919286
R19613 VSS.n11263 VSS.n11261 0.0919286
R19614 VSS.n11422 VSS.n11421 0.0919286
R19615 VSS.n12096 VSS.n12095 0.0919286
R19616 VSS.n12110 VSS.n11772 0.0919286
R19617 VSS.n12140 VSS.n12139 0.0919286
R19618 VSS.n12179 VSS.n11744 0.0919286
R19619 VSS.n12230 VSS.n12229 0.0919286
R19620 VSS.n12006 VSS.n11847 0.0919286
R19621 VSS.n11855 VSS.n11853 0.0919286
R19622 VSS.n12014 VSS.n12013 0.0919286
R19623 VSS.n12688 VSS.n12687 0.0919286
R19624 VSS.n12702 VSS.n12364 0.0919286
R19625 VSS.n12732 VSS.n12731 0.0919286
R19626 VSS.n12771 VSS.n12336 0.0919286
R19627 VSS.n12822 VSS.n12821 0.0919286
R19628 VSS.n12598 VSS.n12439 0.0919286
R19629 VSS.n12447 VSS.n12445 0.0919286
R19630 VSS.n12606 VSS.n12605 0.0919286
R19631 VSS.n13280 VSS.n13279 0.0919286
R19632 VSS.n13294 VSS.n12956 0.0919286
R19633 VSS.n13324 VSS.n13323 0.0919286
R19634 VSS.n13363 VSS.n12928 0.0919286
R19635 VSS.n13414 VSS.n13413 0.0919286
R19636 VSS.n13190 VSS.n13031 0.0919286
R19637 VSS.n13039 VSS.n13037 0.0919286
R19638 VSS.n13198 VSS.n13197 0.0919286
R19639 VSS.n13872 VSS.n13871 0.0919286
R19640 VSS.n13886 VSS.n13548 0.0919286
R19641 VSS.n13916 VSS.n13915 0.0919286
R19642 VSS.n13955 VSS.n13520 0.0919286
R19643 VSS.n14006 VSS.n14005 0.0919286
R19644 VSS.n13782 VSS.n13623 0.0919286
R19645 VSS.n13631 VSS.n13629 0.0919286
R19646 VSS.n13790 VSS.n13789 0.0919286
R19647 VSS.n14464 VSS.n14463 0.0919286
R19648 VSS.n14478 VSS.n14140 0.0919286
R19649 VSS.n14508 VSS.n14507 0.0919286
R19650 VSS.n14547 VSS.n14112 0.0919286
R19651 VSS.n14598 VSS.n14597 0.0919286
R19652 VSS.n14374 VSS.n14215 0.0919286
R19653 VSS.n14223 VSS.n14221 0.0919286
R19654 VSS.n14382 VSS.n14381 0.0919286
R19655 VSS.n15056 VSS.n15055 0.0919286
R19656 VSS.n15070 VSS.n14732 0.0919286
R19657 VSS.n15100 VSS.n15099 0.0919286
R19658 VSS.n15139 VSS.n14704 0.0919286
R19659 VSS.n15190 VSS.n15189 0.0919286
R19660 VSS.n14966 VSS.n14807 0.0919286
R19661 VSS.n14815 VSS.n14813 0.0919286
R19662 VSS.n14974 VSS.n14973 0.0919286
R19663 VSS.n15648 VSS.n15647 0.0919286
R19664 VSS.n15662 VSS.n15324 0.0919286
R19665 VSS.n15692 VSS.n15691 0.0919286
R19666 VSS.n15731 VSS.n15296 0.0919286
R19667 VSS.n15782 VSS.n15781 0.0919286
R19668 VSS.n15558 VSS.n15399 0.0919286
R19669 VSS.n15407 VSS.n15405 0.0919286
R19670 VSS.n15566 VSS.n15565 0.0919286
R19671 VSS.n6793 VSS.n6792 0.0919286
R19672 VSS.n6801 VSS.n6719 0.0919286
R19673 VSS.n15925 VSS.n15924 0.0919286
R19674 VSS.n15886 VSS.n15885 0.0919286
R19675 VSS.n6922 VSS.n6893 0.0919286
R19676 VSS.n6666 VSS.n6507 0.0919286
R19677 VSS.n6515 VSS.n6513 0.0919286
R19678 VSS.n6674 VSS.n6673 0.0919286
R19679 VSS.n7360 VSS.n7359 0.0919286
R19680 VSS.n7374 VSS.n7035 0.0919286
R19681 VSS.n7404 VSS.n7403 0.0919286
R19682 VSS.n7443 VSS.n7007 0.0919286
R19683 VSS.n7494 VSS.n7493 0.0919286
R19684 VSS.n7256 VSS.n7255 0.0919286
R19685 VSS.n7270 VSS.n7110 0.0919286
R19686 VSS.n7278 VSS.n7277 0.0919286
R19687 VSS.n18672 VSS.n18671 0.0919286
R19688 VSS.n18686 VSS.n133 0.0919286
R19689 VSS.n18716 VSS.n18715 0.0919286
R19690 VSS.n18755 VSS.n105 0.0919286
R19691 VSS.n18806 VSS.n18805 0.0919286
R19692 VSS.n396 VSS.n328 0.0919286
R19693 VSS.n405 VSS.n404 0.0919286
R19694 VSS.n18590 VSS.n18589 0.0919286
R19695 VSS.n616 VSS.n615 0.0919286
R19696 VSS.n624 VSS.n539 0.0919286
R19697 VSS.n839 VSS.n838 0.0919286
R19698 VSS.n800 VSS.n799 0.0919286
R19699 VSS.n754 VSS.n716 0.0919286
R19700 VSS.n960 VSS.n959 0.0919286
R19701 VSS.n968 VSS.n886 0.0919286
R19702 VSS.n976 VSS.n975 0.0919286
R19703 VSS.n17914 VSS.n17913 0.0919286
R19704 VSS.n1404 VSS.n1375 0.0919286
R19705 VSS.n18037 VSS.n18036 0.024
R19706 VSS.n18007 VSS.n18006 0.024
R19707 VSS.n17021 VSS.n17020 0.024
R19708 VSS.n17092 VSS.n17091 0.024
R19709 VSS.n17515 VSS.n17514 0.024
R19710 VSS.n17577 VSS.n17576 0.024
R19711 VSS.n17613 VSS.n17612 0.024
R19712 VSS.n17684 VSS.n17683 0.024
R19713 VSS.n18092 VSS.n18091 0.024
R19714 VSS.n18154 VSS.n18153 0.024
R19715 VSS.n18577 VSS.n18576 0.024
R19716 VSS.n18547 VSS.n18546 0.024
R19717 VSS.n9663 VSS.n9662 0.024
R19718 VSS.n9734 VSS.n9733 0.024
R19719 VSS.n16501 VSS.n16500 0.024
R19720 VSS.n16573 VSS.n16572 0.024
R19721 VSS.n16606 VSS.n16605 0.024
R19722 VSS.n16677 VSS.n16676 0.024
R19723 VSS.n1666 VSS.n1665 0.024
R19724 VSS.n1738 VSS.n1737 0.024
R19725 VSS.n16013 VSS.n16012 0.024
R19726 VSS.n16084 VSS.n16083 0.024
R19727 VSS.n1857 VSS.n1856 0.024
R19728 VSS.n1919 VSS.n1918 0.024
R19729 VSS.n2342 VSS.n2341 0.024
R19730 VSS.n2312 VSS.n2311 0.024
R19731 VSS.n3056 VSS.n3055 0.024
R19732 VSS.n3118 VSS.n3117 0.024
R19733 VSS.n3154 VSS.n3153 0.024
R19734 VSS.n3225 VSS.n3224 0.024
R19735 VSS.n3648 VSS.n3647 0.024
R19736 VSS.n3710 VSS.n3709 0.024
R19737 VSS.n3746 VSS.n3745 0.024
R19738 VSS.n3817 VSS.n3816 0.024
R19739 VSS.n4240 VSS.n4239 0.024
R19740 VSS.n4302 VSS.n4301 0.024
R19741 VSS.n4338 VSS.n4337 0.024
R19742 VSS.n4409 VSS.n4408 0.024
R19743 VSS.n4832 VSS.n4831 0.024
R19744 VSS.n4894 VSS.n4893 0.024
R19745 VSS.n4930 VSS.n4929 0.024
R19746 VSS.n5001 VSS.n5000 0.024
R19747 VSS.n2453 VSS.n2452 0.024
R19748 VSS.n2515 VSS.n2514 0.024
R19749 VSS.n5307 VSS.n5306 0.024
R19750 VSS.n5277 VSS.n5276 0.024
R19751 VSS.n5414 VSS.n5413 0.024
R19752 VSS.n5476 VSS.n5475 0.024
R19753 VSS.n5880 VSS.n5879 0.024
R19754 VSS.n5850 VSS.n5849 0.024
R19755 VSS.n5987 VSS.n5986 0.024
R19756 VSS.n6049 VSS.n6048 0.024
R19757 VSS.n6472 VSS.n6471 0.024
R19758 VSS.n6442 VSS.n6441 0.024
R19759 VSS.n7789 VSS.n7788 0.024
R19760 VSS.n7851 VSS.n7850 0.024
R19761 VSS.n7887 VSS.n7886 0.024
R19762 VSS.n7958 VSS.n7957 0.024
R19763 VSS.n8381 VSS.n8380 0.024
R19764 VSS.n8443 VSS.n8442 0.024
R19765 VSS.n8479 VSS.n8478 0.024
R19766 VSS.n8550 VSS.n8549 0.024
R19767 VSS.n8973 VSS.n8972 0.024
R19768 VSS.n9035 VSS.n9034 0.024
R19769 VSS.n9071 VSS.n9070 0.024
R19770 VSS.n9142 VSS.n9141 0.024
R19771 VSS.n10157 VSS.n10156 0.024
R19772 VSS.n10219 VSS.n10218 0.024
R19773 VSS.n10255 VSS.n10254 0.024
R19774 VSS.n10326 VSS.n10325 0.024
R19775 VSS.n10749 VSS.n10748 0.024
R19776 VSS.n10811 VSS.n10810 0.024
R19777 VSS.n10847 VSS.n10846 0.024
R19778 VSS.n10918 VSS.n10917 0.024
R19779 VSS.n11341 VSS.n11340 0.024
R19780 VSS.n11403 VSS.n11402 0.024
R19781 VSS.n11439 VSS.n11438 0.024
R19782 VSS.n11510 VSS.n11509 0.024
R19783 VSS.n11933 VSS.n11932 0.024
R19784 VSS.n11995 VSS.n11994 0.024
R19785 VSS.n12031 VSS.n12030 0.024
R19786 VSS.n12102 VSS.n12101 0.024
R19787 VSS.n12525 VSS.n12524 0.024
R19788 VSS.n12587 VSS.n12586 0.024
R19789 VSS.n12623 VSS.n12622 0.024
R19790 VSS.n12694 VSS.n12693 0.024
R19791 VSS.n13117 VSS.n13116 0.024
R19792 VSS.n13179 VSS.n13178 0.024
R19793 VSS.n13215 VSS.n13214 0.024
R19794 VSS.n13286 VSS.n13285 0.024
R19795 VSS.n13709 VSS.n13708 0.024
R19796 VSS.n13771 VSS.n13770 0.024
R19797 VSS.n13807 VSS.n13806 0.024
R19798 VSS.n13878 VSS.n13877 0.024
R19799 VSS.n14301 VSS.n14300 0.024
R19800 VSS.n14363 VSS.n14362 0.024
R19801 VSS.n14399 VSS.n14398 0.024
R19802 VSS.n14470 VSS.n14469 0.024
R19803 VSS.n14893 VSS.n14892 0.024
R19804 VSS.n14955 VSS.n14954 0.024
R19805 VSS.n14991 VSS.n14990 0.024
R19806 VSS.n15062 VSS.n15061 0.024
R19807 VSS.n15485 VSS.n15484 0.024
R19808 VSS.n15547 VSS.n15546 0.024
R19809 VSS.n15583 VSS.n15582 0.024
R19810 VSS.n15654 VSS.n15653 0.024
R19811 VSS.n6593 VSS.n6592 0.024
R19812 VSS.n6655 VSS.n6654 0.024
R19813 VSS.n15960 VSS.n15959 0.024
R19814 VSS.n15930 VSS.n15929 0.024
R19815 VSS.n7190 VSS.n7189 0.024
R19816 VSS.n7262 VSS.n7261 0.024
R19817 VSS.n7295 VSS.n7294 0.024
R19818 VSS.n7366 VSS.n7365 0.024
R19819 VSS.n446 VSS.n445 0.024
R19820 VSS.n416 VSS.n415 0.024
R19821 VSS.n18607 VSS.n18606 0.024
R19822 VSS.n18678 VSS.n18677 0.024
R19823 VSS.n1011 VSS.n1010 0.024
R19824 VSS.n981 VSS.n980 0.024
R19825 VSS.n874 VSS.n873 0.024
R19826 VSS.n844 VSS.n843 0.024
R19827 VSS.n17988 VSS.n17987 0.024
R19828 VSS.n17958 VSS.n17957 0.024
R19829 VSS.n9565 VSS.n9564 0.0238333
R19830 VSS.n9627 VSS.n9626 0.0238333
R19831 VSS.n17977 VSS.n17976 0.0228214
R19832 VSS.n17969 VSS.n17968 0.0228214
R19833 VSS.n17961 VSS.n1188 0.0228214
R19834 VSS.n1000 VSS.n999 0.0228214
R19835 VSS.n992 VSS.n991 0.0228214
R19836 VSS.n984 VSS.n487 0.0228214
R19837 VSS.n16980 VSS.n16969 0.0228214
R19838 VSS.n17065 VSS.n17064 0.0228214
R19839 VSS.n17073 VSS.n16947 0.0228214
R19840 VSS.n18026 VSS.n18025 0.0228214
R19841 VSS.n18018 VSS.n18017 0.0228214
R19842 VSS.n18010 VSS.n1054 0.0228214
R19843 VSS.n17204 VSS.n16890 0.0228214
R19844 VSS.n17394 VSS.n17383 0.0228214
R19845 VSS.n17657 VSS.n17656 0.0228214
R19846 VSS.n17665 VSS.n17361 0.0228214
R19847 VSS.n17543 VSS.n17542 0.0228214
R19848 VSS.n17464 VSS.n17446 0.0228214
R19849 VSS.n17573 VSS.n17441 0.0228214
R19850 VSS.n17796 VSS.n17304 0.0228214
R19851 VSS.n18120 VSS.n18119 0.0228214
R19852 VSS.n256 VSS.n238 0.0228214
R19853 VSS.n18150 VSS.n233 0.0228214
R19854 VSS.n18566 VSS.n18565 0.0228214
R19855 VSS.n18558 VSS.n18557 0.0228214
R19856 VSS.n18550 VSS.n18205 0.0228214
R19857 VSS.n18489 VSS.n18388 0.0228214
R19858 VSS.n9593 VSS.n9592 0.0228214
R19859 VSS.n9514 VSS.n9496 0.0228214
R19860 VSS.n9623 VSS.n9491 0.0228214
R19861 VSS.n9444 VSS.n9433 0.0228214
R19862 VSS.n9707 VSS.n9706 0.0228214
R19863 VSS.n9715 VSS.n9411 0.0228214
R19864 VSS.n9846 VSS.n9354 0.0228214
R19865 VSS.n16463 VSS.n16450 0.0228214
R19866 VSS.n16545 VSS.n16544 0.0228214
R19867 VSS.n16553 VSS.n16428 0.0228214
R19868 VSS.n16386 VSS.n16375 0.0228214
R19869 VSS.n16650 VSS.n16649 0.0228214
R19870 VSS.n16658 VSS.n16353 0.0228214
R19871 VSS.n16789 VSS.n16296 0.0228214
R19872 VSS.n1628 VSS.n1615 0.0228214
R19873 VSS.n1710 VSS.n1709 0.0228214
R19874 VSS.n1718 VSS.n1593 0.0228214
R19875 VSS.n1558 VSS.n1547 0.0228214
R19876 VSS.n16057 VSS.n16056 0.0228214
R19877 VSS.n16065 VSS.n1525 0.0228214
R19878 VSS.n16196 VSS.n1468 0.0228214
R19879 VSS.n1885 VSS.n1884 0.0228214
R19880 VSS.n1806 VSS.n1788 0.0228214
R19881 VSS.n1915 VSS.n1783 0.0228214
R19882 VSS.n2331 VSS.n2330 0.0228214
R19883 VSS.n2323 VSS.n2322 0.0228214
R19884 VSS.n2315 VSS.n1970 0.0228214
R19885 VSS.n2252 VSS.n2251 0.0228214
R19886 VSS.n3084 VSS.n3083 0.0228214
R19887 VSS.n3005 VSS.n2987 0.0228214
R19888 VSS.n3114 VSS.n2982 0.0228214
R19889 VSS.n2935 VSS.n2924 0.0228214
R19890 VSS.n3198 VSS.n3197 0.0228214
R19891 VSS.n3206 VSS.n2902 0.0228214
R19892 VSS.n3337 VSS.n2845 0.0228214
R19893 VSS.n3676 VSS.n3675 0.0228214
R19894 VSS.n3597 VSS.n3579 0.0228214
R19895 VSS.n3706 VSS.n3574 0.0228214
R19896 VSS.n3527 VSS.n3516 0.0228214
R19897 VSS.n3790 VSS.n3789 0.0228214
R19898 VSS.n3798 VSS.n3494 0.0228214
R19899 VSS.n3929 VSS.n3437 0.0228214
R19900 VSS.n4268 VSS.n4267 0.0228214
R19901 VSS.n4189 VSS.n4171 0.0228214
R19902 VSS.n4298 VSS.n4166 0.0228214
R19903 VSS.n4119 VSS.n4108 0.0228214
R19904 VSS.n4382 VSS.n4381 0.0228214
R19905 VSS.n4390 VSS.n4086 0.0228214
R19906 VSS.n4521 VSS.n4029 0.0228214
R19907 VSS.n4860 VSS.n4859 0.0228214
R19908 VSS.n4781 VSS.n4763 0.0228214
R19909 VSS.n4890 VSS.n4758 0.0228214
R19910 VSS.n4711 VSS.n4700 0.0228214
R19911 VSS.n4974 VSS.n4973 0.0228214
R19912 VSS.n4982 VSS.n4678 0.0228214
R19913 VSS.n5113 VSS.n4621 0.0228214
R19914 VSS.n2481 VSS.n2480 0.0228214
R19915 VSS.n2402 VSS.n2384 0.0228214
R19916 VSS.n2511 VSS.n2379 0.0228214
R19917 VSS.n5296 VSS.n5295 0.0228214
R19918 VSS.n5288 VSS.n5287 0.0228214
R19919 VSS.n5280 VSS.n2566 0.0228214
R19920 VSS.n5217 VSS.n5216 0.0228214
R19921 VSS.n5442 VSS.n5441 0.0228214
R19922 VSS.n5363 VSS.n5345 0.0228214
R19923 VSS.n5472 VSS.n5340 0.0228214
R19924 VSS.n5869 VSS.n5868 0.0228214
R19925 VSS.n5861 VSS.n5860 0.0228214
R19926 VSS.n5853 VSS.n5527 0.0228214
R19927 VSS.n5790 VSS.n5789 0.0228214
R19928 VSS.n6015 VSS.n6014 0.0228214
R19929 VSS.n5936 VSS.n5918 0.0228214
R19930 VSS.n6045 VSS.n5913 0.0228214
R19931 VSS.n6461 VSS.n6460 0.0228214
R19932 VSS.n6453 VSS.n6452 0.0228214
R19933 VSS.n6445 VSS.n6100 0.0228214
R19934 VSS.n6382 VSS.n6381 0.0228214
R19935 VSS.n7817 VSS.n7816 0.0228214
R19936 VSS.n7738 VSS.n7720 0.0228214
R19937 VSS.n7847 VSS.n7715 0.0228214
R19938 VSS.n7668 VSS.n7657 0.0228214
R19939 VSS.n7931 VSS.n7930 0.0228214
R19940 VSS.n7939 VSS.n7635 0.0228214
R19941 VSS.n8070 VSS.n7578 0.0228214
R19942 VSS.n8409 VSS.n8408 0.0228214
R19943 VSS.n8330 VSS.n8312 0.0228214
R19944 VSS.n8439 VSS.n8307 0.0228214
R19945 VSS.n8260 VSS.n8249 0.0228214
R19946 VSS.n8523 VSS.n8522 0.0228214
R19947 VSS.n8531 VSS.n8227 0.0228214
R19948 VSS.n8662 VSS.n8170 0.0228214
R19949 VSS.n9001 VSS.n9000 0.0228214
R19950 VSS.n8922 VSS.n8904 0.0228214
R19951 VSS.n9031 VSS.n8899 0.0228214
R19952 VSS.n8852 VSS.n8841 0.0228214
R19953 VSS.n9115 VSS.n9114 0.0228214
R19954 VSS.n9123 VSS.n8819 0.0228214
R19955 VSS.n9254 VSS.n8762 0.0228214
R19956 VSS.n10185 VSS.n10184 0.0228214
R19957 VSS.n10106 VSS.n10088 0.0228214
R19958 VSS.n10215 VSS.n10083 0.0228214
R19959 VSS.n10036 VSS.n10025 0.0228214
R19960 VSS.n10299 VSS.n10298 0.0228214
R19961 VSS.n10307 VSS.n10003 0.0228214
R19962 VSS.n10438 VSS.n9946 0.0228214
R19963 VSS.n10777 VSS.n10776 0.0228214
R19964 VSS.n10698 VSS.n10680 0.0228214
R19965 VSS.n10807 VSS.n10675 0.0228214
R19966 VSS.n10628 VSS.n10617 0.0228214
R19967 VSS.n10891 VSS.n10890 0.0228214
R19968 VSS.n10899 VSS.n10595 0.0228214
R19969 VSS.n11030 VSS.n10538 0.0228214
R19970 VSS.n11369 VSS.n11368 0.0228214
R19971 VSS.n11290 VSS.n11272 0.0228214
R19972 VSS.n11399 VSS.n11267 0.0228214
R19973 VSS.n11220 VSS.n11209 0.0228214
R19974 VSS.n11483 VSS.n11482 0.0228214
R19975 VSS.n11491 VSS.n11187 0.0228214
R19976 VSS.n11622 VSS.n11130 0.0228214
R19977 VSS.n11961 VSS.n11960 0.0228214
R19978 VSS.n11882 VSS.n11864 0.0228214
R19979 VSS.n11991 VSS.n11859 0.0228214
R19980 VSS.n11812 VSS.n11801 0.0228214
R19981 VSS.n12075 VSS.n12074 0.0228214
R19982 VSS.n12083 VSS.n11779 0.0228214
R19983 VSS.n12214 VSS.n11722 0.0228214
R19984 VSS.n12553 VSS.n12552 0.0228214
R19985 VSS.n12474 VSS.n12456 0.0228214
R19986 VSS.n12583 VSS.n12451 0.0228214
R19987 VSS.n12404 VSS.n12393 0.0228214
R19988 VSS.n12667 VSS.n12666 0.0228214
R19989 VSS.n12675 VSS.n12371 0.0228214
R19990 VSS.n12806 VSS.n12314 0.0228214
R19991 VSS.n13145 VSS.n13144 0.0228214
R19992 VSS.n13066 VSS.n13048 0.0228214
R19993 VSS.n13175 VSS.n13043 0.0228214
R19994 VSS.n12996 VSS.n12985 0.0228214
R19995 VSS.n13259 VSS.n13258 0.0228214
R19996 VSS.n13267 VSS.n12963 0.0228214
R19997 VSS.n13398 VSS.n12906 0.0228214
R19998 VSS.n13737 VSS.n13736 0.0228214
R19999 VSS.n13658 VSS.n13640 0.0228214
R20000 VSS.n13767 VSS.n13635 0.0228214
R20001 VSS.n13588 VSS.n13577 0.0228214
R20002 VSS.n13851 VSS.n13850 0.0228214
R20003 VSS.n13859 VSS.n13555 0.0228214
R20004 VSS.n13990 VSS.n13498 0.0228214
R20005 VSS.n14329 VSS.n14328 0.0228214
R20006 VSS.n14250 VSS.n14232 0.0228214
R20007 VSS.n14359 VSS.n14227 0.0228214
R20008 VSS.n14180 VSS.n14169 0.0228214
R20009 VSS.n14443 VSS.n14442 0.0228214
R20010 VSS.n14451 VSS.n14147 0.0228214
R20011 VSS.n14582 VSS.n14090 0.0228214
R20012 VSS.n14921 VSS.n14920 0.0228214
R20013 VSS.n14842 VSS.n14824 0.0228214
R20014 VSS.n14951 VSS.n14819 0.0228214
R20015 VSS.n14772 VSS.n14761 0.0228214
R20016 VSS.n15035 VSS.n15034 0.0228214
R20017 VSS.n15043 VSS.n14739 0.0228214
R20018 VSS.n15174 VSS.n14682 0.0228214
R20019 VSS.n15513 VSS.n15512 0.0228214
R20020 VSS.n15434 VSS.n15416 0.0228214
R20021 VSS.n15543 VSS.n15411 0.0228214
R20022 VSS.n15364 VSS.n15353 0.0228214
R20023 VSS.n15627 VSS.n15626 0.0228214
R20024 VSS.n15635 VSS.n15331 0.0228214
R20025 VSS.n15766 VSS.n15274 0.0228214
R20026 VSS.n6621 VSS.n6620 0.0228214
R20027 VSS.n6542 VSS.n6524 0.0228214
R20028 VSS.n6651 VSS.n6519 0.0228214
R20029 VSS.n15949 VSS.n15948 0.0228214
R20030 VSS.n15941 VSS.n15940 0.0228214
R20031 VSS.n15933 VSS.n6706 0.0228214
R20032 VSS.n15870 VSS.n15869 0.0228214
R20033 VSS.n7152 VSS.n7139 0.0228214
R20034 VSS.n7234 VSS.n7233 0.0228214
R20035 VSS.n7242 VSS.n7117 0.0228214
R20036 VSS.n7075 VSS.n7064 0.0228214
R20037 VSS.n7339 VSS.n7338 0.0228214
R20038 VSS.n7347 VSS.n7042 0.0228214
R20039 VSS.n7478 VSS.n6985 0.0228214
R20040 VSS.n435 VSS.n434 0.0228214
R20041 VSS.n427 VSS.n426 0.0228214
R20042 VSS.n419 VSS.n321 0.0228214
R20043 VSS.n173 VSS.n162 0.0228214
R20044 VSS.n18651 VSS.n18650 0.0228214
R20045 VSS.n18659 VSS.n140 0.0228214
R20046 VSS.n18790 VSS.n83 0.0228214
R20047 VSS.n863 VSS.n862 0.0228214
R20048 VSS.n855 VSS.n854 0.0228214
R20049 VSS.n847 VSS.n526 0.0228214
R20050 VSS.n784 VSS.n783 0.0228214
R20051 VSS.n17898 VSS.n17897 0.0228214
R20052 VSS.n17984 VSS.n1166 0.0210357
R20053 VSS.n1007 VSS.n464 0.0210357
R20054 VSS.n16993 VSS.n16985 0.0210357
R20055 VSS.n18033 VSS.n1031 0.0210357
R20056 VSS.n17171 VSS.n16911 0.0210357
R20057 VSS.n17211 VSS.n16897 0.0210357
R20058 VSS.n17210 VSS.n16899 0.0210357
R20059 VSS.n17407 VSS.n17399 0.0210357
R20060 VSS.n17487 VSS.n17486 0.0210357
R20061 VSS.n17763 VSS.n17325 0.0210357
R20062 VSS.n17803 VSS.n17311 0.0210357
R20063 VSS.n17802 VSS.n17313 0.0210357
R20064 VSS.n279 VSS.n278 0.0210357
R20065 VSS.n18573 VSS.n18183 0.0210357
R20066 VSS.n18508 VSS.n18507 0.0210357
R20067 VSS.n18401 VSS.n18356 0.0210357
R20068 VSS.n18400 VSS.n18354 0.0210357
R20069 VSS.n9537 VSS.n9536 0.0210357
R20070 VSS.n9457 VSS.n9449 0.0210357
R20071 VSS.n9813 VSS.n9375 0.0210357
R20072 VSS.n9853 VSS.n9361 0.0210357
R20073 VSS.n9852 VSS.n9363 0.0210357
R20074 VSS.n16474 VSS.n16467 0.0210357
R20075 VSS.n16399 VSS.n16391 0.0210357
R20076 VSS.n16756 VSS.n16317 0.0210357
R20077 VSS.n16796 VSS.n16303 0.0210357
R20078 VSS.n16795 VSS.n16305 0.0210357
R20079 VSS.n1639 VSS.n1632 0.0210357
R20080 VSS.n1571 VSS.n1563 0.0210357
R20081 VSS.n16163 VSS.n1489 0.0210357
R20082 VSS.n16203 VSS.n1475 0.0210357
R20083 VSS.n16202 VSS.n1477 0.0210357
R20084 VSS.n1829 VSS.n1828 0.0210357
R20085 VSS.n2338 VSS.n1948 0.0210357
R20086 VSS.n2270 VSS.n2120 0.0210357
R20087 VSS.n2259 VSS.n2127 0.0210357
R20088 VSS.n2258 VSS.n2129 0.0210357
R20089 VSS.n3028 VSS.n3027 0.0210357
R20090 VSS.n2948 VSS.n2940 0.0210357
R20091 VSS.n3304 VSS.n2866 0.0210357
R20092 VSS.n3344 VSS.n2852 0.0210357
R20093 VSS.n3343 VSS.n2854 0.0210357
R20094 VSS.n3620 VSS.n3619 0.0210357
R20095 VSS.n3540 VSS.n3532 0.0210357
R20096 VSS.n3896 VSS.n3458 0.0210357
R20097 VSS.n3936 VSS.n3444 0.0210357
R20098 VSS.n3935 VSS.n3446 0.0210357
R20099 VSS.n4212 VSS.n4211 0.0210357
R20100 VSS.n4132 VSS.n4124 0.0210357
R20101 VSS.n4488 VSS.n4050 0.0210357
R20102 VSS.n4528 VSS.n4036 0.0210357
R20103 VSS.n4527 VSS.n4038 0.0210357
R20104 VSS.n4804 VSS.n4803 0.0210357
R20105 VSS.n4724 VSS.n4716 0.0210357
R20106 VSS.n5080 VSS.n4642 0.0210357
R20107 VSS.n5120 VSS.n4628 0.0210357
R20108 VSS.n5119 VSS.n4630 0.0210357
R20109 VSS.n2425 VSS.n2424 0.0210357
R20110 VSS.n5303 VSS.n2544 0.0210357
R20111 VSS.n5235 VSS.n2716 0.0210357
R20112 VSS.n5224 VSS.n2723 0.0210357
R20113 VSS.n5223 VSS.n2725 0.0210357
R20114 VSS.n5386 VSS.n5385 0.0210357
R20115 VSS.n5876 VSS.n5505 0.0210357
R20116 VSS.n5808 VSS.n5677 0.0210357
R20117 VSS.n5797 VSS.n5684 0.0210357
R20118 VSS.n5796 VSS.n5686 0.0210357
R20119 VSS.n5959 VSS.n5958 0.0210357
R20120 VSS.n6468 VSS.n6078 0.0210357
R20121 VSS.n6400 VSS.n6250 0.0210357
R20122 VSS.n6389 VSS.n6257 0.0210357
R20123 VSS.n6388 VSS.n6259 0.0210357
R20124 VSS.n7761 VSS.n7760 0.0210357
R20125 VSS.n7681 VSS.n7673 0.0210357
R20126 VSS.n8037 VSS.n7599 0.0210357
R20127 VSS.n8077 VSS.n7585 0.0210357
R20128 VSS.n8076 VSS.n7587 0.0210357
R20129 VSS.n8353 VSS.n8352 0.0210357
R20130 VSS.n8273 VSS.n8265 0.0210357
R20131 VSS.n8629 VSS.n8191 0.0210357
R20132 VSS.n8669 VSS.n8177 0.0210357
R20133 VSS.n8668 VSS.n8179 0.0210357
R20134 VSS.n8945 VSS.n8944 0.0210357
R20135 VSS.n8865 VSS.n8857 0.0210357
R20136 VSS.n9221 VSS.n8783 0.0210357
R20137 VSS.n9261 VSS.n8769 0.0210357
R20138 VSS.n9260 VSS.n8771 0.0210357
R20139 VSS.n10129 VSS.n10128 0.0210357
R20140 VSS.n10049 VSS.n10041 0.0210357
R20141 VSS.n10405 VSS.n9967 0.0210357
R20142 VSS.n10445 VSS.n9953 0.0210357
R20143 VSS.n10444 VSS.n9955 0.0210357
R20144 VSS.n10721 VSS.n10720 0.0210357
R20145 VSS.n10641 VSS.n10633 0.0210357
R20146 VSS.n10997 VSS.n10559 0.0210357
R20147 VSS.n11037 VSS.n10545 0.0210357
R20148 VSS.n11036 VSS.n10547 0.0210357
R20149 VSS.n11313 VSS.n11312 0.0210357
R20150 VSS.n11233 VSS.n11225 0.0210357
R20151 VSS.n11589 VSS.n11151 0.0210357
R20152 VSS.n11629 VSS.n11137 0.0210357
R20153 VSS.n11628 VSS.n11139 0.0210357
R20154 VSS.n11905 VSS.n11904 0.0210357
R20155 VSS.n11825 VSS.n11817 0.0210357
R20156 VSS.n12181 VSS.n11743 0.0210357
R20157 VSS.n12221 VSS.n11729 0.0210357
R20158 VSS.n12220 VSS.n11731 0.0210357
R20159 VSS.n12497 VSS.n12496 0.0210357
R20160 VSS.n12417 VSS.n12409 0.0210357
R20161 VSS.n12773 VSS.n12335 0.0210357
R20162 VSS.n12813 VSS.n12321 0.0210357
R20163 VSS.n12812 VSS.n12323 0.0210357
R20164 VSS.n13089 VSS.n13088 0.0210357
R20165 VSS.n13009 VSS.n13001 0.0210357
R20166 VSS.n13365 VSS.n12927 0.0210357
R20167 VSS.n13405 VSS.n12913 0.0210357
R20168 VSS.n13404 VSS.n12915 0.0210357
R20169 VSS.n13681 VSS.n13680 0.0210357
R20170 VSS.n13601 VSS.n13593 0.0210357
R20171 VSS.n13957 VSS.n13519 0.0210357
R20172 VSS.n13997 VSS.n13505 0.0210357
R20173 VSS.n13996 VSS.n13507 0.0210357
R20174 VSS.n14273 VSS.n14272 0.0210357
R20175 VSS.n14193 VSS.n14185 0.0210357
R20176 VSS.n14549 VSS.n14111 0.0210357
R20177 VSS.n14589 VSS.n14097 0.0210357
R20178 VSS.n14588 VSS.n14099 0.0210357
R20179 VSS.n14865 VSS.n14864 0.0210357
R20180 VSS.n14785 VSS.n14777 0.0210357
R20181 VSS.n15141 VSS.n14703 0.0210357
R20182 VSS.n15181 VSS.n14689 0.0210357
R20183 VSS.n15180 VSS.n14691 0.0210357
R20184 VSS.n15457 VSS.n15456 0.0210357
R20185 VSS.n15377 VSS.n15369 0.0210357
R20186 VSS.n15733 VSS.n15295 0.0210357
R20187 VSS.n15773 VSS.n15281 0.0210357
R20188 VSS.n15772 VSS.n15283 0.0210357
R20189 VSS.n6565 VSS.n6564 0.0210357
R20190 VSS.n15956 VSS.n6684 0.0210357
R20191 VSS.n15888 VSS.n6856 0.0210357
R20192 VSS.n15877 VSS.n6863 0.0210357
R20193 VSS.n15876 VSS.n6865 0.0210357
R20194 VSS.n7163 VSS.n7156 0.0210357
R20195 VSS.n7088 VSS.n7080 0.0210357
R20196 VSS.n7445 VSS.n7006 0.0210357
R20197 VSS.n7485 VSS.n6992 0.0210357
R20198 VSS.n7484 VSS.n6994 0.0210357
R20199 VSS.n442 VSS.n298 0.0210357
R20200 VSS.n186 VSS.n178 0.0210357
R20201 VSS.n18757 VSS.n104 0.0210357
R20202 VSS.n18797 VSS.n90 0.0210357
R20203 VSS.n18796 VSS.n92 0.0210357
R20204 VSS.n870 VSS.n504 0.0210357
R20205 VSS.n802 VSS.n679 0.0210357
R20206 VSS.n791 VSS.n686 0.0210357
R20207 VSS.n790 VSS.n688 0.0210357
R20208 VSS.n17916 VSS.n1338 0.0210357
R20209 VSS.n17905 VSS.n1345 0.0210357
R20210 VSS.n17904 VSS.n1347 0.0210357
R20211 VSS.n17187 VSS.n16897 0.0201429
R20212 VSS.n17228 VSS.n16878 0.0201429
R20213 VSS.n17188 VSS.n16899 0.0201429
R20214 VSS.n17779 VSS.n17311 0.0201429
R20215 VSS.n17820 VSS.n17292 0.0201429
R20216 VSS.n17780 VSS.n17313 0.0201429
R20217 VSS.n18500 VSS.n18356 0.0201429
R20218 VSS.n18483 VSS.n18482 0.0201429
R20219 VSS.n18501 VSS.n18354 0.0201429
R20220 VSS.n9829 VSS.n9361 0.0201429
R20221 VSS.n9870 VSS.n9342 0.0201429
R20222 VSS.n9830 VSS.n9363 0.0201429
R20223 VSS.n16772 VSS.n16303 0.0201429
R20224 VSS.n16813 VSS.n16284 0.0201429
R20225 VSS.n16773 VSS.n16305 0.0201429
R20226 VSS.n16179 VSS.n1475 0.0201429
R20227 VSS.n16220 VSS.n1456 0.0201429
R20228 VSS.n16180 VSS.n1477 0.0201429
R20229 VSS.n2147 VSS.n2127 0.0201429
R20230 VSS.n2241 VSS.n2163 0.0201429
R20231 VSS.n2148 VSS.n2129 0.0201429
R20232 VSS.n3320 VSS.n2852 0.0201429
R20233 VSS.n3361 VSS.n2833 0.0201429
R20234 VSS.n3321 VSS.n2854 0.0201429
R20235 VSS.n3912 VSS.n3444 0.0201429
R20236 VSS.n3953 VSS.n3425 0.0201429
R20237 VSS.n3913 VSS.n3446 0.0201429
R20238 VSS.n4504 VSS.n4036 0.0201429
R20239 VSS.n4545 VSS.n4017 0.0201429
R20240 VSS.n4505 VSS.n4038 0.0201429
R20241 VSS.n5096 VSS.n4628 0.0201429
R20242 VSS.n5137 VSS.n4609 0.0201429
R20243 VSS.n5097 VSS.n4630 0.0201429
R20244 VSS.n2743 VSS.n2723 0.0201429
R20245 VSS.n5206 VSS.n2759 0.0201429
R20246 VSS.n2744 VSS.n2725 0.0201429
R20247 VSS.n5704 VSS.n5684 0.0201429
R20248 VSS.n5779 VSS.n5720 0.0201429
R20249 VSS.n5705 VSS.n5686 0.0201429
R20250 VSS.n6277 VSS.n6257 0.0201429
R20251 VSS.n6371 VSS.n6293 0.0201429
R20252 VSS.n6278 VSS.n6259 0.0201429
R20253 VSS.n8053 VSS.n7585 0.0201429
R20254 VSS.n8094 VSS.n7566 0.0201429
R20255 VSS.n8054 VSS.n7587 0.0201429
R20256 VSS.n8645 VSS.n8177 0.0201429
R20257 VSS.n8686 VSS.n8158 0.0201429
R20258 VSS.n8646 VSS.n8179 0.0201429
R20259 VSS.n9237 VSS.n8769 0.0201429
R20260 VSS.n9278 VSS.n8750 0.0201429
R20261 VSS.n9238 VSS.n8771 0.0201429
R20262 VSS.n10421 VSS.n9953 0.0201429
R20263 VSS.n10462 VSS.n9934 0.0201429
R20264 VSS.n10422 VSS.n9955 0.0201429
R20265 VSS.n11013 VSS.n10545 0.0201429
R20266 VSS.n11054 VSS.n10526 0.0201429
R20267 VSS.n11014 VSS.n10547 0.0201429
R20268 VSS.n11605 VSS.n11137 0.0201429
R20269 VSS.n11646 VSS.n11118 0.0201429
R20270 VSS.n11606 VSS.n11139 0.0201429
R20271 VSS.n12197 VSS.n11729 0.0201429
R20272 VSS.n12238 VSS.n11710 0.0201429
R20273 VSS.n12198 VSS.n11731 0.0201429
R20274 VSS.n12789 VSS.n12321 0.0201429
R20275 VSS.n12830 VSS.n12302 0.0201429
R20276 VSS.n12790 VSS.n12323 0.0201429
R20277 VSS.n13381 VSS.n12913 0.0201429
R20278 VSS.n13422 VSS.n12894 0.0201429
R20279 VSS.n13382 VSS.n12915 0.0201429
R20280 VSS.n13973 VSS.n13505 0.0201429
R20281 VSS.n14014 VSS.n13486 0.0201429
R20282 VSS.n13974 VSS.n13507 0.0201429
R20283 VSS.n14565 VSS.n14097 0.0201429
R20284 VSS.n14606 VSS.n14078 0.0201429
R20285 VSS.n14566 VSS.n14099 0.0201429
R20286 VSS.n15157 VSS.n14689 0.0201429
R20287 VSS.n15198 VSS.n14670 0.0201429
R20288 VSS.n15158 VSS.n14691 0.0201429
R20289 VSS.n15749 VSS.n15281 0.0201429
R20290 VSS.n15790 VSS.n15262 0.0201429
R20291 VSS.n15750 VSS.n15283 0.0201429
R20292 VSS.n6883 VSS.n6863 0.0201429
R20293 VSS.n15859 VSS.n6899 0.0201429
R20294 VSS.n6884 VSS.n6865 0.0201429
R20295 VSS.n7461 VSS.n6992 0.0201429
R20296 VSS.n7502 VSS.n6973 0.0201429
R20297 VSS.n7462 VSS.n6994 0.0201429
R20298 VSS.n18773 VSS.n90 0.0201429
R20299 VSS.n18814 VSS.n71 0.0201429
R20300 VSS.n18774 VSS.n92 0.0201429
R20301 VSS.n706 VSS.n686 0.0201429
R20302 VSS.n773 VSS.n722 0.0201429
R20303 VSS.n707 VSS.n688 0.0201429
R20304 VSS.n1365 VSS.n1345 0.0201429
R20305 VSS.n17887 VSS.n1381 0.0201429
R20306 VSS.n1366 VSS.n1347 0.0201429
R20307 VSS.n17154 VSS.n17153 0.01925
R20308 VSS.n17746 VSS.n17745 0.01925
R20309 VSS.n18518 VSS.n18339 0.01925
R20310 VSS.n9796 VSS.n9795 0.01925
R20311 VSS.n16739 VSS.n16738 0.01925
R20312 VSS.n16146 VSS.n16145 0.01925
R20313 VSS.n2115 VSS.n2102 0.01925
R20314 VSS.n3287 VSS.n3286 0.01925
R20315 VSS.n3879 VSS.n3878 0.01925
R20316 VSS.n4471 VSS.n4470 0.01925
R20317 VSS.n5063 VSS.n5062 0.01925
R20318 VSS.n2711 VSS.n2698 0.01925
R20319 VSS.n5672 VSS.n5659 0.01925
R20320 VSS.n6245 VSS.n6232 0.01925
R20321 VSS.n8020 VSS.n8019 0.01925
R20322 VSS.n8612 VSS.n8611 0.01925
R20323 VSS.n9204 VSS.n9203 0.01925
R20324 VSS.n10388 VSS.n10387 0.01925
R20325 VSS.n10980 VSS.n10979 0.01925
R20326 VSS.n11572 VSS.n11571 0.01925
R20327 VSS.n12164 VSS.n12163 0.01925
R20328 VSS.n12756 VSS.n12755 0.01925
R20329 VSS.n13348 VSS.n13347 0.01925
R20330 VSS.n13940 VSS.n13939 0.01925
R20331 VSS.n14532 VSS.n14531 0.01925
R20332 VSS.n15124 VSS.n15123 0.01925
R20333 VSS.n15716 VSS.n15715 0.01925
R20334 VSS.n6851 VSS.n6838 0.01925
R20335 VSS.n7428 VSS.n7427 0.01925
R20336 VSS.n18740 VSS.n18739 0.01925
R20337 VSS.n674 VSS.n661 0.01925
R20338 VSS.n1333 VSS.n1320 0.01925
R20339 VSS.n1179 VSS.n1172 0.0174643
R20340 VSS.n17970 VSS.n1179 0.0174643
R20341 VSS.n17974 VSS.n1175 0.0174643
R20342 VSS.n17971 VSS.n1175 0.0174643
R20343 VSS.n993 VSS.n478 0.0174643
R20344 VSS.n17057 VSS.n17056 0.0174643
R20345 VSS.n17056 VSS.n16963 0.0174643
R20346 VSS.n18019 VSS.n1045 0.0174643
R20347 VSS.n18020 VSS.n1043 0.0174643
R20348 VSS.n17179 VSS.n16902 0.0174643
R20349 VSS.n17058 VSS.n16968 0.0174643
R20350 VSS.n16968 VSS.n16964 0.0174643
R20351 VSS.n17649 VSS.n17648 0.0174643
R20352 VSS.n17648 VSS.n17377 0.0174643
R20353 VSS.n17553 VSS.n17463 0.0174643
R20354 VSS.n17552 VSS.n17551 0.0174643
R20355 VSS.n17771 VSS.n17316 0.0174643
R20356 VSS.n17650 VSS.n17382 0.0174643
R20357 VSS.n17382 VSS.n17378 0.0174643
R20358 VSS.n18130 VSS.n255 0.0174643
R20359 VSS.n18196 VSS.n18189 0.0174643
R20360 VSS.n18559 VSS.n18196 0.0174643
R20361 VSS.n18563 VSS.n18192 0.0174643
R20362 VSS.n18560 VSS.n18192 0.0174643
R20363 VSS.n18353 VSS.n18347 0.0174643
R20364 VSS.n18129 VSS.n18128 0.0174643
R20365 VSS.n9603 VSS.n9513 0.0174643
R20366 VSS.n9699 VSS.n9698 0.0174643
R20367 VSS.n9698 VSS.n9427 0.0174643
R20368 VSS.n9700 VSS.n9432 0.0174643
R20369 VSS.n9432 VSS.n9428 0.0174643
R20370 VSS.n9821 VSS.n9366 0.0174643
R20371 VSS.n9602 VSS.n9601 0.0174643
R20372 VSS.n16452 VSS.n16444 0.0174643
R20373 VSS.n16642 VSS.n16641 0.0174643
R20374 VSS.n16641 VSS.n16369 0.0174643
R20375 VSS.n16643 VSS.n16374 0.0174643
R20376 VSS.n16374 VSS.n16370 0.0174643
R20377 VSS.n16764 VSS.n16308 0.0174643
R20378 VSS.n16451 VSS.n16445 0.0174643
R20379 VSS.n1617 VSS.n1609 0.0174643
R20380 VSS.n16049 VSS.n16048 0.0174643
R20381 VSS.n16048 VSS.n1541 0.0174643
R20382 VSS.n16050 VSS.n1546 0.0174643
R20383 VSS.n1546 VSS.n1542 0.0174643
R20384 VSS.n16171 VSS.n1480 0.0174643
R20385 VSS.n1616 VSS.n1610 0.0174643
R20386 VSS.n1895 VSS.n1805 0.0174643
R20387 VSS.n1961 VSS.n1954 0.0174643
R20388 VSS.n2324 VSS.n1961 0.0174643
R20389 VSS.n2328 VSS.n1957 0.0174643
R20390 VSS.n2325 VSS.n1957 0.0174643
R20391 VSS.n2139 VSS.n2132 0.0174643
R20392 VSS.n1894 VSS.n1893 0.0174643
R20393 VSS.n3094 VSS.n3004 0.0174643
R20394 VSS.n3190 VSS.n3189 0.0174643
R20395 VSS.n3189 VSS.n2918 0.0174643
R20396 VSS.n3191 VSS.n2923 0.0174643
R20397 VSS.n2923 VSS.n2919 0.0174643
R20398 VSS.n3312 VSS.n2857 0.0174643
R20399 VSS.n3093 VSS.n3092 0.0174643
R20400 VSS.n3686 VSS.n3596 0.0174643
R20401 VSS.n3782 VSS.n3781 0.0174643
R20402 VSS.n3781 VSS.n3510 0.0174643
R20403 VSS.n3783 VSS.n3515 0.0174643
R20404 VSS.n3515 VSS.n3511 0.0174643
R20405 VSS.n3904 VSS.n3449 0.0174643
R20406 VSS.n3685 VSS.n3684 0.0174643
R20407 VSS.n4278 VSS.n4188 0.0174643
R20408 VSS.n4374 VSS.n4373 0.0174643
R20409 VSS.n4373 VSS.n4102 0.0174643
R20410 VSS.n4375 VSS.n4107 0.0174643
R20411 VSS.n4107 VSS.n4103 0.0174643
R20412 VSS.n4496 VSS.n4041 0.0174643
R20413 VSS.n4277 VSS.n4276 0.0174643
R20414 VSS.n4870 VSS.n4780 0.0174643
R20415 VSS.n4966 VSS.n4965 0.0174643
R20416 VSS.n4965 VSS.n4694 0.0174643
R20417 VSS.n4967 VSS.n4699 0.0174643
R20418 VSS.n4699 VSS.n4695 0.0174643
R20419 VSS.n5088 VSS.n4633 0.0174643
R20420 VSS.n4869 VSS.n4868 0.0174643
R20421 VSS.n2491 VSS.n2401 0.0174643
R20422 VSS.n2557 VSS.n2550 0.0174643
R20423 VSS.n5289 VSS.n2557 0.0174643
R20424 VSS.n5293 VSS.n2553 0.0174643
R20425 VSS.n5290 VSS.n2553 0.0174643
R20426 VSS.n2735 VSS.n2728 0.0174643
R20427 VSS.n2490 VSS.n2489 0.0174643
R20428 VSS.n5452 VSS.n5362 0.0174643
R20429 VSS.n5518 VSS.n5511 0.0174643
R20430 VSS.n5862 VSS.n5518 0.0174643
R20431 VSS.n5866 VSS.n5514 0.0174643
R20432 VSS.n5863 VSS.n5514 0.0174643
R20433 VSS.n5696 VSS.n5689 0.0174643
R20434 VSS.n5451 VSS.n5450 0.0174643
R20435 VSS.n6025 VSS.n5935 0.0174643
R20436 VSS.n6091 VSS.n6084 0.0174643
R20437 VSS.n6454 VSS.n6091 0.0174643
R20438 VSS.n6458 VSS.n6087 0.0174643
R20439 VSS.n6455 VSS.n6087 0.0174643
R20440 VSS.n6269 VSS.n6262 0.0174643
R20441 VSS.n6024 VSS.n6023 0.0174643
R20442 VSS.n7827 VSS.n7737 0.0174643
R20443 VSS.n7923 VSS.n7922 0.0174643
R20444 VSS.n7922 VSS.n7651 0.0174643
R20445 VSS.n7924 VSS.n7656 0.0174643
R20446 VSS.n7656 VSS.n7652 0.0174643
R20447 VSS.n8045 VSS.n7590 0.0174643
R20448 VSS.n7826 VSS.n7825 0.0174643
R20449 VSS.n8419 VSS.n8329 0.0174643
R20450 VSS.n8515 VSS.n8514 0.0174643
R20451 VSS.n8514 VSS.n8243 0.0174643
R20452 VSS.n8516 VSS.n8248 0.0174643
R20453 VSS.n8248 VSS.n8244 0.0174643
R20454 VSS.n8637 VSS.n8182 0.0174643
R20455 VSS.n8418 VSS.n8417 0.0174643
R20456 VSS.n9011 VSS.n8921 0.0174643
R20457 VSS.n9107 VSS.n9106 0.0174643
R20458 VSS.n9106 VSS.n8835 0.0174643
R20459 VSS.n9108 VSS.n8840 0.0174643
R20460 VSS.n8840 VSS.n8836 0.0174643
R20461 VSS.n9229 VSS.n8774 0.0174643
R20462 VSS.n9010 VSS.n9009 0.0174643
R20463 VSS.n10195 VSS.n10105 0.0174643
R20464 VSS.n10291 VSS.n10290 0.0174643
R20465 VSS.n10290 VSS.n10019 0.0174643
R20466 VSS.n10292 VSS.n10024 0.0174643
R20467 VSS.n10024 VSS.n10020 0.0174643
R20468 VSS.n10413 VSS.n9958 0.0174643
R20469 VSS.n10194 VSS.n10193 0.0174643
R20470 VSS.n10787 VSS.n10697 0.0174643
R20471 VSS.n10883 VSS.n10882 0.0174643
R20472 VSS.n10882 VSS.n10611 0.0174643
R20473 VSS.n10884 VSS.n10616 0.0174643
R20474 VSS.n10616 VSS.n10612 0.0174643
R20475 VSS.n11005 VSS.n10550 0.0174643
R20476 VSS.n10786 VSS.n10785 0.0174643
R20477 VSS.n11379 VSS.n11289 0.0174643
R20478 VSS.n11475 VSS.n11474 0.0174643
R20479 VSS.n11474 VSS.n11203 0.0174643
R20480 VSS.n11476 VSS.n11208 0.0174643
R20481 VSS.n11208 VSS.n11204 0.0174643
R20482 VSS.n11597 VSS.n11142 0.0174643
R20483 VSS.n11378 VSS.n11377 0.0174643
R20484 VSS.n11971 VSS.n11881 0.0174643
R20485 VSS.n12067 VSS.n12066 0.0174643
R20486 VSS.n12066 VSS.n11795 0.0174643
R20487 VSS.n12068 VSS.n11800 0.0174643
R20488 VSS.n11800 VSS.n11796 0.0174643
R20489 VSS.n12189 VSS.n11734 0.0174643
R20490 VSS.n11970 VSS.n11969 0.0174643
R20491 VSS.n12563 VSS.n12473 0.0174643
R20492 VSS.n12659 VSS.n12658 0.0174643
R20493 VSS.n12658 VSS.n12387 0.0174643
R20494 VSS.n12660 VSS.n12392 0.0174643
R20495 VSS.n12392 VSS.n12388 0.0174643
R20496 VSS.n12781 VSS.n12326 0.0174643
R20497 VSS.n12562 VSS.n12561 0.0174643
R20498 VSS.n13155 VSS.n13065 0.0174643
R20499 VSS.n13251 VSS.n13250 0.0174643
R20500 VSS.n13250 VSS.n12979 0.0174643
R20501 VSS.n13252 VSS.n12984 0.0174643
R20502 VSS.n12984 VSS.n12980 0.0174643
R20503 VSS.n13373 VSS.n12918 0.0174643
R20504 VSS.n13154 VSS.n13153 0.0174643
R20505 VSS.n13747 VSS.n13657 0.0174643
R20506 VSS.n13843 VSS.n13842 0.0174643
R20507 VSS.n13842 VSS.n13571 0.0174643
R20508 VSS.n13844 VSS.n13576 0.0174643
R20509 VSS.n13576 VSS.n13572 0.0174643
R20510 VSS.n13965 VSS.n13510 0.0174643
R20511 VSS.n13746 VSS.n13745 0.0174643
R20512 VSS.n14339 VSS.n14249 0.0174643
R20513 VSS.n14435 VSS.n14434 0.0174643
R20514 VSS.n14434 VSS.n14163 0.0174643
R20515 VSS.n14436 VSS.n14168 0.0174643
R20516 VSS.n14168 VSS.n14164 0.0174643
R20517 VSS.n14557 VSS.n14102 0.0174643
R20518 VSS.n14338 VSS.n14337 0.0174643
R20519 VSS.n14931 VSS.n14841 0.0174643
R20520 VSS.n15027 VSS.n15026 0.0174643
R20521 VSS.n15026 VSS.n14755 0.0174643
R20522 VSS.n15028 VSS.n14760 0.0174643
R20523 VSS.n14760 VSS.n14756 0.0174643
R20524 VSS.n15149 VSS.n14694 0.0174643
R20525 VSS.n14930 VSS.n14929 0.0174643
R20526 VSS.n15523 VSS.n15433 0.0174643
R20527 VSS.n15619 VSS.n15618 0.0174643
R20528 VSS.n15618 VSS.n15347 0.0174643
R20529 VSS.n15620 VSS.n15352 0.0174643
R20530 VSS.n15352 VSS.n15348 0.0174643
R20531 VSS.n15741 VSS.n15286 0.0174643
R20532 VSS.n15522 VSS.n15521 0.0174643
R20533 VSS.n6631 VSS.n6541 0.0174643
R20534 VSS.n6697 VSS.n6690 0.0174643
R20535 VSS.n15942 VSS.n6697 0.0174643
R20536 VSS.n15946 VSS.n6693 0.0174643
R20537 VSS.n15943 VSS.n6693 0.0174643
R20538 VSS.n6875 VSS.n6868 0.0174643
R20539 VSS.n6630 VSS.n6629 0.0174643
R20540 VSS.n7141 VSS.n7133 0.0174643
R20541 VSS.n7331 VSS.n7330 0.0174643
R20542 VSS.n7330 VSS.n7058 0.0174643
R20543 VSS.n7332 VSS.n7063 0.0174643
R20544 VSS.n7063 VSS.n7059 0.0174643
R20545 VSS.n7453 VSS.n6997 0.0174643
R20546 VSS.n7140 VSS.n7134 0.0174643
R20547 VSS.n428 VSS.n312 0.0174643
R20548 VSS.n18643 VSS.n18642 0.0174643
R20549 VSS.n18642 VSS.n156 0.0174643
R20550 VSS.n18644 VSS.n161 0.0174643
R20551 VSS.n161 VSS.n157 0.0174643
R20552 VSS.n18765 VSS.n95 0.0174643
R20553 VSS.n429 VSS.n310 0.0174643
R20554 VSS.n517 VSS.n510 0.0174643
R20555 VSS.n856 VSS.n517 0.0174643
R20556 VSS.n860 VSS.n513 0.0174643
R20557 VSS.n857 VSS.n513 0.0174643
R20558 VSS.n698 VSS.n691 0.0174643
R20559 VSS.n994 VSS.n476 0.0174643
R20560 VSS.n1357 VSS.n1350 0.0174643
R20561 VSS.n1231 VSS.n1230 0.0165714
R20562 VSS.n17963 VSS.n17962 0.0165714
R20563 VSS.n1280 VSS.n1278 0.0165714
R20564 VSS.n895 VSS.n470 0.0165714
R20565 VSS.n1076 VSS.n1037 0.0165714
R20566 VSS.n1098 VSS.n1097 0.0165714
R20567 VSS.n18032 VSS.n18031 0.0165714
R20568 VSS.n18031 VSS.n1032 0.0165714
R20569 VSS.n18023 VSS.n1040 0.0165714
R20570 VSS.n1146 VSS.n1144 0.0165714
R20571 VSS.n17189 VSS.n16902 0.0165714
R20572 VSS.n17209 VSS.n16900 0.0165714
R20573 VSS.n17197 VSS.n17193 0.0165714
R20574 VSS.n17014 VSS.n17013 0.0165714
R20575 VSS.n17070 VSS.n16960 0.0165714
R20576 VSS.n17097 VSS.n16943 0.0165714
R20577 VSS.n17554 VSS.n17461 0.0165714
R20578 VSS.n17508 VSS.n17507 0.0165714
R20579 VSS.n17536 VSS.n17471 0.0165714
R20580 VSS.n17536 VSS.n17535 0.0165714
R20581 VSS.n17545 VSS.n17462 0.0165714
R20582 VSS.n17584 VSS.n17583 0.0165714
R20583 VSS.n17781 VSS.n17316 0.0165714
R20584 VSS.n17801 VSS.n17314 0.0165714
R20585 VSS.n17789 VSS.n17785 0.0165714
R20586 VSS.n17606 VSS.n17605 0.0165714
R20587 VSS.n17662 VSS.n17374 0.0165714
R20588 VSS.n17689 VSS.n17357 0.0165714
R20589 VSS.n18131 VSS.n253 0.0165714
R20590 VSS.n18248 VSS.n18247 0.0165714
R20591 VSS.n18552 VSS.n18551 0.0165714
R20592 VSS.n18297 VSS.n18295 0.0165714
R20593 VSS.n18502 VSS.n18353 0.0165714
R20594 VSS.n18399 VSS.n18397 0.0165714
R20595 VSS.n18395 VSS.n18393 0.0165714
R20596 VSS.n18085 VSS.n18084 0.0165714
R20597 VSS.n18113 VSS.n263 0.0165714
R20598 VSS.n18113 VSS.n18112 0.0165714
R20599 VSS.n18122 VSS.n254 0.0165714
R20600 VSS.n18161 VSS.n18160 0.0165714
R20601 VSS.n9604 VSS.n9511 0.0165714
R20602 VSS.n9656 VSS.n9655 0.0165714
R20603 VSS.n9712 VSS.n9424 0.0165714
R20604 VSS.n9739 VSS.n9407 0.0165714
R20605 VSS.n9831 VSS.n9366 0.0165714
R20606 VSS.n9851 VSS.n9364 0.0165714
R20607 VSS.n9839 VSS.n9835 0.0165714
R20608 VSS.n9558 VSS.n9557 0.0165714
R20609 VSS.n9586 VSS.n9521 0.0165714
R20610 VSS.n9586 VSS.n9585 0.0165714
R20611 VSS.n9595 VSS.n9512 0.0165714
R20612 VSS.n9634 VSS.n9633 0.0165714
R20613 VSS.n16537 VSS.n16536 0.0165714
R20614 VSS.n16599 VSS.n16598 0.0165714
R20615 VSS.n16655 VSS.n16366 0.0165714
R20616 VSS.n16682 VSS.n16349 0.0165714
R20617 VSS.n16774 VSS.n16308 0.0165714
R20618 VSS.n16794 VSS.n16306 0.0165714
R20619 VSS.n16782 VSS.n16778 0.0165714
R20620 VSS.n16494 VSS.n16493 0.0165714
R20621 VSS.n16517 VSS.n16466 0.0165714
R20622 VSS.n16517 VSS.n16516 0.0165714
R20623 VSS.n16538 VSS.n16449 0.0165714
R20624 VSS.n16578 VSS.n16424 0.0165714
R20625 VSS.n1702 VSS.n1701 0.0165714
R20626 VSS.n16006 VSS.n16005 0.0165714
R20627 VSS.n16062 VSS.n1538 0.0165714
R20628 VSS.n16089 VSS.n1521 0.0165714
R20629 VSS.n16181 VSS.n1480 0.0165714
R20630 VSS.n16201 VSS.n1478 0.0165714
R20631 VSS.n16189 VSS.n16185 0.0165714
R20632 VSS.n1659 VSS.n1658 0.0165714
R20633 VSS.n1682 VSS.n1631 0.0165714
R20634 VSS.n1682 VSS.n1681 0.0165714
R20635 VSS.n1703 VSS.n1614 0.0165714
R20636 VSS.n1743 VSS.n1589 0.0165714
R20637 VSS.n1896 VSS.n1803 0.0165714
R20638 VSS.n2013 VSS.n2012 0.0165714
R20639 VSS.n2317 VSS.n2316 0.0165714
R20640 VSS.n2062 VSS.n2060 0.0165714
R20641 VSS.n2149 VSS.n2132 0.0165714
R20642 VSS.n2257 VSS.n2130 0.0165714
R20643 VSS.n2182 VSS.n2153 0.0165714
R20644 VSS.n1850 VSS.n1849 0.0165714
R20645 VSS.n1878 VSS.n1813 0.0165714
R20646 VSS.n1878 VSS.n1877 0.0165714
R20647 VSS.n1887 VSS.n1804 0.0165714
R20648 VSS.n1926 VSS.n1925 0.0165714
R20649 VSS.n3095 VSS.n3002 0.0165714
R20650 VSS.n3147 VSS.n3146 0.0165714
R20651 VSS.n3203 VSS.n2915 0.0165714
R20652 VSS.n3230 VSS.n2898 0.0165714
R20653 VSS.n3322 VSS.n2857 0.0165714
R20654 VSS.n3342 VSS.n2855 0.0165714
R20655 VSS.n3330 VSS.n3326 0.0165714
R20656 VSS.n3049 VSS.n3048 0.0165714
R20657 VSS.n3077 VSS.n3012 0.0165714
R20658 VSS.n3077 VSS.n3076 0.0165714
R20659 VSS.n3086 VSS.n3003 0.0165714
R20660 VSS.n3125 VSS.n3124 0.0165714
R20661 VSS.n3687 VSS.n3594 0.0165714
R20662 VSS.n3739 VSS.n3738 0.0165714
R20663 VSS.n3795 VSS.n3507 0.0165714
R20664 VSS.n3822 VSS.n3490 0.0165714
R20665 VSS.n3914 VSS.n3449 0.0165714
R20666 VSS.n3934 VSS.n3447 0.0165714
R20667 VSS.n3922 VSS.n3918 0.0165714
R20668 VSS.n3641 VSS.n3640 0.0165714
R20669 VSS.n3669 VSS.n3604 0.0165714
R20670 VSS.n3669 VSS.n3668 0.0165714
R20671 VSS.n3678 VSS.n3595 0.0165714
R20672 VSS.n3717 VSS.n3716 0.0165714
R20673 VSS.n4279 VSS.n4186 0.0165714
R20674 VSS.n4331 VSS.n4330 0.0165714
R20675 VSS.n4387 VSS.n4099 0.0165714
R20676 VSS.n4414 VSS.n4082 0.0165714
R20677 VSS.n4506 VSS.n4041 0.0165714
R20678 VSS.n4526 VSS.n4039 0.0165714
R20679 VSS.n4514 VSS.n4510 0.0165714
R20680 VSS.n4233 VSS.n4232 0.0165714
R20681 VSS.n4261 VSS.n4196 0.0165714
R20682 VSS.n4261 VSS.n4260 0.0165714
R20683 VSS.n4270 VSS.n4187 0.0165714
R20684 VSS.n4309 VSS.n4308 0.0165714
R20685 VSS.n4871 VSS.n4778 0.0165714
R20686 VSS.n4923 VSS.n4922 0.0165714
R20687 VSS.n4979 VSS.n4691 0.0165714
R20688 VSS.n5006 VSS.n4674 0.0165714
R20689 VSS.n5098 VSS.n4633 0.0165714
R20690 VSS.n5118 VSS.n4631 0.0165714
R20691 VSS.n5106 VSS.n5102 0.0165714
R20692 VSS.n4825 VSS.n4824 0.0165714
R20693 VSS.n4853 VSS.n4788 0.0165714
R20694 VSS.n4853 VSS.n4852 0.0165714
R20695 VSS.n4862 VSS.n4779 0.0165714
R20696 VSS.n4901 VSS.n4900 0.0165714
R20697 VSS.n2492 VSS.n2399 0.0165714
R20698 VSS.n2609 VSS.n2608 0.0165714
R20699 VSS.n5282 VSS.n5281 0.0165714
R20700 VSS.n2658 VSS.n2656 0.0165714
R20701 VSS.n2745 VSS.n2728 0.0165714
R20702 VSS.n5222 VSS.n2726 0.0165714
R20703 VSS.n2778 VSS.n2749 0.0165714
R20704 VSS.n2446 VSS.n2445 0.0165714
R20705 VSS.n2474 VSS.n2409 0.0165714
R20706 VSS.n2474 VSS.n2473 0.0165714
R20707 VSS.n2483 VSS.n2400 0.0165714
R20708 VSS.n2522 VSS.n2521 0.0165714
R20709 VSS.n5453 VSS.n5360 0.0165714
R20710 VSS.n5570 VSS.n5569 0.0165714
R20711 VSS.n5855 VSS.n5854 0.0165714
R20712 VSS.n5619 VSS.n5617 0.0165714
R20713 VSS.n5706 VSS.n5689 0.0165714
R20714 VSS.n5795 VSS.n5687 0.0165714
R20715 VSS.n5752 VSS.n5710 0.0165714
R20716 VSS.n5407 VSS.n5406 0.0165714
R20717 VSS.n5435 VSS.n5370 0.0165714
R20718 VSS.n5435 VSS.n5434 0.0165714
R20719 VSS.n5444 VSS.n5361 0.0165714
R20720 VSS.n5483 VSS.n5482 0.0165714
R20721 VSS.n6026 VSS.n5933 0.0165714
R20722 VSS.n6143 VSS.n6142 0.0165714
R20723 VSS.n6447 VSS.n6446 0.0165714
R20724 VSS.n6192 VSS.n6190 0.0165714
R20725 VSS.n6279 VSS.n6262 0.0165714
R20726 VSS.n6387 VSS.n6260 0.0165714
R20727 VSS.n6312 VSS.n6283 0.0165714
R20728 VSS.n5980 VSS.n5979 0.0165714
R20729 VSS.n6008 VSS.n5943 0.0165714
R20730 VSS.n6008 VSS.n6007 0.0165714
R20731 VSS.n6017 VSS.n5934 0.0165714
R20732 VSS.n6056 VSS.n6055 0.0165714
R20733 VSS.n7828 VSS.n7735 0.0165714
R20734 VSS.n7880 VSS.n7879 0.0165714
R20735 VSS.n7936 VSS.n7648 0.0165714
R20736 VSS.n7963 VSS.n7631 0.0165714
R20737 VSS.n8055 VSS.n7590 0.0165714
R20738 VSS.n8075 VSS.n7588 0.0165714
R20739 VSS.n8063 VSS.n8059 0.0165714
R20740 VSS.n7782 VSS.n7781 0.0165714
R20741 VSS.n7810 VSS.n7745 0.0165714
R20742 VSS.n7810 VSS.n7809 0.0165714
R20743 VSS.n7819 VSS.n7736 0.0165714
R20744 VSS.n7858 VSS.n7857 0.0165714
R20745 VSS.n8420 VSS.n8327 0.0165714
R20746 VSS.n8472 VSS.n8471 0.0165714
R20747 VSS.n8528 VSS.n8240 0.0165714
R20748 VSS.n8555 VSS.n8223 0.0165714
R20749 VSS.n8647 VSS.n8182 0.0165714
R20750 VSS.n8667 VSS.n8180 0.0165714
R20751 VSS.n8655 VSS.n8651 0.0165714
R20752 VSS.n8374 VSS.n8373 0.0165714
R20753 VSS.n8402 VSS.n8337 0.0165714
R20754 VSS.n8402 VSS.n8401 0.0165714
R20755 VSS.n8411 VSS.n8328 0.0165714
R20756 VSS.n8450 VSS.n8449 0.0165714
R20757 VSS.n9012 VSS.n8919 0.0165714
R20758 VSS.n9064 VSS.n9063 0.0165714
R20759 VSS.n9120 VSS.n8832 0.0165714
R20760 VSS.n9147 VSS.n8815 0.0165714
R20761 VSS.n9239 VSS.n8774 0.0165714
R20762 VSS.n9259 VSS.n8772 0.0165714
R20763 VSS.n9247 VSS.n9243 0.0165714
R20764 VSS.n8966 VSS.n8965 0.0165714
R20765 VSS.n8994 VSS.n8929 0.0165714
R20766 VSS.n8994 VSS.n8993 0.0165714
R20767 VSS.n9003 VSS.n8920 0.0165714
R20768 VSS.n9042 VSS.n9041 0.0165714
R20769 VSS.n10196 VSS.n10103 0.0165714
R20770 VSS.n10248 VSS.n10247 0.0165714
R20771 VSS.n10304 VSS.n10016 0.0165714
R20772 VSS.n10331 VSS.n9999 0.0165714
R20773 VSS.n10423 VSS.n9958 0.0165714
R20774 VSS.n10443 VSS.n9956 0.0165714
R20775 VSS.n10431 VSS.n10427 0.0165714
R20776 VSS.n10150 VSS.n10149 0.0165714
R20777 VSS.n10178 VSS.n10113 0.0165714
R20778 VSS.n10178 VSS.n10177 0.0165714
R20779 VSS.n10187 VSS.n10104 0.0165714
R20780 VSS.n10226 VSS.n10225 0.0165714
R20781 VSS.n10788 VSS.n10695 0.0165714
R20782 VSS.n10840 VSS.n10839 0.0165714
R20783 VSS.n10896 VSS.n10608 0.0165714
R20784 VSS.n10923 VSS.n10591 0.0165714
R20785 VSS.n11015 VSS.n10550 0.0165714
R20786 VSS.n11035 VSS.n10548 0.0165714
R20787 VSS.n11023 VSS.n11019 0.0165714
R20788 VSS.n10742 VSS.n10741 0.0165714
R20789 VSS.n10770 VSS.n10705 0.0165714
R20790 VSS.n10770 VSS.n10769 0.0165714
R20791 VSS.n10779 VSS.n10696 0.0165714
R20792 VSS.n10818 VSS.n10817 0.0165714
R20793 VSS.n11380 VSS.n11287 0.0165714
R20794 VSS.n11432 VSS.n11431 0.0165714
R20795 VSS.n11488 VSS.n11200 0.0165714
R20796 VSS.n11515 VSS.n11183 0.0165714
R20797 VSS.n11607 VSS.n11142 0.0165714
R20798 VSS.n11627 VSS.n11140 0.0165714
R20799 VSS.n11615 VSS.n11611 0.0165714
R20800 VSS.n11334 VSS.n11333 0.0165714
R20801 VSS.n11362 VSS.n11297 0.0165714
R20802 VSS.n11362 VSS.n11361 0.0165714
R20803 VSS.n11371 VSS.n11288 0.0165714
R20804 VSS.n11410 VSS.n11409 0.0165714
R20805 VSS.n11972 VSS.n11879 0.0165714
R20806 VSS.n12024 VSS.n12023 0.0165714
R20807 VSS.n12080 VSS.n11792 0.0165714
R20808 VSS.n12107 VSS.n11775 0.0165714
R20809 VSS.n12199 VSS.n11734 0.0165714
R20810 VSS.n12219 VSS.n11732 0.0165714
R20811 VSS.n12207 VSS.n12203 0.0165714
R20812 VSS.n11926 VSS.n11925 0.0165714
R20813 VSS.n11954 VSS.n11889 0.0165714
R20814 VSS.n11954 VSS.n11953 0.0165714
R20815 VSS.n11963 VSS.n11880 0.0165714
R20816 VSS.n12002 VSS.n12001 0.0165714
R20817 VSS.n12564 VSS.n12471 0.0165714
R20818 VSS.n12616 VSS.n12615 0.0165714
R20819 VSS.n12672 VSS.n12384 0.0165714
R20820 VSS.n12699 VSS.n12367 0.0165714
R20821 VSS.n12791 VSS.n12326 0.0165714
R20822 VSS.n12811 VSS.n12324 0.0165714
R20823 VSS.n12799 VSS.n12795 0.0165714
R20824 VSS.n12518 VSS.n12517 0.0165714
R20825 VSS.n12546 VSS.n12481 0.0165714
R20826 VSS.n12546 VSS.n12545 0.0165714
R20827 VSS.n12555 VSS.n12472 0.0165714
R20828 VSS.n12594 VSS.n12593 0.0165714
R20829 VSS.n13156 VSS.n13063 0.0165714
R20830 VSS.n13208 VSS.n13207 0.0165714
R20831 VSS.n13264 VSS.n12976 0.0165714
R20832 VSS.n13291 VSS.n12959 0.0165714
R20833 VSS.n13383 VSS.n12918 0.0165714
R20834 VSS.n13403 VSS.n12916 0.0165714
R20835 VSS.n13391 VSS.n13387 0.0165714
R20836 VSS.n13110 VSS.n13109 0.0165714
R20837 VSS.n13138 VSS.n13073 0.0165714
R20838 VSS.n13138 VSS.n13137 0.0165714
R20839 VSS.n13147 VSS.n13064 0.0165714
R20840 VSS.n13186 VSS.n13185 0.0165714
R20841 VSS.n13748 VSS.n13655 0.0165714
R20842 VSS.n13800 VSS.n13799 0.0165714
R20843 VSS.n13856 VSS.n13568 0.0165714
R20844 VSS.n13883 VSS.n13551 0.0165714
R20845 VSS.n13975 VSS.n13510 0.0165714
R20846 VSS.n13995 VSS.n13508 0.0165714
R20847 VSS.n13983 VSS.n13979 0.0165714
R20848 VSS.n13702 VSS.n13701 0.0165714
R20849 VSS.n13730 VSS.n13665 0.0165714
R20850 VSS.n13730 VSS.n13729 0.0165714
R20851 VSS.n13739 VSS.n13656 0.0165714
R20852 VSS.n13778 VSS.n13777 0.0165714
R20853 VSS.n14340 VSS.n14247 0.0165714
R20854 VSS.n14392 VSS.n14391 0.0165714
R20855 VSS.n14448 VSS.n14160 0.0165714
R20856 VSS.n14475 VSS.n14143 0.0165714
R20857 VSS.n14567 VSS.n14102 0.0165714
R20858 VSS.n14587 VSS.n14100 0.0165714
R20859 VSS.n14575 VSS.n14571 0.0165714
R20860 VSS.n14294 VSS.n14293 0.0165714
R20861 VSS.n14322 VSS.n14257 0.0165714
R20862 VSS.n14322 VSS.n14321 0.0165714
R20863 VSS.n14331 VSS.n14248 0.0165714
R20864 VSS.n14370 VSS.n14369 0.0165714
R20865 VSS.n14932 VSS.n14839 0.0165714
R20866 VSS.n14984 VSS.n14983 0.0165714
R20867 VSS.n15040 VSS.n14752 0.0165714
R20868 VSS.n15067 VSS.n14735 0.0165714
R20869 VSS.n15159 VSS.n14694 0.0165714
R20870 VSS.n15179 VSS.n14692 0.0165714
R20871 VSS.n15167 VSS.n15163 0.0165714
R20872 VSS.n14886 VSS.n14885 0.0165714
R20873 VSS.n14914 VSS.n14849 0.0165714
R20874 VSS.n14914 VSS.n14913 0.0165714
R20875 VSS.n14923 VSS.n14840 0.0165714
R20876 VSS.n14962 VSS.n14961 0.0165714
R20877 VSS.n15524 VSS.n15431 0.0165714
R20878 VSS.n15576 VSS.n15575 0.0165714
R20879 VSS.n15632 VSS.n15344 0.0165714
R20880 VSS.n15659 VSS.n15327 0.0165714
R20881 VSS.n15751 VSS.n15286 0.0165714
R20882 VSS.n15771 VSS.n15284 0.0165714
R20883 VSS.n15759 VSS.n15755 0.0165714
R20884 VSS.n15478 VSS.n15477 0.0165714
R20885 VSS.n15506 VSS.n15441 0.0165714
R20886 VSS.n15506 VSS.n15505 0.0165714
R20887 VSS.n15515 VSS.n15432 0.0165714
R20888 VSS.n15554 VSS.n15553 0.0165714
R20889 VSS.n6632 VSS.n6539 0.0165714
R20890 VSS.n6749 VSS.n6748 0.0165714
R20891 VSS.n15935 VSS.n15934 0.0165714
R20892 VSS.n6798 VSS.n6796 0.0165714
R20893 VSS.n6885 VSS.n6868 0.0165714
R20894 VSS.n15875 VSS.n6866 0.0165714
R20895 VSS.n6918 VSS.n6889 0.0165714
R20896 VSS.n6586 VSS.n6585 0.0165714
R20897 VSS.n6614 VSS.n6549 0.0165714
R20898 VSS.n6614 VSS.n6613 0.0165714
R20899 VSS.n6623 VSS.n6540 0.0165714
R20900 VSS.n6662 VSS.n6661 0.0165714
R20901 VSS.n7226 VSS.n7225 0.0165714
R20902 VSS.n7288 VSS.n7287 0.0165714
R20903 VSS.n7344 VSS.n7055 0.0165714
R20904 VSS.n7371 VSS.n7038 0.0165714
R20905 VSS.n7463 VSS.n6997 0.0165714
R20906 VSS.n7483 VSS.n6995 0.0165714
R20907 VSS.n7471 VSS.n7467 0.0165714
R20908 VSS.n7183 VSS.n7182 0.0165714
R20909 VSS.n7206 VSS.n7155 0.0165714
R20910 VSS.n7206 VSS.n7205 0.0165714
R20911 VSS.n7227 VSS.n7138 0.0165714
R20912 VSS.n7267 VSS.n7113 0.0165714
R20913 VSS.n378 VSS.n304 0.0165714
R20914 VSS.n18600 VSS.n18599 0.0165714
R20915 VSS.n18656 VSS.n153 0.0165714
R20916 VSS.n18683 VSS.n136 0.0165714
R20917 VSS.n18775 VSS.n95 0.0165714
R20918 VSS.n18795 VSS.n93 0.0165714
R20919 VSS.n18783 VSS.n18779 0.0165714
R20920 VSS.n353 VSS.n351 0.0165714
R20921 VSS.n441 VSS.n440 0.0165714
R20922 VSS.n440 VSS.n299 0.0165714
R20923 VSS.n432 VSS.n307 0.0165714
R20924 VSS.n409 VSS.n408 0.0165714
R20925 VSS.n572 VSS.n571 0.0165714
R20926 VSS.n849 VSS.n848 0.0165714
R20927 VSS.n621 VSS.n619 0.0165714
R20928 VSS.n708 VSS.n691 0.0165714
R20929 VSS.n789 VSS.n689 0.0165714
R20930 VSS.n750 VSS.n712 0.0165714
R20931 VSS.n917 VSS.n916 0.0165714
R20932 VSS.n1006 VSS.n1005 0.0165714
R20933 VSS.n1005 VSS.n465 0.0165714
R20934 VSS.n997 VSS.n473 0.0165714
R20935 VSS.n965 VSS.n963 0.0165714
R20936 VSS.n1367 VSS.n1350 0.0165714
R20937 VSS.n17903 VSS.n1348 0.0165714
R20938 VSS.n1400 VSS.n1371 0.0165714
R20939 VSS.n17983 VSS.n17982 0.0156786
R20940 VSS.n18012 VSS.n18011 0.0156786
R20941 VSS.n17142 VSS.n17138 0.0156786
R20942 VSS.n17147 VSS.n16926 0.0156786
R20943 VSS.n16926 VSS.n16920 0.0156786
R20944 VSS.n17229 VSS.n16876 0.0156786
R20945 VSS.n17244 VSS.n16876 0.0156786
R20946 VSS.n17037 VSS.n16983 0.0156786
R20947 VSS.n17572 VSS.n17571 0.0156786
R20948 VSS.n17734 VSS.n17730 0.0156786
R20949 VSS.n17739 VSS.n17340 0.0156786
R20950 VSS.n17340 VSS.n17334 0.0156786
R20951 VSS.n17821 VSS.n17290 0.0156786
R20952 VSS.n17836 VSS.n17290 0.0156786
R20953 VSS.n17629 VSS.n17397 0.0156786
R20954 VSS.n18572 VSS.n18571 0.0156786
R20955 VSS.n18334 VSS.n18332 0.0156786
R20956 VSS.n18523 VSS.n18317 0.0156786
R20957 VSS.n18519 VSS.n18317 0.0156786
R20958 VSS.n18484 VSS.n18417 0.0156786
R20959 VSS.n18424 VSS.n18417 0.0156786
R20960 VSS.n18149 VSS.n18148 0.0156786
R20961 VSS.n9679 VSS.n9447 0.0156786
R20962 VSS.n9784 VSS.n9780 0.0156786
R20963 VSS.n9789 VSS.n9390 0.0156786
R20964 VSS.n9390 VSS.n9384 0.0156786
R20965 VSS.n9871 VSS.n9341 0.0156786
R20966 VSS.n9886 VSS.n9341 0.0156786
R20967 VSS.n9622 VSS.n9621 0.0156786
R20968 VSS.n16622 VSS.n16389 0.0156786
R20969 VSS.n16727 VSS.n16723 0.0156786
R20970 VSS.n16732 VSS.n16332 0.0156786
R20971 VSS.n16332 VSS.n16326 0.0156786
R20972 VSS.n16814 VSS.n16283 0.0156786
R20973 VSS.n16829 VSS.n16283 0.0156786
R20974 VSS.n16550 VSS.n16441 0.0156786
R20975 VSS.n16029 VSS.n1561 0.0156786
R20976 VSS.n16134 VSS.n16130 0.0156786
R20977 VSS.n16139 VSS.n1504 0.0156786
R20978 VSS.n1504 VSS.n1498 0.0156786
R20979 VSS.n16221 VSS.n1455 0.0156786
R20980 VSS.n16236 VSS.n1455 0.0156786
R20981 VSS.n1715 VSS.n1606 0.0156786
R20982 VSS.n2337 VSS.n2336 0.0156786
R20983 VSS.n2098 VSS.n2096 0.0156786
R20984 VSS.n2288 VSS.n2082 0.0156786
R20985 VSS.n2116 VSS.n2082 0.0156786
R20986 VSS.n2240 VSS.n2164 0.0156786
R20987 VSS.n2236 VSS.n2164 0.0156786
R20988 VSS.n1914 VSS.n1913 0.0156786
R20989 VSS.n3170 VSS.n2938 0.0156786
R20990 VSS.n3275 VSS.n3271 0.0156786
R20991 VSS.n3280 VSS.n2881 0.0156786
R20992 VSS.n2881 VSS.n2875 0.0156786
R20993 VSS.n3362 VSS.n2832 0.0156786
R20994 VSS.n3377 VSS.n2832 0.0156786
R20995 VSS.n3113 VSS.n3112 0.0156786
R20996 VSS.n3762 VSS.n3530 0.0156786
R20997 VSS.n3867 VSS.n3863 0.0156786
R20998 VSS.n3872 VSS.n3473 0.0156786
R20999 VSS.n3473 VSS.n3467 0.0156786
R21000 VSS.n3954 VSS.n3424 0.0156786
R21001 VSS.n3969 VSS.n3424 0.0156786
R21002 VSS.n3705 VSS.n3704 0.0156786
R21003 VSS.n4354 VSS.n4122 0.0156786
R21004 VSS.n4459 VSS.n4455 0.0156786
R21005 VSS.n4464 VSS.n4065 0.0156786
R21006 VSS.n4065 VSS.n4059 0.0156786
R21007 VSS.n4546 VSS.n4016 0.0156786
R21008 VSS.n4561 VSS.n4016 0.0156786
R21009 VSS.n4297 VSS.n4296 0.0156786
R21010 VSS.n4946 VSS.n4714 0.0156786
R21011 VSS.n5051 VSS.n5047 0.0156786
R21012 VSS.n5056 VSS.n4657 0.0156786
R21013 VSS.n4657 VSS.n4651 0.0156786
R21014 VSS.n5138 VSS.n4608 0.0156786
R21015 VSS.n5153 VSS.n4608 0.0156786
R21016 VSS.n4889 VSS.n4888 0.0156786
R21017 VSS.n5302 VSS.n5301 0.0156786
R21018 VSS.n2694 VSS.n2692 0.0156786
R21019 VSS.n5253 VSS.n2678 0.0156786
R21020 VSS.n2712 VSS.n2678 0.0156786
R21021 VSS.n5205 VSS.n2760 0.0156786
R21022 VSS.n5201 VSS.n2760 0.0156786
R21023 VSS.n2510 VSS.n2509 0.0156786
R21024 VSS.n5875 VSS.n5874 0.0156786
R21025 VSS.n5655 VSS.n5653 0.0156786
R21026 VSS.n5826 VSS.n5639 0.0156786
R21027 VSS.n5673 VSS.n5639 0.0156786
R21028 VSS.n5778 VSS.n5721 0.0156786
R21029 VSS.n5774 VSS.n5721 0.0156786
R21030 VSS.n5471 VSS.n5470 0.0156786
R21031 VSS.n6467 VSS.n6466 0.0156786
R21032 VSS.n6228 VSS.n6226 0.0156786
R21033 VSS.n6418 VSS.n6212 0.0156786
R21034 VSS.n6246 VSS.n6212 0.0156786
R21035 VSS.n6370 VSS.n6294 0.0156786
R21036 VSS.n6366 VSS.n6294 0.0156786
R21037 VSS.n6044 VSS.n6043 0.0156786
R21038 VSS.n7903 VSS.n7671 0.0156786
R21039 VSS.n8008 VSS.n8004 0.0156786
R21040 VSS.n8013 VSS.n7614 0.0156786
R21041 VSS.n7614 VSS.n7608 0.0156786
R21042 VSS.n8095 VSS.n7565 0.0156786
R21043 VSS.n8110 VSS.n7565 0.0156786
R21044 VSS.n7846 VSS.n7845 0.0156786
R21045 VSS.n8495 VSS.n8263 0.0156786
R21046 VSS.n8600 VSS.n8596 0.0156786
R21047 VSS.n8605 VSS.n8206 0.0156786
R21048 VSS.n8206 VSS.n8200 0.0156786
R21049 VSS.n8687 VSS.n8157 0.0156786
R21050 VSS.n8702 VSS.n8157 0.0156786
R21051 VSS.n8438 VSS.n8437 0.0156786
R21052 VSS.n9087 VSS.n8855 0.0156786
R21053 VSS.n9192 VSS.n9188 0.0156786
R21054 VSS.n9197 VSS.n8798 0.0156786
R21055 VSS.n8798 VSS.n8792 0.0156786
R21056 VSS.n9279 VSS.n8749 0.0156786
R21057 VSS.n9294 VSS.n8749 0.0156786
R21058 VSS.n9030 VSS.n9029 0.0156786
R21059 VSS.n10271 VSS.n10039 0.0156786
R21060 VSS.n10376 VSS.n10372 0.0156786
R21061 VSS.n10381 VSS.n9982 0.0156786
R21062 VSS.n9982 VSS.n9976 0.0156786
R21063 VSS.n10463 VSS.n9933 0.0156786
R21064 VSS.n10478 VSS.n9933 0.0156786
R21065 VSS.n10214 VSS.n10213 0.0156786
R21066 VSS.n10863 VSS.n10631 0.0156786
R21067 VSS.n10968 VSS.n10964 0.0156786
R21068 VSS.n10973 VSS.n10574 0.0156786
R21069 VSS.n10574 VSS.n10568 0.0156786
R21070 VSS.n11055 VSS.n10525 0.0156786
R21071 VSS.n11070 VSS.n10525 0.0156786
R21072 VSS.n10806 VSS.n10805 0.0156786
R21073 VSS.n11455 VSS.n11223 0.0156786
R21074 VSS.n11560 VSS.n11556 0.0156786
R21075 VSS.n11565 VSS.n11166 0.0156786
R21076 VSS.n11166 VSS.n11160 0.0156786
R21077 VSS.n11647 VSS.n11117 0.0156786
R21078 VSS.n11662 VSS.n11117 0.0156786
R21079 VSS.n11398 VSS.n11397 0.0156786
R21080 VSS.n12047 VSS.n11815 0.0156786
R21081 VSS.n12152 VSS.n12148 0.0156786
R21082 VSS.n12157 VSS.n11758 0.0156786
R21083 VSS.n11758 VSS.n11752 0.0156786
R21084 VSS.n12239 VSS.n11709 0.0156786
R21085 VSS.n12254 VSS.n11709 0.0156786
R21086 VSS.n11990 VSS.n11989 0.0156786
R21087 VSS.n12639 VSS.n12407 0.0156786
R21088 VSS.n12744 VSS.n12740 0.0156786
R21089 VSS.n12749 VSS.n12350 0.0156786
R21090 VSS.n12350 VSS.n12344 0.0156786
R21091 VSS.n12831 VSS.n12301 0.0156786
R21092 VSS.n12846 VSS.n12301 0.0156786
R21093 VSS.n12582 VSS.n12581 0.0156786
R21094 VSS.n13231 VSS.n12999 0.0156786
R21095 VSS.n13336 VSS.n13332 0.0156786
R21096 VSS.n13341 VSS.n12942 0.0156786
R21097 VSS.n12942 VSS.n12936 0.0156786
R21098 VSS.n13423 VSS.n12893 0.0156786
R21099 VSS.n13438 VSS.n12893 0.0156786
R21100 VSS.n13174 VSS.n13173 0.0156786
R21101 VSS.n13823 VSS.n13591 0.0156786
R21102 VSS.n13928 VSS.n13924 0.0156786
R21103 VSS.n13933 VSS.n13534 0.0156786
R21104 VSS.n13534 VSS.n13528 0.0156786
R21105 VSS.n14015 VSS.n13485 0.0156786
R21106 VSS.n14030 VSS.n13485 0.0156786
R21107 VSS.n13766 VSS.n13765 0.0156786
R21108 VSS.n14415 VSS.n14183 0.0156786
R21109 VSS.n14520 VSS.n14516 0.0156786
R21110 VSS.n14525 VSS.n14126 0.0156786
R21111 VSS.n14126 VSS.n14120 0.0156786
R21112 VSS.n14607 VSS.n14077 0.0156786
R21113 VSS.n14622 VSS.n14077 0.0156786
R21114 VSS.n14358 VSS.n14357 0.0156786
R21115 VSS.n15007 VSS.n14775 0.0156786
R21116 VSS.n15112 VSS.n15108 0.0156786
R21117 VSS.n15117 VSS.n14718 0.0156786
R21118 VSS.n14718 VSS.n14712 0.0156786
R21119 VSS.n15199 VSS.n14669 0.0156786
R21120 VSS.n15214 VSS.n14669 0.0156786
R21121 VSS.n14950 VSS.n14949 0.0156786
R21122 VSS.n15599 VSS.n15367 0.0156786
R21123 VSS.n15704 VSS.n15700 0.0156786
R21124 VSS.n15709 VSS.n15310 0.0156786
R21125 VSS.n15310 VSS.n15304 0.0156786
R21126 VSS.n15791 VSS.n15261 0.0156786
R21127 VSS.n15806 VSS.n15261 0.0156786
R21128 VSS.n15542 VSS.n15541 0.0156786
R21129 VSS.n15955 VSS.n15954 0.0156786
R21130 VSS.n6834 VSS.n6832 0.0156786
R21131 VSS.n15906 VSS.n6818 0.0156786
R21132 VSS.n6852 VSS.n6818 0.0156786
R21133 VSS.n15858 VSS.n6900 0.0156786
R21134 VSS.n15854 VSS.n6900 0.0156786
R21135 VSS.n6650 VSS.n6649 0.0156786
R21136 VSS.n7311 VSS.n7078 0.0156786
R21137 VSS.n7416 VSS.n7412 0.0156786
R21138 VSS.n7421 VSS.n7021 0.0156786
R21139 VSS.n7021 VSS.n7015 0.0156786
R21140 VSS.n7503 VSS.n6972 0.0156786
R21141 VSS.n7518 VSS.n6972 0.0156786
R21142 VSS.n7239 VSS.n7130 0.0156786
R21143 VSS.n18623 VSS.n176 0.0156786
R21144 VSS.n18728 VSS.n18724 0.0156786
R21145 VSS.n18733 VSS.n119 0.0156786
R21146 VSS.n119 VSS.n113 0.0156786
R21147 VSS.n18815 VSS.n70 0.0156786
R21148 VSS.n18830 VSS.n70 0.0156786
R21149 VSS.n421 VSS.n420 0.0156786
R21150 VSS.n869 VSS.n868 0.0156786
R21151 VSS.n657 VSS.n655 0.0156786
R21152 VSS.n820 VSS.n641 0.0156786
R21153 VSS.n675 VSS.n641 0.0156786
R21154 VSS.n772 VSS.n723 0.0156786
R21155 VSS.n768 VSS.n723 0.0156786
R21156 VSS.n986 VSS.n985 0.0156786
R21157 VSS.n1316 VSS.n1314 0.0156786
R21158 VSS.n17934 VSS.n1300 0.0156786
R21159 VSS.n1334 VSS.n1300 0.0156786
R21160 VSS.n17886 VSS.n1382 0.0156786
R21161 VSS.n17882 VSS.n1382 0.0156786
R21162 VSS.n18030 VSS.n18029 0.0152714
R21163 VSS.n18014 VSS.n18013 0.0152714
R21164 VSS.n17042 VSS.n17038 0.0152714
R21165 VSS.n17069 VSS.n17068 0.0152714
R21166 VSS.n17190 VSS.n16901 0.0152714
R21167 VSS.n17208 VSS.n17207 0.0152714
R21168 VSS.n17538 VSS.n17537 0.0152714
R21169 VSS.n17570 VSS.n17569 0.0152714
R21170 VSS.n17634 VSS.n17630 0.0152714
R21171 VSS.n17661 VSS.n17660 0.0152714
R21172 VSS.n17782 VSS.n17315 0.0152714
R21173 VSS.n17800 VSS.n17799 0.0152714
R21174 VSS.n18115 VSS.n18114 0.0152714
R21175 VSS.n18147 VSS.n18146 0.0152714
R21176 VSS.n18570 VSS.n18569 0.0152714
R21177 VSS.n18554 VSS.n18553 0.0152714
R21178 VSS.n18504 VSS.n18503 0.0152714
R21179 VSS.n18398 VSS.n18392 0.0152714
R21180 VSS.n9684 VSS.n9680 0.0152714
R21181 VSS.n9711 VSS.n9710 0.0152714
R21182 VSS.n9832 VSS.n9365 0.0152714
R21183 VSS.n9850 VSS.n9849 0.0152714
R21184 VSS.n16522 VSS.n16518 0.0152714
R21185 VSS.n16549 VSS.n16548 0.0152714
R21186 VSS.n16627 VSS.n16623 0.0152714
R21187 VSS.n16654 VSS.n16653 0.0152714
R21188 VSS.n16775 VSS.n16307 0.0152714
R21189 VSS.n16793 VSS.n16792 0.0152714
R21190 VSS.n1687 VSS.n1683 0.0152714
R21191 VSS.n1714 VSS.n1713 0.0152714
R21192 VSS.n16034 VSS.n16030 0.0152714
R21193 VSS.n16061 VSS.n16060 0.0152714
R21194 VSS.n16182 VSS.n1479 0.0152714
R21195 VSS.n16200 VSS.n16199 0.0152714
R21196 VSS.n1880 VSS.n1879 0.0152714
R21197 VSS.n1912 VSS.n1911 0.0152714
R21198 VSS.n2335 VSS.n2334 0.0152714
R21199 VSS.n2319 VSS.n2318 0.0152714
R21200 VSS.n2150 VSS.n2131 0.0152714
R21201 VSS.n2256 VSS.n2255 0.0152714
R21202 VSS.n3079 VSS.n3078 0.0152714
R21203 VSS.n3111 VSS.n3110 0.0152714
R21204 VSS.n3175 VSS.n3171 0.0152714
R21205 VSS.n3202 VSS.n3201 0.0152714
R21206 VSS.n3323 VSS.n2856 0.0152714
R21207 VSS.n3341 VSS.n3340 0.0152714
R21208 VSS.n3671 VSS.n3670 0.0152714
R21209 VSS.n3703 VSS.n3702 0.0152714
R21210 VSS.n3767 VSS.n3763 0.0152714
R21211 VSS.n3794 VSS.n3793 0.0152714
R21212 VSS.n3915 VSS.n3448 0.0152714
R21213 VSS.n3933 VSS.n3932 0.0152714
R21214 VSS.n4263 VSS.n4262 0.0152714
R21215 VSS.n4295 VSS.n4294 0.0152714
R21216 VSS.n4359 VSS.n4355 0.0152714
R21217 VSS.n4386 VSS.n4385 0.0152714
R21218 VSS.n4507 VSS.n4040 0.0152714
R21219 VSS.n4525 VSS.n4524 0.0152714
R21220 VSS.n4855 VSS.n4854 0.0152714
R21221 VSS.n4887 VSS.n4886 0.0152714
R21222 VSS.n4951 VSS.n4947 0.0152714
R21223 VSS.n4978 VSS.n4977 0.0152714
R21224 VSS.n5099 VSS.n4632 0.0152714
R21225 VSS.n5117 VSS.n5116 0.0152714
R21226 VSS.n2476 VSS.n2475 0.0152714
R21227 VSS.n2508 VSS.n2507 0.0152714
R21228 VSS.n5300 VSS.n5299 0.0152714
R21229 VSS.n5284 VSS.n5283 0.0152714
R21230 VSS.n2746 VSS.n2727 0.0152714
R21231 VSS.n5221 VSS.n5220 0.0152714
R21232 VSS.n5437 VSS.n5436 0.0152714
R21233 VSS.n5469 VSS.n5468 0.0152714
R21234 VSS.n5873 VSS.n5872 0.0152714
R21235 VSS.n5857 VSS.n5856 0.0152714
R21236 VSS.n5707 VSS.n5688 0.0152714
R21237 VSS.n5794 VSS.n5793 0.0152714
R21238 VSS.n6010 VSS.n6009 0.0152714
R21239 VSS.n6042 VSS.n6041 0.0152714
R21240 VSS.n6465 VSS.n6464 0.0152714
R21241 VSS.n6449 VSS.n6448 0.0152714
R21242 VSS.n6280 VSS.n6261 0.0152714
R21243 VSS.n6386 VSS.n6385 0.0152714
R21244 VSS.n7812 VSS.n7811 0.0152714
R21245 VSS.n7844 VSS.n7843 0.0152714
R21246 VSS.n7908 VSS.n7904 0.0152714
R21247 VSS.n7935 VSS.n7934 0.0152714
R21248 VSS.n8056 VSS.n7589 0.0152714
R21249 VSS.n8074 VSS.n8073 0.0152714
R21250 VSS.n8404 VSS.n8403 0.0152714
R21251 VSS.n8436 VSS.n8435 0.0152714
R21252 VSS.n8500 VSS.n8496 0.0152714
R21253 VSS.n8527 VSS.n8526 0.0152714
R21254 VSS.n8648 VSS.n8181 0.0152714
R21255 VSS.n8666 VSS.n8665 0.0152714
R21256 VSS.n8996 VSS.n8995 0.0152714
R21257 VSS.n9028 VSS.n9027 0.0152714
R21258 VSS.n9092 VSS.n9088 0.0152714
R21259 VSS.n9119 VSS.n9118 0.0152714
R21260 VSS.n9240 VSS.n8773 0.0152714
R21261 VSS.n9258 VSS.n9257 0.0152714
R21262 VSS.n10180 VSS.n10179 0.0152714
R21263 VSS.n10212 VSS.n10211 0.0152714
R21264 VSS.n10276 VSS.n10272 0.0152714
R21265 VSS.n10303 VSS.n10302 0.0152714
R21266 VSS.n10424 VSS.n9957 0.0152714
R21267 VSS.n10442 VSS.n10441 0.0152714
R21268 VSS.n10772 VSS.n10771 0.0152714
R21269 VSS.n10804 VSS.n10803 0.0152714
R21270 VSS.n10868 VSS.n10864 0.0152714
R21271 VSS.n10895 VSS.n10894 0.0152714
R21272 VSS.n11016 VSS.n10549 0.0152714
R21273 VSS.n11034 VSS.n11033 0.0152714
R21274 VSS.n11364 VSS.n11363 0.0152714
R21275 VSS.n11396 VSS.n11395 0.0152714
R21276 VSS.n11460 VSS.n11456 0.0152714
R21277 VSS.n11487 VSS.n11486 0.0152714
R21278 VSS.n11608 VSS.n11141 0.0152714
R21279 VSS.n11626 VSS.n11625 0.0152714
R21280 VSS.n11956 VSS.n11955 0.0152714
R21281 VSS.n11988 VSS.n11987 0.0152714
R21282 VSS.n12052 VSS.n12048 0.0152714
R21283 VSS.n12079 VSS.n12078 0.0152714
R21284 VSS.n12200 VSS.n11733 0.0152714
R21285 VSS.n12218 VSS.n12217 0.0152714
R21286 VSS.n12548 VSS.n12547 0.0152714
R21287 VSS.n12580 VSS.n12579 0.0152714
R21288 VSS.n12644 VSS.n12640 0.0152714
R21289 VSS.n12671 VSS.n12670 0.0152714
R21290 VSS.n12792 VSS.n12325 0.0152714
R21291 VSS.n12810 VSS.n12809 0.0152714
R21292 VSS.n13140 VSS.n13139 0.0152714
R21293 VSS.n13172 VSS.n13171 0.0152714
R21294 VSS.n13236 VSS.n13232 0.0152714
R21295 VSS.n13263 VSS.n13262 0.0152714
R21296 VSS.n13384 VSS.n12917 0.0152714
R21297 VSS.n13402 VSS.n13401 0.0152714
R21298 VSS.n13732 VSS.n13731 0.0152714
R21299 VSS.n13764 VSS.n13763 0.0152714
R21300 VSS.n13828 VSS.n13824 0.0152714
R21301 VSS.n13855 VSS.n13854 0.0152714
R21302 VSS.n13976 VSS.n13509 0.0152714
R21303 VSS.n13994 VSS.n13993 0.0152714
R21304 VSS.n14324 VSS.n14323 0.0152714
R21305 VSS.n14356 VSS.n14355 0.0152714
R21306 VSS.n14420 VSS.n14416 0.0152714
R21307 VSS.n14447 VSS.n14446 0.0152714
R21308 VSS.n14568 VSS.n14101 0.0152714
R21309 VSS.n14586 VSS.n14585 0.0152714
R21310 VSS.n14916 VSS.n14915 0.0152714
R21311 VSS.n14948 VSS.n14947 0.0152714
R21312 VSS.n15012 VSS.n15008 0.0152714
R21313 VSS.n15039 VSS.n15038 0.0152714
R21314 VSS.n15160 VSS.n14693 0.0152714
R21315 VSS.n15178 VSS.n15177 0.0152714
R21316 VSS.n15508 VSS.n15507 0.0152714
R21317 VSS.n15540 VSS.n15539 0.0152714
R21318 VSS.n15604 VSS.n15600 0.0152714
R21319 VSS.n15631 VSS.n15630 0.0152714
R21320 VSS.n15752 VSS.n15285 0.0152714
R21321 VSS.n15770 VSS.n15769 0.0152714
R21322 VSS.n6616 VSS.n6615 0.0152714
R21323 VSS.n6648 VSS.n6647 0.0152714
R21324 VSS.n15953 VSS.n15952 0.0152714
R21325 VSS.n15937 VSS.n15936 0.0152714
R21326 VSS.n6886 VSS.n6867 0.0152714
R21327 VSS.n15874 VSS.n15873 0.0152714
R21328 VSS.n7211 VSS.n7207 0.0152714
R21329 VSS.n7238 VSS.n7237 0.0152714
R21330 VSS.n7316 VSS.n7312 0.0152714
R21331 VSS.n7343 VSS.n7342 0.0152714
R21332 VSS.n7464 VSS.n6996 0.0152714
R21333 VSS.n7482 VSS.n7481 0.0152714
R21334 VSS.n439 VSS.n438 0.0152714
R21335 VSS.n423 VSS.n422 0.0152714
R21336 VSS.n18628 VSS.n18624 0.0152714
R21337 VSS.n18655 VSS.n18654 0.0152714
R21338 VSS.n18776 VSS.n94 0.0152714
R21339 VSS.n18794 VSS.n18793 0.0152714
R21340 VSS.n1004 VSS.n1003 0.0152714
R21341 VSS.n988 VSS.n987 0.0152714
R21342 VSS.n867 VSS.n866 0.0152714
R21343 VSS.n851 VSS.n850 0.0152714
R21344 VSS.n709 VSS.n690 0.0152714
R21345 VSS.n788 VSS.n787 0.0152714
R21346 VSS.n17981 VSS.n17980 0.0152714
R21347 VSS.n17965 VSS.n17964 0.0152714
R21348 VSS.n1368 VSS.n1349 0.0152714
R21349 VSS.n17902 VSS.n17901 0.0152714
R21350 VSS.n9588 VSS.n9587 0.0151667
R21351 VSS.n9620 VSS.n9619 0.0151667
R21352 VSS.n17177 VSS.n16906 0.0147857
R21353 VSS.n17194 VSS.n16888 0.0147857
R21354 VSS.n17769 VSS.n17320 0.0147857
R21355 VSS.n17786 VSS.n17302 0.0147857
R21356 VSS.n18349 VSS.n18346 0.0147857
R21357 VSS.n18412 VSS.n18390 0.0147857
R21358 VSS.n9819 VSS.n9370 0.0147857
R21359 VSS.n9836 VSS.n9352 0.0147857
R21360 VSS.n16762 VSS.n16312 0.0147857
R21361 VSS.n16779 VSS.n16294 0.0147857
R21362 VSS.n16169 VSS.n1484 0.0147857
R21363 VSS.n16186 VSS.n1466 0.0147857
R21364 VSS.n2137 VSS.n2111 0.0147857
R21365 VSS.n2166 VSS.n2165 0.0147857
R21366 VSS.n3310 VSS.n2861 0.0147857
R21367 VSS.n3327 VSS.n2843 0.0147857
R21368 VSS.n3902 VSS.n3453 0.0147857
R21369 VSS.n3919 VSS.n3435 0.0147857
R21370 VSS.n4494 VSS.n4045 0.0147857
R21371 VSS.n4511 VSS.n4027 0.0147857
R21372 VSS.n5086 VSS.n4637 0.0147857
R21373 VSS.n5103 VSS.n4619 0.0147857
R21374 VSS.n2733 VSS.n2707 0.0147857
R21375 VSS.n2762 VSS.n2761 0.0147857
R21376 VSS.n5694 VSS.n5668 0.0147857
R21377 VSS.n5723 VSS.n5722 0.0147857
R21378 VSS.n6267 VSS.n6241 0.0147857
R21379 VSS.n6296 VSS.n6295 0.0147857
R21380 VSS.n8043 VSS.n7594 0.0147857
R21381 VSS.n8060 VSS.n7576 0.0147857
R21382 VSS.n8635 VSS.n8186 0.0147857
R21383 VSS.n8652 VSS.n8168 0.0147857
R21384 VSS.n9227 VSS.n8778 0.0147857
R21385 VSS.n9244 VSS.n8760 0.0147857
R21386 VSS.n10411 VSS.n9962 0.0147857
R21387 VSS.n10428 VSS.n9944 0.0147857
R21388 VSS.n11003 VSS.n10554 0.0147857
R21389 VSS.n11020 VSS.n10536 0.0147857
R21390 VSS.n11595 VSS.n11146 0.0147857
R21391 VSS.n11612 VSS.n11128 0.0147857
R21392 VSS.n12187 VSS.n11738 0.0147857
R21393 VSS.n12204 VSS.n11720 0.0147857
R21394 VSS.n12779 VSS.n12330 0.0147857
R21395 VSS.n12796 VSS.n12312 0.0147857
R21396 VSS.n13371 VSS.n12922 0.0147857
R21397 VSS.n13388 VSS.n12904 0.0147857
R21398 VSS.n13963 VSS.n13514 0.0147857
R21399 VSS.n13980 VSS.n13496 0.0147857
R21400 VSS.n14555 VSS.n14106 0.0147857
R21401 VSS.n14572 VSS.n14088 0.0147857
R21402 VSS.n15147 VSS.n14698 0.0147857
R21403 VSS.n15164 VSS.n14680 0.0147857
R21404 VSS.n15739 VSS.n15290 0.0147857
R21405 VSS.n15756 VSS.n15272 0.0147857
R21406 VSS.n6873 VSS.n6847 0.0147857
R21407 VSS.n6902 VSS.n6901 0.0147857
R21408 VSS.n7451 VSS.n7001 0.0147857
R21409 VSS.n7468 VSS.n6983 0.0147857
R21410 VSS.n18763 VSS.n99 0.0147857
R21411 VSS.n18780 VSS.n81 0.0147857
R21412 VSS.n696 VSS.n670 0.0147857
R21413 VSS.n725 VSS.n724 0.0147857
R21414 VSS.n1355 VSS.n1329 0.0147857
R21415 VSS.n1384 VSS.n1383 0.0147857
R21416 VSS.n17250 VSS.n17249 0.0138929
R21417 VSS.n17842 VSS.n17841 0.0138929
R21418 VSS.n18433 VSS.n18426 0.0138929
R21419 VSS.n9893 VSS.n9892 0.0138929
R21420 VSS.n16836 VSS.n16835 0.0138929
R21421 VSS.n16243 VSS.n16242 0.0138929
R21422 VSS.n2213 VSS.n2200 0.0138929
R21423 VSS.n3384 VSS.n3383 0.0138929
R21424 VSS.n3976 VSS.n3975 0.0138929
R21425 VSS.n4568 VSS.n4567 0.0138929
R21426 VSS.n5160 VSS.n5159 0.0138929
R21427 VSS.n2809 VSS.n2796 0.0138929
R21428 VSS.n5735 VSS.n5734 0.0138929
R21429 VSS.n6343 VSS.n6330 0.0138929
R21430 VSS.n8117 VSS.n8116 0.0138929
R21431 VSS.n8709 VSS.n8708 0.0138929
R21432 VSS.n9301 VSS.n9300 0.0138929
R21433 VSS.n10485 VSS.n10484 0.0138929
R21434 VSS.n11077 VSS.n11076 0.0138929
R21435 VSS.n11669 VSS.n11668 0.0138929
R21436 VSS.n12261 VSS.n12260 0.0138929
R21437 VSS.n12853 VSS.n12852 0.0138929
R21438 VSS.n13445 VSS.n13444 0.0138929
R21439 VSS.n14037 VSS.n14036 0.0138929
R21440 VSS.n14629 VSS.n14628 0.0138929
R21441 VSS.n15221 VSS.n15220 0.0138929
R21442 VSS.n15813 VSS.n15812 0.0138929
R21443 VSS.n6949 VSS.n6936 0.0138929
R21444 VSS.n7525 VSS.n7524 0.0138929
R21445 VSS.n18837 VSS.n18836 0.0138929
R21446 VSS.n736 VSS.n49 0.0138929
R21447 VSS.n1431 VSS.n1418 0.0138929
R21448 VSS.n18022 VSS.n18021 0.0132571
R21449 VSS.n17060 VSS.n17059 0.0132571
R21450 VSS.n17146 VSS.n17144 0.0132571
R21451 VSS.n17174 VSS.n16907 0.0132571
R21452 VSS.n17227 VSS.n17226 0.0132571
R21453 VSS.n17247 VSS.n17245 0.0132571
R21454 VSS.n17550 VSS.n17546 0.0132571
R21455 VSS.n17652 VSS.n17651 0.0132571
R21456 VSS.n17738 VSS.n17736 0.0132571
R21457 VSS.n17766 VSS.n17321 0.0132571
R21458 VSS.n17819 VSS.n17818 0.0132571
R21459 VSS.n17839 VSS.n17837 0.0132571
R21460 VSS.n18127 VSS.n18123 0.0132571
R21461 VSS.n18562 VSS.n18561 0.0132571
R21462 VSS.n18522 VSS.n18336 0.0132571
R21463 VSS.n18520 VSS.n18337 0.0132571
R21464 VSS.n18486 VSS.n18485 0.0132571
R21465 VSS.n18470 VSS.n18428 0.0132571
R21466 VSS.n9702 VSS.n9701 0.0132571
R21467 VSS.n9788 VSS.n9786 0.0132571
R21468 VSS.n9816 VSS.n9371 0.0132571
R21469 VSS.n9869 VSS.n9868 0.0132571
R21470 VSS.n9888 VSS.n9887 0.0132571
R21471 VSS.n16540 VSS.n16539 0.0132571
R21472 VSS.n16645 VSS.n16644 0.0132571
R21473 VSS.n16731 VSS.n16729 0.0132571
R21474 VSS.n16759 VSS.n16313 0.0132571
R21475 VSS.n16812 VSS.n16811 0.0132571
R21476 VSS.n16831 VSS.n16830 0.0132571
R21477 VSS.n1705 VSS.n1704 0.0132571
R21478 VSS.n16052 VSS.n16051 0.0132571
R21479 VSS.n16138 VSS.n16136 0.0132571
R21480 VSS.n16166 VSS.n1485 0.0132571
R21481 VSS.n16219 VSS.n16218 0.0132571
R21482 VSS.n16238 VSS.n16237 0.0132571
R21483 VSS.n1892 VSS.n1888 0.0132571
R21484 VSS.n2327 VSS.n2326 0.0132571
R21485 VSS.n2101 VSS.n2100 0.0132571
R21486 VSS.n2118 VSS.n2117 0.0132571
R21487 VSS.n2239 VSS.n2168 0.0132571
R21488 VSS.n2237 VSS.n2169 0.0132571
R21489 VSS.n3091 VSS.n3087 0.0132571
R21490 VSS.n3193 VSS.n3192 0.0132571
R21491 VSS.n3279 VSS.n3277 0.0132571
R21492 VSS.n3307 VSS.n2862 0.0132571
R21493 VSS.n3360 VSS.n3359 0.0132571
R21494 VSS.n3379 VSS.n3378 0.0132571
R21495 VSS.n3683 VSS.n3679 0.0132571
R21496 VSS.n3785 VSS.n3784 0.0132571
R21497 VSS.n3871 VSS.n3869 0.0132571
R21498 VSS.n3899 VSS.n3454 0.0132571
R21499 VSS.n3952 VSS.n3951 0.0132571
R21500 VSS.n3971 VSS.n3970 0.0132571
R21501 VSS.n4275 VSS.n4271 0.0132571
R21502 VSS.n4377 VSS.n4376 0.0132571
R21503 VSS.n4463 VSS.n4461 0.0132571
R21504 VSS.n4491 VSS.n4046 0.0132571
R21505 VSS.n4544 VSS.n4543 0.0132571
R21506 VSS.n4563 VSS.n4562 0.0132571
R21507 VSS.n4867 VSS.n4863 0.0132571
R21508 VSS.n4969 VSS.n4968 0.0132571
R21509 VSS.n5055 VSS.n5053 0.0132571
R21510 VSS.n5083 VSS.n4638 0.0132571
R21511 VSS.n5136 VSS.n5135 0.0132571
R21512 VSS.n5155 VSS.n5154 0.0132571
R21513 VSS.n2488 VSS.n2484 0.0132571
R21514 VSS.n5292 VSS.n5291 0.0132571
R21515 VSS.n2697 VSS.n2696 0.0132571
R21516 VSS.n2714 VSS.n2713 0.0132571
R21517 VSS.n5204 VSS.n2764 0.0132571
R21518 VSS.n5202 VSS.n2765 0.0132571
R21519 VSS.n5449 VSS.n5445 0.0132571
R21520 VSS.n5865 VSS.n5864 0.0132571
R21521 VSS.n5658 VSS.n5657 0.0132571
R21522 VSS.n5675 VSS.n5674 0.0132571
R21523 VSS.n5777 VSS.n5725 0.0132571
R21524 VSS.n5775 VSS.n5726 0.0132571
R21525 VSS.n6022 VSS.n6018 0.0132571
R21526 VSS.n6457 VSS.n6456 0.0132571
R21527 VSS.n6231 VSS.n6230 0.0132571
R21528 VSS.n6248 VSS.n6247 0.0132571
R21529 VSS.n6369 VSS.n6298 0.0132571
R21530 VSS.n6367 VSS.n6299 0.0132571
R21531 VSS.n7824 VSS.n7820 0.0132571
R21532 VSS.n7926 VSS.n7925 0.0132571
R21533 VSS.n8012 VSS.n8010 0.0132571
R21534 VSS.n8040 VSS.n7595 0.0132571
R21535 VSS.n8093 VSS.n8092 0.0132571
R21536 VSS.n8112 VSS.n8111 0.0132571
R21537 VSS.n8416 VSS.n8412 0.0132571
R21538 VSS.n8518 VSS.n8517 0.0132571
R21539 VSS.n8604 VSS.n8602 0.0132571
R21540 VSS.n8632 VSS.n8187 0.0132571
R21541 VSS.n8685 VSS.n8684 0.0132571
R21542 VSS.n8704 VSS.n8703 0.0132571
R21543 VSS.n9008 VSS.n9004 0.0132571
R21544 VSS.n9110 VSS.n9109 0.0132571
R21545 VSS.n9196 VSS.n9194 0.0132571
R21546 VSS.n9224 VSS.n8779 0.0132571
R21547 VSS.n9277 VSS.n9276 0.0132571
R21548 VSS.n9296 VSS.n9295 0.0132571
R21549 VSS.n10192 VSS.n10188 0.0132571
R21550 VSS.n10294 VSS.n10293 0.0132571
R21551 VSS.n10380 VSS.n10378 0.0132571
R21552 VSS.n10408 VSS.n9963 0.0132571
R21553 VSS.n10461 VSS.n10460 0.0132571
R21554 VSS.n10480 VSS.n10479 0.0132571
R21555 VSS.n10784 VSS.n10780 0.0132571
R21556 VSS.n10886 VSS.n10885 0.0132571
R21557 VSS.n10972 VSS.n10970 0.0132571
R21558 VSS.n11000 VSS.n10555 0.0132571
R21559 VSS.n11053 VSS.n11052 0.0132571
R21560 VSS.n11072 VSS.n11071 0.0132571
R21561 VSS.n11376 VSS.n11372 0.0132571
R21562 VSS.n11478 VSS.n11477 0.0132571
R21563 VSS.n11564 VSS.n11562 0.0132571
R21564 VSS.n11592 VSS.n11147 0.0132571
R21565 VSS.n11645 VSS.n11644 0.0132571
R21566 VSS.n11664 VSS.n11663 0.0132571
R21567 VSS.n11968 VSS.n11964 0.0132571
R21568 VSS.n12070 VSS.n12069 0.0132571
R21569 VSS.n12156 VSS.n12154 0.0132571
R21570 VSS.n12184 VSS.n11739 0.0132571
R21571 VSS.n12237 VSS.n12236 0.0132571
R21572 VSS.n12256 VSS.n12255 0.0132571
R21573 VSS.n12560 VSS.n12556 0.0132571
R21574 VSS.n12662 VSS.n12661 0.0132571
R21575 VSS.n12748 VSS.n12746 0.0132571
R21576 VSS.n12776 VSS.n12331 0.0132571
R21577 VSS.n12829 VSS.n12828 0.0132571
R21578 VSS.n12848 VSS.n12847 0.0132571
R21579 VSS.n13152 VSS.n13148 0.0132571
R21580 VSS.n13254 VSS.n13253 0.0132571
R21581 VSS.n13340 VSS.n13338 0.0132571
R21582 VSS.n13368 VSS.n12923 0.0132571
R21583 VSS.n13421 VSS.n13420 0.0132571
R21584 VSS.n13440 VSS.n13439 0.0132571
R21585 VSS.n13744 VSS.n13740 0.0132571
R21586 VSS.n13846 VSS.n13845 0.0132571
R21587 VSS.n13932 VSS.n13930 0.0132571
R21588 VSS.n13960 VSS.n13515 0.0132571
R21589 VSS.n14013 VSS.n14012 0.0132571
R21590 VSS.n14032 VSS.n14031 0.0132571
R21591 VSS.n14336 VSS.n14332 0.0132571
R21592 VSS.n14438 VSS.n14437 0.0132571
R21593 VSS.n14524 VSS.n14522 0.0132571
R21594 VSS.n14552 VSS.n14107 0.0132571
R21595 VSS.n14605 VSS.n14604 0.0132571
R21596 VSS.n14624 VSS.n14623 0.0132571
R21597 VSS.n14928 VSS.n14924 0.0132571
R21598 VSS.n15030 VSS.n15029 0.0132571
R21599 VSS.n15116 VSS.n15114 0.0132571
R21600 VSS.n15144 VSS.n14699 0.0132571
R21601 VSS.n15197 VSS.n15196 0.0132571
R21602 VSS.n15216 VSS.n15215 0.0132571
R21603 VSS.n15520 VSS.n15516 0.0132571
R21604 VSS.n15622 VSS.n15621 0.0132571
R21605 VSS.n15708 VSS.n15706 0.0132571
R21606 VSS.n15736 VSS.n15291 0.0132571
R21607 VSS.n15789 VSS.n15788 0.0132571
R21608 VSS.n15808 VSS.n15807 0.0132571
R21609 VSS.n6628 VSS.n6624 0.0132571
R21610 VSS.n15945 VSS.n15944 0.0132571
R21611 VSS.n6837 VSS.n6836 0.0132571
R21612 VSS.n6854 VSS.n6853 0.0132571
R21613 VSS.n15857 VSS.n6904 0.0132571
R21614 VSS.n15855 VSS.n6905 0.0132571
R21615 VSS.n7229 VSS.n7228 0.0132571
R21616 VSS.n7334 VSS.n7333 0.0132571
R21617 VSS.n7420 VSS.n7418 0.0132571
R21618 VSS.n7448 VSS.n7002 0.0132571
R21619 VSS.n7501 VSS.n7500 0.0132571
R21620 VSS.n7520 VSS.n7519 0.0132571
R21621 VSS.n431 VSS.n430 0.0132571
R21622 VSS.n18646 VSS.n18645 0.0132571
R21623 VSS.n18732 VSS.n18730 0.0132571
R21624 VSS.n18760 VSS.n100 0.0132571
R21625 VSS.n18813 VSS.n18812 0.0132571
R21626 VSS.n18832 VSS.n18831 0.0132571
R21627 VSS.n996 VSS.n995 0.0132571
R21628 VSS.n859 VSS.n858 0.0132571
R21629 VSS.n660 VSS.n659 0.0132571
R21630 VSS.n677 VSS.n676 0.0132571
R21631 VSS.n771 VSS.n727 0.0132571
R21632 VSS.n769 VSS.n728 0.0132571
R21633 VSS.n17973 VSS.n17972 0.0132571
R21634 VSS.n1319 VSS.n1318 0.0132571
R21635 VSS.n1336 VSS.n1335 0.0132571
R21636 VSS.n17885 VSS.n1386 0.0132571
R21637 VSS.n17883 VSS.n1387 0.0132571
R21638 VSS.n9600 VSS.n9596 0.0131667
R21639 VSS.n1281 VSS.n1203 0.013
R21640 VSS.n17955 VSS.n17954 0.013
R21641 VSS.n1280 VSS.n1279 0.013
R21642 VSS.n1015 VSS.n457 0.013
R21643 VSS.n915 VSS.n913 0.013
R21644 VSS.n17098 VSS.n16942 0.013
R21645 VSS.n17131 VSS.n16934 0.013
R21646 VSS.n18041 VSS.n1024 0.013
R21647 VSS.n1096 VSS.n1094 0.013
R21648 VSS.n1097 VSS.n1091 0.013
R21649 VSS.n17097 VSS.n17096 0.013
R21650 VSS.n17690 VSS.n17356 0.013
R21651 VSS.n17723 VSS.n17348 0.013
R21652 VSS.n17512 VSS.n17504 0.013
R21653 VSS.n17510 VSS.n17506 0.013
R21654 VSS.n17509 VSS.n17508 0.013
R21655 VSS.n17689 VSS.n17688 0.013
R21656 VSS.n18089 VSS.n18081 0.013
R21657 VSS.n18087 VSS.n18083 0.013
R21658 VSS.n18298 VSS.n18220 0.013
R21659 VSS.n18544 VSS.n18543 0.013
R21660 VSS.n18297 VSS.n18296 0.013
R21661 VSS.n18086 VSS.n18085 0.013
R21662 VSS.n9562 VSS.n9554 0.013
R21663 VSS.n9560 VSS.n9556 0.013
R21664 VSS.n9740 VSS.n9406 0.013
R21665 VSS.n9773 VSS.n9398 0.013
R21666 VSS.n9739 VSS.n9738 0.013
R21667 VSS.n9559 VSS.n9558 0.013
R21668 VSS.n16498 VSS.n16490 0.013
R21669 VSS.n16496 VSS.n16492 0.013
R21670 VSS.n16683 VSS.n16348 0.013
R21671 VSS.n16716 VSS.n16340 0.013
R21672 VSS.n16682 VSS.n16681 0.013
R21673 VSS.n16495 VSS.n16494 0.013
R21674 VSS.n1663 VSS.n1655 0.013
R21675 VSS.n1661 VSS.n1657 0.013
R21676 VSS.n16090 VSS.n1520 0.013
R21677 VSS.n16123 VSS.n1512 0.013
R21678 VSS.n16089 VSS.n16088 0.013
R21679 VSS.n1660 VSS.n1659 0.013
R21680 VSS.n1854 VSS.n1846 0.013
R21681 VSS.n1852 VSS.n1848 0.013
R21682 VSS.n2063 VSS.n1985 0.013
R21683 VSS.n2309 VSS.n2308 0.013
R21684 VSS.n2062 VSS.n2061 0.013
R21685 VSS.n1851 VSS.n1850 0.013
R21686 VSS.n3053 VSS.n3045 0.013
R21687 VSS.n3051 VSS.n3047 0.013
R21688 VSS.n3231 VSS.n2897 0.013
R21689 VSS.n3264 VSS.n2889 0.013
R21690 VSS.n3230 VSS.n3229 0.013
R21691 VSS.n3050 VSS.n3049 0.013
R21692 VSS.n3645 VSS.n3637 0.013
R21693 VSS.n3643 VSS.n3639 0.013
R21694 VSS.n3823 VSS.n3489 0.013
R21695 VSS.n3856 VSS.n3481 0.013
R21696 VSS.n3822 VSS.n3821 0.013
R21697 VSS.n3642 VSS.n3641 0.013
R21698 VSS.n4237 VSS.n4229 0.013
R21699 VSS.n4235 VSS.n4231 0.013
R21700 VSS.n4415 VSS.n4081 0.013
R21701 VSS.n4448 VSS.n4073 0.013
R21702 VSS.n4414 VSS.n4413 0.013
R21703 VSS.n4234 VSS.n4233 0.013
R21704 VSS.n4829 VSS.n4821 0.013
R21705 VSS.n4827 VSS.n4823 0.013
R21706 VSS.n5007 VSS.n4673 0.013
R21707 VSS.n5040 VSS.n4665 0.013
R21708 VSS.n5006 VSS.n5005 0.013
R21709 VSS.n4826 VSS.n4825 0.013
R21710 VSS.n2450 VSS.n2442 0.013
R21711 VSS.n2448 VSS.n2444 0.013
R21712 VSS.n2659 VSS.n2581 0.013
R21713 VSS.n5274 VSS.n5273 0.013
R21714 VSS.n2658 VSS.n2657 0.013
R21715 VSS.n2447 VSS.n2446 0.013
R21716 VSS.n5411 VSS.n5403 0.013
R21717 VSS.n5409 VSS.n5405 0.013
R21718 VSS.n5620 VSS.n5542 0.013
R21719 VSS.n5847 VSS.n5846 0.013
R21720 VSS.n5619 VSS.n5618 0.013
R21721 VSS.n5408 VSS.n5407 0.013
R21722 VSS.n5984 VSS.n5976 0.013
R21723 VSS.n5982 VSS.n5978 0.013
R21724 VSS.n6193 VSS.n6115 0.013
R21725 VSS.n6439 VSS.n6438 0.013
R21726 VSS.n6192 VSS.n6191 0.013
R21727 VSS.n5981 VSS.n5980 0.013
R21728 VSS.n7786 VSS.n7778 0.013
R21729 VSS.n7784 VSS.n7780 0.013
R21730 VSS.n7964 VSS.n7630 0.013
R21731 VSS.n7997 VSS.n7622 0.013
R21732 VSS.n7963 VSS.n7962 0.013
R21733 VSS.n7783 VSS.n7782 0.013
R21734 VSS.n8378 VSS.n8370 0.013
R21735 VSS.n8376 VSS.n8372 0.013
R21736 VSS.n8556 VSS.n8222 0.013
R21737 VSS.n8589 VSS.n8214 0.013
R21738 VSS.n8555 VSS.n8554 0.013
R21739 VSS.n8375 VSS.n8374 0.013
R21740 VSS.n8970 VSS.n8962 0.013
R21741 VSS.n8968 VSS.n8964 0.013
R21742 VSS.n9148 VSS.n8814 0.013
R21743 VSS.n9181 VSS.n8806 0.013
R21744 VSS.n9147 VSS.n9146 0.013
R21745 VSS.n8967 VSS.n8966 0.013
R21746 VSS.n10154 VSS.n10146 0.013
R21747 VSS.n10152 VSS.n10148 0.013
R21748 VSS.n10332 VSS.n9998 0.013
R21749 VSS.n10365 VSS.n9990 0.013
R21750 VSS.n10331 VSS.n10330 0.013
R21751 VSS.n10151 VSS.n10150 0.013
R21752 VSS.n10746 VSS.n10738 0.013
R21753 VSS.n10744 VSS.n10740 0.013
R21754 VSS.n10924 VSS.n10590 0.013
R21755 VSS.n10957 VSS.n10582 0.013
R21756 VSS.n10923 VSS.n10922 0.013
R21757 VSS.n10743 VSS.n10742 0.013
R21758 VSS.n11338 VSS.n11330 0.013
R21759 VSS.n11336 VSS.n11332 0.013
R21760 VSS.n11516 VSS.n11182 0.013
R21761 VSS.n11549 VSS.n11174 0.013
R21762 VSS.n11515 VSS.n11514 0.013
R21763 VSS.n11335 VSS.n11334 0.013
R21764 VSS.n11930 VSS.n11922 0.013
R21765 VSS.n11928 VSS.n11924 0.013
R21766 VSS.n12108 VSS.n11774 0.013
R21767 VSS.n12141 VSS.n11766 0.013
R21768 VSS.n12107 VSS.n12106 0.013
R21769 VSS.n11927 VSS.n11926 0.013
R21770 VSS.n12522 VSS.n12514 0.013
R21771 VSS.n12520 VSS.n12516 0.013
R21772 VSS.n12700 VSS.n12366 0.013
R21773 VSS.n12733 VSS.n12358 0.013
R21774 VSS.n12699 VSS.n12698 0.013
R21775 VSS.n12519 VSS.n12518 0.013
R21776 VSS.n13114 VSS.n13106 0.013
R21777 VSS.n13112 VSS.n13108 0.013
R21778 VSS.n13292 VSS.n12958 0.013
R21779 VSS.n13325 VSS.n12950 0.013
R21780 VSS.n13291 VSS.n13290 0.013
R21781 VSS.n13111 VSS.n13110 0.013
R21782 VSS.n13706 VSS.n13698 0.013
R21783 VSS.n13704 VSS.n13700 0.013
R21784 VSS.n13884 VSS.n13550 0.013
R21785 VSS.n13917 VSS.n13542 0.013
R21786 VSS.n13883 VSS.n13882 0.013
R21787 VSS.n13703 VSS.n13702 0.013
R21788 VSS.n14298 VSS.n14290 0.013
R21789 VSS.n14296 VSS.n14292 0.013
R21790 VSS.n14476 VSS.n14142 0.013
R21791 VSS.n14509 VSS.n14134 0.013
R21792 VSS.n14475 VSS.n14474 0.013
R21793 VSS.n14295 VSS.n14294 0.013
R21794 VSS.n14890 VSS.n14882 0.013
R21795 VSS.n14888 VSS.n14884 0.013
R21796 VSS.n15068 VSS.n14734 0.013
R21797 VSS.n15101 VSS.n14726 0.013
R21798 VSS.n15067 VSS.n15066 0.013
R21799 VSS.n14887 VSS.n14886 0.013
R21800 VSS.n15482 VSS.n15474 0.013
R21801 VSS.n15480 VSS.n15476 0.013
R21802 VSS.n15660 VSS.n15326 0.013
R21803 VSS.n15693 VSS.n15318 0.013
R21804 VSS.n15659 VSS.n15658 0.013
R21805 VSS.n15479 VSS.n15478 0.013
R21806 VSS.n6590 VSS.n6582 0.013
R21807 VSS.n6588 VSS.n6584 0.013
R21808 VSS.n6799 VSS.n6721 0.013
R21809 VSS.n15927 VSS.n15926 0.013
R21810 VSS.n6798 VSS.n6797 0.013
R21811 VSS.n6587 VSS.n6586 0.013
R21812 VSS.n7187 VSS.n7179 0.013
R21813 VSS.n7185 VSS.n7181 0.013
R21814 VSS.n7372 VSS.n7037 0.013
R21815 VSS.n7405 VSS.n7029 0.013
R21816 VSS.n7371 VSS.n7370 0.013
R21817 VSS.n7184 VSS.n7183 0.013
R21818 VSS.n450 VSS.n291 0.013
R21819 VSS.n349 VSS.n345 0.013
R21820 VSS.n18684 VSS.n135 0.013
R21821 VSS.n18717 VSS.n127 0.013
R21822 VSS.n18683 VSS.n18682 0.013
R21823 VSS.n351 VSS.n350 0.013
R21824 VSS.n622 VSS.n541 0.013
R21825 VSS.n841 VSS.n840 0.013
R21826 VSS.n621 VSS.n620 0.013
R21827 VSS.n916 VSS.n910 0.013
R21828 VSS.n17992 VSS.n1159 0.0121071
R21829 VSS.n1229 VSS.n1227 0.0121071
R21830 VSS.n1230 VSS.n1224 0.0121071
R21831 VSS.n1204 VSS.n1190 0.0121071
R21832 VSS.n919 VSS.n463 0.0121071
R21833 VSS.n966 VSS.n888 0.0121071
R21834 VSS.n978 VSS.n977 0.0121071
R21835 VSS.n17018 VSS.n17010 0.0121071
R21836 VSS.n17016 VSS.n17012 0.0121071
R21837 VSS.n1100 VSS.n1030 0.0121071
R21838 VSS.n1147 VSS.n1069 0.0121071
R21839 VSS.n18004 VSS.n18003 0.0121071
R21840 VSS.n1099 VSS.n1028 0.0121071
R21841 VSS.n1146 VSS.n1145 0.0121071
R21842 VSS.n17138 VSS.n16930 0.0121071
R21843 VSS.n17015 VSS.n17014 0.0121071
R21844 VSS.n16949 VSS.n16946 0.0121071
R21845 VSS.n17610 VSS.n17602 0.0121071
R21846 VSS.n17608 VSS.n17604 0.0121071
R21847 VSS.n17519 VSS.n17518 0.0121071
R21848 VSS.n17582 VSS.n17581 0.0121071
R21849 VSS.n17597 VSS.n17423 0.0121071
R21850 VSS.n17517 VSS.n17485 0.0121071
R21851 VSS.n17583 VSS.n17433 0.0121071
R21852 VSS.n17730 VSS.n17344 0.0121071
R21853 VSS.n17607 VSS.n17606 0.0121071
R21854 VSS.n17363 VSS.n17360 0.0121071
R21855 VSS.n18096 VSS.n18095 0.0121071
R21856 VSS.n18159 VSS.n18158 0.0121071
R21857 VSS.n18174 VSS.n215 0.0121071
R21858 VSS.n18581 VSS.n212 0.0121071
R21859 VSS.n18246 VSS.n18244 0.0121071
R21860 VSS.n18247 VSS.n18241 0.0121071
R21861 VSS.n18221 VSS.n18207 0.0121071
R21862 VSS.n18332 VSS.n18323 0.0121071
R21863 VSS.n18094 VSS.n277 0.0121071
R21864 VSS.n18160 VSS.n225 0.0121071
R21865 VSS.n9569 VSS.n9568 0.0121071
R21866 VSS.n9632 VSS.n9631 0.0121071
R21867 VSS.n9647 VSS.n9473 0.0121071
R21868 VSS.n9660 VSS.n9652 0.0121071
R21869 VSS.n9658 VSS.n9654 0.0121071
R21870 VSS.n9657 VSS.n9656 0.0121071
R21871 VSS.n9413 VSS.n9410 0.0121071
R21872 VSS.n9780 VSS.n9394 0.0121071
R21873 VSS.n9567 VSS.n9535 0.0121071
R21874 VSS.n9633 VSS.n9483 0.0121071
R21875 VSS.n16505 VSS.n16504 0.0121071
R21876 VSS.n16579 VSS.n16423 0.0121071
R21877 VSS.n16590 VSS.n16415 0.0121071
R21878 VSS.n16603 VSS.n16595 0.0121071
R21879 VSS.n16601 VSS.n16597 0.0121071
R21880 VSS.n16600 VSS.n16599 0.0121071
R21881 VSS.n16355 VSS.n16352 0.0121071
R21882 VSS.n16723 VSS.n16336 0.0121071
R21883 VSS.n16503 VSS.n16473 0.0121071
R21884 VSS.n16578 VSS.n16577 0.0121071
R21885 VSS.n1670 VSS.n1669 0.0121071
R21886 VSS.n1744 VSS.n1588 0.0121071
R21887 VSS.n15997 VSS.n1580 0.0121071
R21888 VSS.n16010 VSS.n16002 0.0121071
R21889 VSS.n16008 VSS.n16004 0.0121071
R21890 VSS.n16007 VSS.n16006 0.0121071
R21891 VSS.n1527 VSS.n1524 0.0121071
R21892 VSS.n16130 VSS.n1508 0.0121071
R21893 VSS.n1668 VSS.n1638 0.0121071
R21894 VSS.n1743 VSS.n1742 0.0121071
R21895 VSS.n1861 VSS.n1860 0.0121071
R21896 VSS.n1924 VSS.n1923 0.0121071
R21897 VSS.n1939 VSS.n1765 0.0121071
R21898 VSS.n2346 VSS.n1762 0.0121071
R21899 VSS.n2011 VSS.n2009 0.0121071
R21900 VSS.n2012 VSS.n2006 0.0121071
R21901 VSS.n1986 VSS.n1972 0.0121071
R21902 VSS.n2096 VSS.n2087 0.0121071
R21903 VSS.n1859 VSS.n1827 0.0121071
R21904 VSS.n1925 VSS.n1775 0.0121071
R21905 VSS.n3060 VSS.n3059 0.0121071
R21906 VSS.n3123 VSS.n3122 0.0121071
R21907 VSS.n3138 VSS.n2964 0.0121071
R21908 VSS.n3151 VSS.n3143 0.0121071
R21909 VSS.n3149 VSS.n3145 0.0121071
R21910 VSS.n3148 VSS.n3147 0.0121071
R21911 VSS.n2904 VSS.n2901 0.0121071
R21912 VSS.n3271 VSS.n2885 0.0121071
R21913 VSS.n3058 VSS.n3026 0.0121071
R21914 VSS.n3124 VSS.n2974 0.0121071
R21915 VSS.n3652 VSS.n3651 0.0121071
R21916 VSS.n3715 VSS.n3714 0.0121071
R21917 VSS.n3730 VSS.n3556 0.0121071
R21918 VSS.n3743 VSS.n3735 0.0121071
R21919 VSS.n3741 VSS.n3737 0.0121071
R21920 VSS.n3740 VSS.n3739 0.0121071
R21921 VSS.n3496 VSS.n3493 0.0121071
R21922 VSS.n3863 VSS.n3477 0.0121071
R21923 VSS.n3650 VSS.n3618 0.0121071
R21924 VSS.n3716 VSS.n3566 0.0121071
R21925 VSS.n4244 VSS.n4243 0.0121071
R21926 VSS.n4307 VSS.n4306 0.0121071
R21927 VSS.n4322 VSS.n4148 0.0121071
R21928 VSS.n4335 VSS.n4327 0.0121071
R21929 VSS.n4333 VSS.n4329 0.0121071
R21930 VSS.n4332 VSS.n4331 0.0121071
R21931 VSS.n4088 VSS.n4085 0.0121071
R21932 VSS.n4455 VSS.n4069 0.0121071
R21933 VSS.n4242 VSS.n4210 0.0121071
R21934 VSS.n4308 VSS.n4158 0.0121071
R21935 VSS.n4836 VSS.n4835 0.0121071
R21936 VSS.n4899 VSS.n4898 0.0121071
R21937 VSS.n4914 VSS.n4740 0.0121071
R21938 VSS.n4927 VSS.n4919 0.0121071
R21939 VSS.n4925 VSS.n4921 0.0121071
R21940 VSS.n4924 VSS.n4923 0.0121071
R21941 VSS.n4680 VSS.n4677 0.0121071
R21942 VSS.n5047 VSS.n4661 0.0121071
R21943 VSS.n4834 VSS.n4802 0.0121071
R21944 VSS.n4900 VSS.n4750 0.0121071
R21945 VSS.n2457 VSS.n2456 0.0121071
R21946 VSS.n2520 VSS.n2519 0.0121071
R21947 VSS.n2535 VSS.n2361 0.0121071
R21948 VSS.n5311 VSS.n2358 0.0121071
R21949 VSS.n2607 VSS.n2605 0.0121071
R21950 VSS.n2608 VSS.n2602 0.0121071
R21951 VSS.n2582 VSS.n2568 0.0121071
R21952 VSS.n2692 VSS.n2683 0.0121071
R21953 VSS.n2455 VSS.n2423 0.0121071
R21954 VSS.n2521 VSS.n2371 0.0121071
R21955 VSS.n5418 VSS.n5417 0.0121071
R21956 VSS.n5481 VSS.n5480 0.0121071
R21957 VSS.n5496 VSS.n5322 0.0121071
R21958 VSS.n5884 VSS.n5319 0.0121071
R21959 VSS.n5568 VSS.n5566 0.0121071
R21960 VSS.n5569 VSS.n5563 0.0121071
R21961 VSS.n5543 VSS.n5529 0.0121071
R21962 VSS.n5653 VSS.n5644 0.0121071
R21963 VSS.n5416 VSS.n5384 0.0121071
R21964 VSS.n5482 VSS.n5332 0.0121071
R21965 VSS.n5991 VSS.n5990 0.0121071
R21966 VSS.n6054 VSS.n6053 0.0121071
R21967 VSS.n6069 VSS.n5895 0.0121071
R21968 VSS.n6476 VSS.n5892 0.0121071
R21969 VSS.n6141 VSS.n6139 0.0121071
R21970 VSS.n6142 VSS.n6136 0.0121071
R21971 VSS.n6116 VSS.n6102 0.0121071
R21972 VSS.n6226 VSS.n6217 0.0121071
R21973 VSS.n5989 VSS.n5957 0.0121071
R21974 VSS.n6055 VSS.n5905 0.0121071
R21975 VSS.n7793 VSS.n7792 0.0121071
R21976 VSS.n7856 VSS.n7855 0.0121071
R21977 VSS.n7871 VSS.n7697 0.0121071
R21978 VSS.n7884 VSS.n7876 0.0121071
R21979 VSS.n7882 VSS.n7878 0.0121071
R21980 VSS.n7881 VSS.n7880 0.0121071
R21981 VSS.n7637 VSS.n7634 0.0121071
R21982 VSS.n8004 VSS.n7618 0.0121071
R21983 VSS.n7791 VSS.n7759 0.0121071
R21984 VSS.n7857 VSS.n7707 0.0121071
R21985 VSS.n8385 VSS.n8384 0.0121071
R21986 VSS.n8448 VSS.n8447 0.0121071
R21987 VSS.n8463 VSS.n8289 0.0121071
R21988 VSS.n8476 VSS.n8468 0.0121071
R21989 VSS.n8474 VSS.n8470 0.0121071
R21990 VSS.n8473 VSS.n8472 0.0121071
R21991 VSS.n8229 VSS.n8226 0.0121071
R21992 VSS.n8596 VSS.n8210 0.0121071
R21993 VSS.n8383 VSS.n8351 0.0121071
R21994 VSS.n8449 VSS.n8299 0.0121071
R21995 VSS.n8977 VSS.n8976 0.0121071
R21996 VSS.n9040 VSS.n9039 0.0121071
R21997 VSS.n9055 VSS.n8881 0.0121071
R21998 VSS.n9068 VSS.n9060 0.0121071
R21999 VSS.n9066 VSS.n9062 0.0121071
R22000 VSS.n9065 VSS.n9064 0.0121071
R22001 VSS.n8821 VSS.n8818 0.0121071
R22002 VSS.n9188 VSS.n8802 0.0121071
R22003 VSS.n8975 VSS.n8943 0.0121071
R22004 VSS.n9041 VSS.n8891 0.0121071
R22005 VSS.n10161 VSS.n10160 0.0121071
R22006 VSS.n10224 VSS.n10223 0.0121071
R22007 VSS.n10239 VSS.n10065 0.0121071
R22008 VSS.n10252 VSS.n10244 0.0121071
R22009 VSS.n10250 VSS.n10246 0.0121071
R22010 VSS.n10249 VSS.n10248 0.0121071
R22011 VSS.n10005 VSS.n10002 0.0121071
R22012 VSS.n10372 VSS.n9986 0.0121071
R22013 VSS.n10159 VSS.n10127 0.0121071
R22014 VSS.n10225 VSS.n10075 0.0121071
R22015 VSS.n10753 VSS.n10752 0.0121071
R22016 VSS.n10816 VSS.n10815 0.0121071
R22017 VSS.n10831 VSS.n10657 0.0121071
R22018 VSS.n10844 VSS.n10836 0.0121071
R22019 VSS.n10842 VSS.n10838 0.0121071
R22020 VSS.n10841 VSS.n10840 0.0121071
R22021 VSS.n10597 VSS.n10594 0.0121071
R22022 VSS.n10964 VSS.n10578 0.0121071
R22023 VSS.n10751 VSS.n10719 0.0121071
R22024 VSS.n10817 VSS.n10667 0.0121071
R22025 VSS.n11345 VSS.n11344 0.0121071
R22026 VSS.n11408 VSS.n11407 0.0121071
R22027 VSS.n11423 VSS.n11249 0.0121071
R22028 VSS.n11436 VSS.n11428 0.0121071
R22029 VSS.n11434 VSS.n11430 0.0121071
R22030 VSS.n11433 VSS.n11432 0.0121071
R22031 VSS.n11189 VSS.n11186 0.0121071
R22032 VSS.n11556 VSS.n11170 0.0121071
R22033 VSS.n11343 VSS.n11311 0.0121071
R22034 VSS.n11409 VSS.n11259 0.0121071
R22035 VSS.n11937 VSS.n11936 0.0121071
R22036 VSS.n12000 VSS.n11999 0.0121071
R22037 VSS.n12015 VSS.n11841 0.0121071
R22038 VSS.n12028 VSS.n12020 0.0121071
R22039 VSS.n12026 VSS.n12022 0.0121071
R22040 VSS.n12025 VSS.n12024 0.0121071
R22041 VSS.n11781 VSS.n11778 0.0121071
R22042 VSS.n12148 VSS.n11762 0.0121071
R22043 VSS.n11935 VSS.n11903 0.0121071
R22044 VSS.n12001 VSS.n11851 0.0121071
R22045 VSS.n12529 VSS.n12528 0.0121071
R22046 VSS.n12592 VSS.n12591 0.0121071
R22047 VSS.n12607 VSS.n12433 0.0121071
R22048 VSS.n12620 VSS.n12612 0.0121071
R22049 VSS.n12618 VSS.n12614 0.0121071
R22050 VSS.n12617 VSS.n12616 0.0121071
R22051 VSS.n12373 VSS.n12370 0.0121071
R22052 VSS.n12740 VSS.n12354 0.0121071
R22053 VSS.n12527 VSS.n12495 0.0121071
R22054 VSS.n12593 VSS.n12443 0.0121071
R22055 VSS.n13121 VSS.n13120 0.0121071
R22056 VSS.n13184 VSS.n13183 0.0121071
R22057 VSS.n13199 VSS.n13025 0.0121071
R22058 VSS.n13212 VSS.n13204 0.0121071
R22059 VSS.n13210 VSS.n13206 0.0121071
R22060 VSS.n13209 VSS.n13208 0.0121071
R22061 VSS.n12965 VSS.n12962 0.0121071
R22062 VSS.n13332 VSS.n12946 0.0121071
R22063 VSS.n13119 VSS.n13087 0.0121071
R22064 VSS.n13185 VSS.n13035 0.0121071
R22065 VSS.n13713 VSS.n13712 0.0121071
R22066 VSS.n13776 VSS.n13775 0.0121071
R22067 VSS.n13791 VSS.n13617 0.0121071
R22068 VSS.n13804 VSS.n13796 0.0121071
R22069 VSS.n13802 VSS.n13798 0.0121071
R22070 VSS.n13801 VSS.n13800 0.0121071
R22071 VSS.n13557 VSS.n13554 0.0121071
R22072 VSS.n13924 VSS.n13538 0.0121071
R22073 VSS.n13711 VSS.n13679 0.0121071
R22074 VSS.n13777 VSS.n13627 0.0121071
R22075 VSS.n14305 VSS.n14304 0.0121071
R22076 VSS.n14368 VSS.n14367 0.0121071
R22077 VSS.n14383 VSS.n14209 0.0121071
R22078 VSS.n14396 VSS.n14388 0.0121071
R22079 VSS.n14394 VSS.n14390 0.0121071
R22080 VSS.n14393 VSS.n14392 0.0121071
R22081 VSS.n14149 VSS.n14146 0.0121071
R22082 VSS.n14516 VSS.n14130 0.0121071
R22083 VSS.n14303 VSS.n14271 0.0121071
R22084 VSS.n14369 VSS.n14219 0.0121071
R22085 VSS.n14897 VSS.n14896 0.0121071
R22086 VSS.n14960 VSS.n14959 0.0121071
R22087 VSS.n14975 VSS.n14801 0.0121071
R22088 VSS.n14988 VSS.n14980 0.0121071
R22089 VSS.n14986 VSS.n14982 0.0121071
R22090 VSS.n14985 VSS.n14984 0.0121071
R22091 VSS.n14741 VSS.n14738 0.0121071
R22092 VSS.n15108 VSS.n14722 0.0121071
R22093 VSS.n14895 VSS.n14863 0.0121071
R22094 VSS.n14961 VSS.n14811 0.0121071
R22095 VSS.n15489 VSS.n15488 0.0121071
R22096 VSS.n15552 VSS.n15551 0.0121071
R22097 VSS.n15567 VSS.n15393 0.0121071
R22098 VSS.n15580 VSS.n15572 0.0121071
R22099 VSS.n15578 VSS.n15574 0.0121071
R22100 VSS.n15577 VSS.n15576 0.0121071
R22101 VSS.n15333 VSS.n15330 0.0121071
R22102 VSS.n15700 VSS.n15314 0.0121071
R22103 VSS.n15487 VSS.n15455 0.0121071
R22104 VSS.n15553 VSS.n15403 0.0121071
R22105 VSS.n6597 VSS.n6596 0.0121071
R22106 VSS.n6660 VSS.n6659 0.0121071
R22107 VSS.n6675 VSS.n6501 0.0121071
R22108 VSS.n15964 VSS.n6498 0.0121071
R22109 VSS.n6747 VSS.n6745 0.0121071
R22110 VSS.n6748 VSS.n6742 0.0121071
R22111 VSS.n6722 VSS.n6708 0.0121071
R22112 VSS.n6832 VSS.n6823 0.0121071
R22113 VSS.n6595 VSS.n6563 0.0121071
R22114 VSS.n6661 VSS.n6511 0.0121071
R22115 VSS.n7194 VSS.n7193 0.0121071
R22116 VSS.n7268 VSS.n7112 0.0121071
R22117 VSS.n7279 VSS.n7104 0.0121071
R22118 VSS.n7292 VSS.n7284 0.0121071
R22119 VSS.n7290 VSS.n7286 0.0121071
R22120 VSS.n7289 VSS.n7288 0.0121071
R22121 VSS.n7044 VSS.n7041 0.0121071
R22122 VSS.n7412 VSS.n7025 0.0121071
R22123 VSS.n7192 VSS.n7162 0.0121071
R22124 VSS.n7267 VSS.n7266 0.0121071
R22125 VSS.n346 VSS.n297 0.0121071
R22126 VSS.n411 VSS.n410 0.0121071
R22127 VSS.n18591 VSS.n195 0.0121071
R22128 VSS.n18604 VSS.n18596 0.0121071
R22129 VSS.n18602 VSS.n18598 0.0121071
R22130 VSS.n18601 VSS.n18600 0.0121071
R22131 VSS.n142 VSS.n139 0.0121071
R22132 VSS.n18724 VSS.n123 0.0121071
R22133 VSS.n352 VSS.n295 0.0121071
R22134 VSS.n409 VSS.n324 0.0121071
R22135 VSS.n877 VSS.n876 0.0121071
R22136 VSS.n570 VSS.n568 0.0121071
R22137 VSS.n571 VSS.n567 0.0121071
R22138 VSS.n542 VSS.n528 0.0121071
R22139 VSS.n655 VSS.n646 0.0121071
R22140 VSS.n918 VSS.n461 0.0121071
R22141 VSS.n965 VSS.n964 0.0121071
R22142 VSS.n1314 VSS.n1305 0.0121071
R22143 VSS.n1229 VSS.n1228 0.0112143
R22144 VSS.n1233 VSS.n1165 0.0112143
R22145 VSS.n1205 VSS.n1189 0.0112143
R22146 VSS.n1232 VSS.n1163 0.0112143
R22147 VSS.n967 VSS.n966 0.0112143
R22148 VSS.n17012 VSS.n17011 0.0112143
R22149 VSS.n17025 VSS.n17024 0.0112143
R22150 VSS.n17088 VSS.n17087 0.0112143
R22151 VSS.n1148 VSS.n1147 0.0112143
R22152 VSS.n1070 VSS.n1056 0.0112143
R22153 VSS.n17181 VSS.n17180 0.0112143
R22154 VSS.n17203 VSS.n17202 0.0112143
R22155 VSS.n17232 VSS.n16885 0.0112143
R22156 VSS.n17249 VSS.n16863 0.0112143
R22157 VSS.n17231 VSS.n17230 0.0112143
R22158 VSS.n17023 VSS.n16992 0.0112143
R22159 VSS.n17604 VSS.n17603 0.0112143
R22160 VSS.n17617 VSS.n17616 0.0112143
R22161 VSS.n17680 VSS.n17679 0.0112143
R22162 VSS.n17582 VSS.n17438 0.0112143
R22163 VSS.n17585 VSS.n17432 0.0112143
R22164 VSS.n17773 VSS.n17772 0.0112143
R22165 VSS.n17795 VSS.n17794 0.0112143
R22166 VSS.n17824 VSS.n17299 0.0112143
R22167 VSS.n17841 VSS.n17277 0.0112143
R22168 VSS.n17823 VSS.n17822 0.0112143
R22169 VSS.n17615 VSS.n17406 0.0112143
R22170 VSS.n18159 VSS.n230 0.0112143
R22171 VSS.n18246 VSS.n18245 0.0112143
R22172 VSS.n18250 VSS.n18182 0.0112143
R22173 VSS.n18222 VSS.n18206 0.0112143
R22174 VSS.n18249 VSS.n18180 0.0112143
R22175 VSS.n18378 VSS.n18345 0.0112143
R22176 VSS.n18408 VSS.n18407 0.0112143
R22177 VSS.n18446 VSS.n18418 0.0112143
R22178 VSS.n18434 VSS.n18433 0.0112143
R22179 VSS.n18445 VSS.n18416 0.0112143
R22180 VSS.n18162 VSS.n224 0.0112143
R22181 VSS.n9632 VSS.n9488 0.0112143
R22182 VSS.n9654 VSS.n9653 0.0112143
R22183 VSS.n9667 VSS.n9666 0.0112143
R22184 VSS.n9730 VSS.n9729 0.0112143
R22185 VSS.n9665 VSS.n9456 0.0112143
R22186 VSS.n9823 VSS.n9822 0.0112143
R22187 VSS.n9845 VSS.n9844 0.0112143
R22188 VSS.n9874 VSS.n9349 0.0112143
R22189 VSS.n9892 VSS.n9328 0.0112143
R22190 VSS.n9873 VSS.n9872 0.0112143
R22191 VSS.n9635 VSS.n9482 0.0112143
R22192 VSS.n16580 VSS.n16579 0.0112143
R22193 VSS.n16597 VSS.n16596 0.0112143
R22194 VSS.n16610 VSS.n16609 0.0112143
R22195 VSS.n16673 VSS.n16672 0.0112143
R22196 VSS.n16608 VSS.n16398 0.0112143
R22197 VSS.n16766 VSS.n16765 0.0112143
R22198 VSS.n16788 VSS.n16787 0.0112143
R22199 VSS.n16817 VSS.n16291 0.0112143
R22200 VSS.n16835 VSS.n16270 0.0112143
R22201 VSS.n16816 VSS.n16815 0.0112143
R22202 VSS.n16430 VSS.n16427 0.0112143
R22203 VSS.n1745 VSS.n1744 0.0112143
R22204 VSS.n16004 VSS.n16003 0.0112143
R22205 VSS.n16017 VSS.n16016 0.0112143
R22206 VSS.n16080 VSS.n16079 0.0112143
R22207 VSS.n16015 VSS.n1570 0.0112143
R22208 VSS.n16173 VSS.n16172 0.0112143
R22209 VSS.n16195 VSS.n16194 0.0112143
R22210 VSS.n16224 VSS.n1463 0.0112143
R22211 VSS.n16242 VSS.n1442 0.0112143
R22212 VSS.n16223 VSS.n16222 0.0112143
R22213 VSS.n1595 VSS.n1592 0.0112143
R22214 VSS.n1924 VSS.n1780 0.0112143
R22215 VSS.n2011 VSS.n2010 0.0112143
R22216 VSS.n2015 VSS.n1947 0.0112143
R22217 VSS.n1987 VSS.n1971 0.0112143
R22218 VSS.n2014 VSS.n1945 0.0112143
R22219 VSS.n2141 VSS.n2140 0.0112143
R22220 VSS.n2184 VSS.n2155 0.0112143
R22221 VSS.n2243 VSS.n2242 0.0112143
R22222 VSS.n2224 VSS.n2200 0.0112143
R22223 VSS.n2244 VSS.n2161 0.0112143
R22224 VSS.n1927 VSS.n1774 0.0112143
R22225 VSS.n3123 VSS.n2979 0.0112143
R22226 VSS.n3145 VSS.n3144 0.0112143
R22227 VSS.n3158 VSS.n3157 0.0112143
R22228 VSS.n3221 VSS.n3220 0.0112143
R22229 VSS.n3156 VSS.n2947 0.0112143
R22230 VSS.n3314 VSS.n3313 0.0112143
R22231 VSS.n3336 VSS.n3335 0.0112143
R22232 VSS.n3365 VSS.n2840 0.0112143
R22233 VSS.n3383 VSS.n2819 0.0112143
R22234 VSS.n3364 VSS.n3363 0.0112143
R22235 VSS.n3126 VSS.n2973 0.0112143
R22236 VSS.n3715 VSS.n3571 0.0112143
R22237 VSS.n3737 VSS.n3736 0.0112143
R22238 VSS.n3750 VSS.n3749 0.0112143
R22239 VSS.n3813 VSS.n3812 0.0112143
R22240 VSS.n3748 VSS.n3539 0.0112143
R22241 VSS.n3906 VSS.n3905 0.0112143
R22242 VSS.n3928 VSS.n3927 0.0112143
R22243 VSS.n3957 VSS.n3432 0.0112143
R22244 VSS.n3975 VSS.n3411 0.0112143
R22245 VSS.n3956 VSS.n3955 0.0112143
R22246 VSS.n3718 VSS.n3565 0.0112143
R22247 VSS.n4307 VSS.n4163 0.0112143
R22248 VSS.n4329 VSS.n4328 0.0112143
R22249 VSS.n4342 VSS.n4341 0.0112143
R22250 VSS.n4405 VSS.n4404 0.0112143
R22251 VSS.n4340 VSS.n4131 0.0112143
R22252 VSS.n4498 VSS.n4497 0.0112143
R22253 VSS.n4520 VSS.n4519 0.0112143
R22254 VSS.n4549 VSS.n4024 0.0112143
R22255 VSS.n4567 VSS.n4003 0.0112143
R22256 VSS.n4548 VSS.n4547 0.0112143
R22257 VSS.n4310 VSS.n4157 0.0112143
R22258 VSS.n4899 VSS.n4755 0.0112143
R22259 VSS.n4921 VSS.n4920 0.0112143
R22260 VSS.n4934 VSS.n4933 0.0112143
R22261 VSS.n4997 VSS.n4996 0.0112143
R22262 VSS.n4932 VSS.n4723 0.0112143
R22263 VSS.n5090 VSS.n5089 0.0112143
R22264 VSS.n5112 VSS.n5111 0.0112143
R22265 VSS.n5141 VSS.n4616 0.0112143
R22266 VSS.n5159 VSS.n4595 0.0112143
R22267 VSS.n5140 VSS.n5139 0.0112143
R22268 VSS.n4902 VSS.n4749 0.0112143
R22269 VSS.n2520 VSS.n2376 0.0112143
R22270 VSS.n2607 VSS.n2606 0.0112143
R22271 VSS.n2611 VSS.n2543 0.0112143
R22272 VSS.n2583 VSS.n2567 0.0112143
R22273 VSS.n2610 VSS.n2541 0.0112143
R22274 VSS.n2737 VSS.n2736 0.0112143
R22275 VSS.n2780 VSS.n2751 0.0112143
R22276 VSS.n5208 VSS.n5207 0.0112143
R22277 VSS.n5189 VSS.n2796 0.0112143
R22278 VSS.n5209 VSS.n2757 0.0112143
R22279 VSS.n2523 VSS.n2370 0.0112143
R22280 VSS.n5481 VSS.n5337 0.0112143
R22281 VSS.n5568 VSS.n5567 0.0112143
R22282 VSS.n5572 VSS.n5504 0.0112143
R22283 VSS.n5544 VSS.n5528 0.0112143
R22284 VSS.n5571 VSS.n5502 0.0112143
R22285 VSS.n5698 VSS.n5697 0.0112143
R22286 VSS.n5754 VSS.n5712 0.0112143
R22287 VSS.n5781 VSS.n5780 0.0112143
R22288 VSS.n5734 VSS.n4 0.0112143
R22289 VSS.n5782 VSS.n5718 0.0112143
R22290 VSS.n5484 VSS.n5331 0.0112143
R22291 VSS.n6054 VSS.n5910 0.0112143
R22292 VSS.n6141 VSS.n6140 0.0112143
R22293 VSS.n6145 VSS.n6077 0.0112143
R22294 VSS.n6117 VSS.n6101 0.0112143
R22295 VSS.n6144 VSS.n6075 0.0112143
R22296 VSS.n6271 VSS.n6270 0.0112143
R22297 VSS.n6314 VSS.n6285 0.0112143
R22298 VSS.n6373 VSS.n6372 0.0112143
R22299 VSS.n6354 VSS.n6330 0.0112143
R22300 VSS.n6374 VSS.n6291 0.0112143
R22301 VSS.n6057 VSS.n5904 0.0112143
R22302 VSS.n7856 VSS.n7712 0.0112143
R22303 VSS.n7878 VSS.n7877 0.0112143
R22304 VSS.n7891 VSS.n7890 0.0112143
R22305 VSS.n7954 VSS.n7953 0.0112143
R22306 VSS.n7889 VSS.n7680 0.0112143
R22307 VSS.n8047 VSS.n8046 0.0112143
R22308 VSS.n8069 VSS.n8068 0.0112143
R22309 VSS.n8098 VSS.n7573 0.0112143
R22310 VSS.n8116 VSS.n7552 0.0112143
R22311 VSS.n8097 VSS.n8096 0.0112143
R22312 VSS.n7859 VSS.n7706 0.0112143
R22313 VSS.n8448 VSS.n8304 0.0112143
R22314 VSS.n8470 VSS.n8469 0.0112143
R22315 VSS.n8483 VSS.n8482 0.0112143
R22316 VSS.n8546 VSS.n8545 0.0112143
R22317 VSS.n8481 VSS.n8272 0.0112143
R22318 VSS.n8639 VSS.n8638 0.0112143
R22319 VSS.n8661 VSS.n8660 0.0112143
R22320 VSS.n8690 VSS.n8165 0.0112143
R22321 VSS.n8708 VSS.n8144 0.0112143
R22322 VSS.n8689 VSS.n8688 0.0112143
R22323 VSS.n8451 VSS.n8298 0.0112143
R22324 VSS.n9040 VSS.n8896 0.0112143
R22325 VSS.n9062 VSS.n9061 0.0112143
R22326 VSS.n9075 VSS.n9074 0.0112143
R22327 VSS.n9138 VSS.n9137 0.0112143
R22328 VSS.n9073 VSS.n8864 0.0112143
R22329 VSS.n9231 VSS.n9230 0.0112143
R22330 VSS.n9253 VSS.n9252 0.0112143
R22331 VSS.n9282 VSS.n8757 0.0112143
R22332 VSS.n9300 VSS.n8736 0.0112143
R22333 VSS.n9281 VSS.n9280 0.0112143
R22334 VSS.n9043 VSS.n8890 0.0112143
R22335 VSS.n10224 VSS.n10080 0.0112143
R22336 VSS.n10246 VSS.n10245 0.0112143
R22337 VSS.n10259 VSS.n10258 0.0112143
R22338 VSS.n10322 VSS.n10321 0.0112143
R22339 VSS.n10257 VSS.n10048 0.0112143
R22340 VSS.n10415 VSS.n10414 0.0112143
R22341 VSS.n10437 VSS.n10436 0.0112143
R22342 VSS.n10466 VSS.n9941 0.0112143
R22343 VSS.n10484 VSS.n9920 0.0112143
R22344 VSS.n10465 VSS.n10464 0.0112143
R22345 VSS.n10227 VSS.n10074 0.0112143
R22346 VSS.n10816 VSS.n10672 0.0112143
R22347 VSS.n10838 VSS.n10837 0.0112143
R22348 VSS.n10851 VSS.n10850 0.0112143
R22349 VSS.n10914 VSS.n10913 0.0112143
R22350 VSS.n10849 VSS.n10640 0.0112143
R22351 VSS.n11007 VSS.n11006 0.0112143
R22352 VSS.n11029 VSS.n11028 0.0112143
R22353 VSS.n11058 VSS.n10533 0.0112143
R22354 VSS.n11076 VSS.n10512 0.0112143
R22355 VSS.n11057 VSS.n11056 0.0112143
R22356 VSS.n10819 VSS.n10666 0.0112143
R22357 VSS.n11408 VSS.n11264 0.0112143
R22358 VSS.n11430 VSS.n11429 0.0112143
R22359 VSS.n11443 VSS.n11442 0.0112143
R22360 VSS.n11506 VSS.n11505 0.0112143
R22361 VSS.n11441 VSS.n11232 0.0112143
R22362 VSS.n11599 VSS.n11598 0.0112143
R22363 VSS.n11621 VSS.n11620 0.0112143
R22364 VSS.n11650 VSS.n11125 0.0112143
R22365 VSS.n11668 VSS.n11104 0.0112143
R22366 VSS.n11649 VSS.n11648 0.0112143
R22367 VSS.n11411 VSS.n11258 0.0112143
R22368 VSS.n12000 VSS.n11856 0.0112143
R22369 VSS.n12022 VSS.n12021 0.0112143
R22370 VSS.n12035 VSS.n12034 0.0112143
R22371 VSS.n12098 VSS.n12097 0.0112143
R22372 VSS.n12033 VSS.n11824 0.0112143
R22373 VSS.n12191 VSS.n12190 0.0112143
R22374 VSS.n12213 VSS.n12212 0.0112143
R22375 VSS.n12242 VSS.n11717 0.0112143
R22376 VSS.n12260 VSS.n11696 0.0112143
R22377 VSS.n12241 VSS.n12240 0.0112143
R22378 VSS.n12003 VSS.n11850 0.0112143
R22379 VSS.n12592 VSS.n12448 0.0112143
R22380 VSS.n12614 VSS.n12613 0.0112143
R22381 VSS.n12627 VSS.n12626 0.0112143
R22382 VSS.n12690 VSS.n12689 0.0112143
R22383 VSS.n12625 VSS.n12416 0.0112143
R22384 VSS.n12783 VSS.n12782 0.0112143
R22385 VSS.n12805 VSS.n12804 0.0112143
R22386 VSS.n12834 VSS.n12309 0.0112143
R22387 VSS.n12852 VSS.n12288 0.0112143
R22388 VSS.n12833 VSS.n12832 0.0112143
R22389 VSS.n12595 VSS.n12442 0.0112143
R22390 VSS.n13184 VSS.n13040 0.0112143
R22391 VSS.n13206 VSS.n13205 0.0112143
R22392 VSS.n13219 VSS.n13218 0.0112143
R22393 VSS.n13282 VSS.n13281 0.0112143
R22394 VSS.n13217 VSS.n13008 0.0112143
R22395 VSS.n13375 VSS.n13374 0.0112143
R22396 VSS.n13397 VSS.n13396 0.0112143
R22397 VSS.n13426 VSS.n12901 0.0112143
R22398 VSS.n13444 VSS.n12880 0.0112143
R22399 VSS.n13425 VSS.n13424 0.0112143
R22400 VSS.n13187 VSS.n13034 0.0112143
R22401 VSS.n13776 VSS.n13632 0.0112143
R22402 VSS.n13798 VSS.n13797 0.0112143
R22403 VSS.n13811 VSS.n13810 0.0112143
R22404 VSS.n13874 VSS.n13873 0.0112143
R22405 VSS.n13809 VSS.n13600 0.0112143
R22406 VSS.n13967 VSS.n13966 0.0112143
R22407 VSS.n13989 VSS.n13988 0.0112143
R22408 VSS.n14018 VSS.n13493 0.0112143
R22409 VSS.n14036 VSS.n13472 0.0112143
R22410 VSS.n14017 VSS.n14016 0.0112143
R22411 VSS.n13779 VSS.n13626 0.0112143
R22412 VSS.n14368 VSS.n14224 0.0112143
R22413 VSS.n14390 VSS.n14389 0.0112143
R22414 VSS.n14403 VSS.n14402 0.0112143
R22415 VSS.n14466 VSS.n14465 0.0112143
R22416 VSS.n14401 VSS.n14192 0.0112143
R22417 VSS.n14559 VSS.n14558 0.0112143
R22418 VSS.n14581 VSS.n14580 0.0112143
R22419 VSS.n14610 VSS.n14085 0.0112143
R22420 VSS.n14628 VSS.n14064 0.0112143
R22421 VSS.n14609 VSS.n14608 0.0112143
R22422 VSS.n14371 VSS.n14218 0.0112143
R22423 VSS.n14960 VSS.n14816 0.0112143
R22424 VSS.n14982 VSS.n14981 0.0112143
R22425 VSS.n14995 VSS.n14994 0.0112143
R22426 VSS.n15058 VSS.n15057 0.0112143
R22427 VSS.n14993 VSS.n14784 0.0112143
R22428 VSS.n15151 VSS.n15150 0.0112143
R22429 VSS.n15173 VSS.n15172 0.0112143
R22430 VSS.n15202 VSS.n14677 0.0112143
R22431 VSS.n15220 VSS.n14656 0.0112143
R22432 VSS.n15201 VSS.n15200 0.0112143
R22433 VSS.n14963 VSS.n14810 0.0112143
R22434 VSS.n15552 VSS.n15408 0.0112143
R22435 VSS.n15574 VSS.n15573 0.0112143
R22436 VSS.n15587 VSS.n15586 0.0112143
R22437 VSS.n15650 VSS.n15649 0.0112143
R22438 VSS.n15585 VSS.n15376 0.0112143
R22439 VSS.n15743 VSS.n15742 0.0112143
R22440 VSS.n15765 VSS.n15764 0.0112143
R22441 VSS.n15794 VSS.n15269 0.0112143
R22442 VSS.n15812 VSS.n15248 0.0112143
R22443 VSS.n15793 VSS.n15792 0.0112143
R22444 VSS.n15555 VSS.n15402 0.0112143
R22445 VSS.n6660 VSS.n6516 0.0112143
R22446 VSS.n6747 VSS.n6746 0.0112143
R22447 VSS.n6751 VSS.n6683 0.0112143
R22448 VSS.n6723 VSS.n6707 0.0112143
R22449 VSS.n6750 VSS.n6681 0.0112143
R22450 VSS.n6877 VSS.n6876 0.0112143
R22451 VSS.n6920 VSS.n6891 0.0112143
R22452 VSS.n15861 VSS.n15860 0.0112143
R22453 VSS.n15842 VSS.n6936 0.0112143
R22454 VSS.n15862 VSS.n6897 0.0112143
R22455 VSS.n6663 VSS.n6510 0.0112143
R22456 VSS.n7269 VSS.n7268 0.0112143
R22457 VSS.n7286 VSS.n7285 0.0112143
R22458 VSS.n7299 VSS.n7298 0.0112143
R22459 VSS.n7362 VSS.n7361 0.0112143
R22460 VSS.n7297 VSS.n7087 0.0112143
R22461 VSS.n7455 VSS.n7454 0.0112143
R22462 VSS.n7477 VSS.n7476 0.0112143
R22463 VSS.n7506 VSS.n6980 0.0112143
R22464 VSS.n7524 VSS.n6959 0.0112143
R22465 VSS.n7505 VSS.n7504 0.0112143
R22466 VSS.n7119 VSS.n7116 0.0112143
R22467 VSS.n410 VSS.n325 0.0112143
R22468 VSS.n18598 VSS.n18597 0.0112143
R22469 VSS.n18611 VSS.n18610 0.0112143
R22470 VSS.n18674 VSS.n18673 0.0112143
R22471 VSS.n18609 VSS.n185 0.0112143
R22472 VSS.n18767 VSS.n18766 0.0112143
R22473 VSS.n18789 VSS.n18788 0.0112143
R22474 VSS.n18818 VSS.n78 0.0112143
R22475 VSS.n18836 VSS.n57 0.0112143
R22476 VSS.n18817 VSS.n18816 0.0112143
R22477 VSS.n326 VSS.n323 0.0112143
R22478 VSS.n570 VSS.n569 0.0112143
R22479 VSS.n574 VSS.n503 0.0112143
R22480 VSS.n543 VSS.n527 0.0112143
R22481 VSS.n573 VSS.n501 0.0112143
R22482 VSS.n700 VSS.n699 0.0112143
R22483 VSS.n752 VSS.n714 0.0112143
R22484 VSS.n775 VSS.n774 0.0112143
R22485 VSS.n18865 VSS.n49 0.0112143
R22486 VSS.n776 VSS.n720 0.0112143
R22487 VSS.n889 VSS.n489 0.0112143
R22488 VSS.n1359 VSS.n1358 0.0112143
R22489 VSS.n1402 VSS.n1373 0.0112143
R22490 VSS.n17889 VSS.n17888 0.0112143
R22491 VSS.n17870 VSS.n1418 0.0112143
R22492 VSS.n17890 VSS.n1379 0.0112143
R22493 VSS.n1233 VSS.n1223 0.0103214
R22494 VSS.n17985 VSS.n17984 0.0103214
R22495 VSS.n17978 VSS.n1171 0.0103214
R22496 VSS.n1260 VSS.n1180 0.0103214
R22497 VSS.n1282 VSS.n1281 0.0103214
R22498 VSS.n1232 VSS.n1231 0.0103214
R22499 VSS.n17979 VSS.n1169 0.0103214
R22500 VSS.n17975 VSS.n1174 0.0103214
R22501 VSS.n17966 VSS.n1183 0.0103214
R22502 VSS.n1264 VSS.n1186 0.0103214
R22503 VSS.n915 VSS.n914 0.0103214
R22504 VSS.n1001 VSS.n469 0.0103214
R22505 VSS.n944 VSS.n479 0.0103214
R22506 VSS.n984 VSS.n983 0.0103214
R22507 VSS.n890 VSS.n488 0.0103214
R22508 VSS.n962 VSS.n961 0.0103214
R22509 VSS.n17025 VSS.n16991 0.0103214
R22510 VSS.n16994 VSS.n16993 0.0103214
R22511 VSS.n17045 VSS.n16978 0.0103214
R22512 VSS.n17066 VSS.n16957 0.0103214
R22513 VSS.n17099 VSS.n17098 0.0103214
R22514 VSS.n1096 VSS.n1095 0.0103214
R22515 VSS.n18027 VSS.n1036 0.0103214
R22516 VSS.n1125 VSS.n1046 0.0103214
R22517 VSS.n18010 VSS.n18009 0.0103214
R22518 VSS.n1071 VSS.n1055 0.0103214
R22519 VSS.n1143 VSS.n1142 0.0103214
R22520 VSS.n18028 VSS.n1034 0.0103214
R22521 VSS.n1047 VSS.n1044 0.0103214
R22522 VSS.n18015 VSS.n1049 0.0103214
R22523 VSS.n1144 VSS.n1070 0.0103214
R22524 VSS.n17149 VSS.n16923 0.0103214
R22525 VSS.n17153 VSS.n16921 0.0103214
R22526 VSS.n17155 VSS.n16919 0.0103214
R22527 VSS.n17148 VSS.n16925 0.0103214
R22528 VSS.n17157 VSS.n17156 0.0103214
R22529 VSS.n17013 VSS.n16992 0.0103214
R22530 VSS.n17044 VSS.n17043 0.0103214
R22531 VSS.n17039 VSS.n16967 0.0103214
R22532 VSS.n17067 VSS.n16959 0.0103214
R22533 VSS.n17075 VSS.n17074 0.0103214
R22534 VSS.n17617 VSS.n17405 0.0103214
R22535 VSS.n17408 VSS.n17407 0.0103214
R22536 VSS.n17637 VSS.n17392 0.0103214
R22537 VSS.n17658 VSS.n17371 0.0103214
R22538 VSS.n17691 VSS.n17690 0.0103214
R22539 VSS.n17506 VSS.n17505 0.0103214
R22540 VSS.n17475 VSS.n17468 0.0103214
R22541 VSS.n17567 VSS.n17566 0.0103214
R22542 VSS.n17574 VSS.n17573 0.0103214
R22543 VSS.n17587 VSS.n17430 0.0103214
R22544 VSS.n17586 VSS.n17431 0.0103214
R22545 VSS.n17474 VSS.n17469 0.0103214
R22546 VSS.n17548 VSS.n17465 0.0103214
R22547 VSS.n17568 VSS.n17445 0.0103214
R22548 VSS.n17585 VSS.n17584 0.0103214
R22549 VSS.n17741 VSS.n17337 0.0103214
R22550 VSS.n17745 VSS.n17335 0.0103214
R22551 VSS.n17747 VSS.n17333 0.0103214
R22552 VSS.n17740 VSS.n17339 0.0103214
R22553 VSS.n17749 VSS.n17748 0.0103214
R22554 VSS.n17605 VSS.n17406 0.0103214
R22555 VSS.n17636 VSS.n17635 0.0103214
R22556 VSS.n17631 VSS.n17381 0.0103214
R22557 VSS.n17659 VSS.n17373 0.0103214
R22558 VSS.n17667 VSS.n17666 0.0103214
R22559 VSS.n18083 VSS.n18082 0.0103214
R22560 VSS.n267 VSS.n260 0.0103214
R22561 VSS.n18144 VSS.n18143 0.0103214
R22562 VSS.n18151 VSS.n18150 0.0103214
R22563 VSS.n18164 VSS.n222 0.0103214
R22564 VSS.n18163 VSS.n223 0.0103214
R22565 VSS.n18250 VSS.n18240 0.0103214
R22566 VSS.n18574 VSS.n18573 0.0103214
R22567 VSS.n18567 VSS.n18188 0.0103214
R22568 VSS.n18277 VSS.n18197 0.0103214
R22569 VSS.n18299 VSS.n18298 0.0103214
R22570 VSS.n18249 VSS.n18248 0.0103214
R22571 VSS.n18568 VSS.n18186 0.0103214
R22572 VSS.n18564 VSS.n18191 0.0103214
R22573 VSS.n18555 VSS.n18200 0.0103214
R22574 VSS.n18281 VSS.n18203 0.0103214
R22575 VSS.n18526 VSS.n18525 0.0103214
R22576 VSS.n18363 VSS.n18339 0.0103214
R22577 VSS.n18517 VSS.n18516 0.0103214
R22578 VSS.n18524 VSS.n18315 0.0103214
R22579 VSS.n18515 VSS.n18338 0.0103214
R22580 VSS.n266 VSS.n261 0.0103214
R22581 VSS.n18125 VSS.n257 0.0103214
R22582 VSS.n18145 VSS.n237 0.0103214
R22583 VSS.n18162 VSS.n18161 0.0103214
R22584 VSS.n9556 VSS.n9555 0.0103214
R22585 VSS.n9525 VSS.n9518 0.0103214
R22586 VSS.n9617 VSS.n9616 0.0103214
R22587 VSS.n9624 VSS.n9623 0.0103214
R22588 VSS.n9637 VSS.n9480 0.0103214
R22589 VSS.n9636 VSS.n9481 0.0103214
R22590 VSS.n9667 VSS.n9455 0.0103214
R22591 VSS.n9458 VSS.n9457 0.0103214
R22592 VSS.n9687 VSS.n9442 0.0103214
R22593 VSS.n9708 VSS.n9421 0.0103214
R22594 VSS.n9741 VSS.n9740 0.0103214
R22595 VSS.n9655 VSS.n9456 0.0103214
R22596 VSS.n9686 VSS.n9685 0.0103214
R22597 VSS.n9681 VSS.n9431 0.0103214
R22598 VSS.n9709 VSS.n9423 0.0103214
R22599 VSS.n9717 VSS.n9716 0.0103214
R22600 VSS.n9791 VSS.n9387 0.0103214
R22601 VSS.n9795 VSS.n9385 0.0103214
R22602 VSS.n9797 VSS.n9383 0.0103214
R22603 VSS.n9790 VSS.n9389 0.0103214
R22604 VSS.n9799 VSS.n9798 0.0103214
R22605 VSS.n9524 VSS.n9519 0.0103214
R22606 VSS.n9598 VSS.n9515 0.0103214
R22607 VSS.n9618 VSS.n9495 0.0103214
R22608 VSS.n9635 VSS.n9634 0.0103214
R22609 VSS.n16492 VSS.n16491 0.0103214
R22610 VSS.n16525 VSS.n16461 0.0103214
R22611 VSS.n16546 VSS.n16438 0.0103214
R22612 VSS.n16570 VSS.n16428 0.0103214
R22613 VSS.n16569 VSS.n16568 0.0103214
R22614 VSS.n16431 VSS.n16429 0.0103214
R22615 VSS.n16610 VSS.n16397 0.0103214
R22616 VSS.n16400 VSS.n16399 0.0103214
R22617 VSS.n16630 VSS.n16384 0.0103214
R22618 VSS.n16651 VSS.n16363 0.0103214
R22619 VSS.n16684 VSS.n16683 0.0103214
R22620 VSS.n16598 VSS.n16398 0.0103214
R22621 VSS.n16629 VSS.n16628 0.0103214
R22622 VSS.n16624 VSS.n16373 0.0103214
R22623 VSS.n16652 VSS.n16365 0.0103214
R22624 VSS.n16660 VSS.n16659 0.0103214
R22625 VSS.n16734 VSS.n16329 0.0103214
R22626 VSS.n16738 VSS.n16327 0.0103214
R22627 VSS.n16740 VSS.n16325 0.0103214
R22628 VSS.n16733 VSS.n16331 0.0103214
R22629 VSS.n16742 VSS.n16741 0.0103214
R22630 VSS.n16524 VSS.n16523 0.0103214
R22631 VSS.n16543 VSS.n16542 0.0103214
R22632 VSS.n16547 VSS.n16440 0.0103214
R22633 VSS.n16430 VSS.n16424 0.0103214
R22634 VSS.n1657 VSS.n1656 0.0103214
R22635 VSS.n1690 VSS.n1626 0.0103214
R22636 VSS.n1711 VSS.n1603 0.0103214
R22637 VSS.n1735 VSS.n1593 0.0103214
R22638 VSS.n1734 VSS.n1733 0.0103214
R22639 VSS.n1596 VSS.n1594 0.0103214
R22640 VSS.n16017 VSS.n1569 0.0103214
R22641 VSS.n1572 VSS.n1571 0.0103214
R22642 VSS.n16037 VSS.n1556 0.0103214
R22643 VSS.n16058 VSS.n1535 0.0103214
R22644 VSS.n16091 VSS.n16090 0.0103214
R22645 VSS.n16005 VSS.n1570 0.0103214
R22646 VSS.n16036 VSS.n16035 0.0103214
R22647 VSS.n16031 VSS.n1545 0.0103214
R22648 VSS.n16059 VSS.n1537 0.0103214
R22649 VSS.n16067 VSS.n16066 0.0103214
R22650 VSS.n16141 VSS.n1501 0.0103214
R22651 VSS.n16145 VSS.n1499 0.0103214
R22652 VSS.n16147 VSS.n1497 0.0103214
R22653 VSS.n16140 VSS.n1503 0.0103214
R22654 VSS.n16149 VSS.n16148 0.0103214
R22655 VSS.n1689 VSS.n1688 0.0103214
R22656 VSS.n1708 VSS.n1707 0.0103214
R22657 VSS.n1712 VSS.n1605 0.0103214
R22658 VSS.n1595 VSS.n1589 0.0103214
R22659 VSS.n1848 VSS.n1847 0.0103214
R22660 VSS.n1817 VSS.n1810 0.0103214
R22661 VSS.n1909 VSS.n1908 0.0103214
R22662 VSS.n1916 VSS.n1915 0.0103214
R22663 VSS.n1929 VSS.n1772 0.0103214
R22664 VSS.n1928 VSS.n1773 0.0103214
R22665 VSS.n2015 VSS.n2005 0.0103214
R22666 VSS.n2339 VSS.n2338 0.0103214
R22667 VSS.n2332 VSS.n1953 0.0103214
R22668 VSS.n2042 VSS.n1962 0.0103214
R22669 VSS.n2064 VSS.n2063 0.0103214
R22670 VSS.n2014 VSS.n2013 0.0103214
R22671 VSS.n2333 VSS.n1951 0.0103214
R22672 VSS.n2329 VSS.n1956 0.0103214
R22673 VSS.n2320 VSS.n1965 0.0103214
R22674 VSS.n2046 VSS.n1968 0.0103214
R22675 VSS.n2291 VSS.n2080 0.0103214
R22676 VSS.n2286 VSS.n2102 0.0103214
R22677 VSS.n2114 VSS.n2108 0.0103214
R22678 VSS.n2290 VSS.n2289 0.0103214
R22679 VSS.n2113 VSS.n2110 0.0103214
R22680 VSS.n1816 VSS.n1811 0.0103214
R22681 VSS.n1890 VSS.n1807 0.0103214
R22682 VSS.n1910 VSS.n1787 0.0103214
R22683 VSS.n1927 VSS.n1926 0.0103214
R22684 VSS.n3047 VSS.n3046 0.0103214
R22685 VSS.n3016 VSS.n3009 0.0103214
R22686 VSS.n3108 VSS.n3107 0.0103214
R22687 VSS.n3115 VSS.n3114 0.0103214
R22688 VSS.n3128 VSS.n2971 0.0103214
R22689 VSS.n3127 VSS.n2972 0.0103214
R22690 VSS.n3158 VSS.n2946 0.0103214
R22691 VSS.n2949 VSS.n2948 0.0103214
R22692 VSS.n3178 VSS.n2933 0.0103214
R22693 VSS.n3199 VSS.n2912 0.0103214
R22694 VSS.n3232 VSS.n3231 0.0103214
R22695 VSS.n3146 VSS.n2947 0.0103214
R22696 VSS.n3177 VSS.n3176 0.0103214
R22697 VSS.n3172 VSS.n2922 0.0103214
R22698 VSS.n3200 VSS.n2914 0.0103214
R22699 VSS.n3208 VSS.n3207 0.0103214
R22700 VSS.n3282 VSS.n2878 0.0103214
R22701 VSS.n3286 VSS.n2876 0.0103214
R22702 VSS.n3288 VSS.n2874 0.0103214
R22703 VSS.n3281 VSS.n2880 0.0103214
R22704 VSS.n3290 VSS.n3289 0.0103214
R22705 VSS.n3015 VSS.n3010 0.0103214
R22706 VSS.n3089 VSS.n3006 0.0103214
R22707 VSS.n3109 VSS.n2986 0.0103214
R22708 VSS.n3126 VSS.n3125 0.0103214
R22709 VSS.n3639 VSS.n3638 0.0103214
R22710 VSS.n3608 VSS.n3601 0.0103214
R22711 VSS.n3700 VSS.n3699 0.0103214
R22712 VSS.n3707 VSS.n3706 0.0103214
R22713 VSS.n3720 VSS.n3563 0.0103214
R22714 VSS.n3719 VSS.n3564 0.0103214
R22715 VSS.n3750 VSS.n3538 0.0103214
R22716 VSS.n3541 VSS.n3540 0.0103214
R22717 VSS.n3770 VSS.n3525 0.0103214
R22718 VSS.n3791 VSS.n3504 0.0103214
R22719 VSS.n3824 VSS.n3823 0.0103214
R22720 VSS.n3738 VSS.n3539 0.0103214
R22721 VSS.n3769 VSS.n3768 0.0103214
R22722 VSS.n3764 VSS.n3514 0.0103214
R22723 VSS.n3792 VSS.n3506 0.0103214
R22724 VSS.n3800 VSS.n3799 0.0103214
R22725 VSS.n3874 VSS.n3470 0.0103214
R22726 VSS.n3878 VSS.n3468 0.0103214
R22727 VSS.n3880 VSS.n3466 0.0103214
R22728 VSS.n3873 VSS.n3472 0.0103214
R22729 VSS.n3882 VSS.n3881 0.0103214
R22730 VSS.n3607 VSS.n3602 0.0103214
R22731 VSS.n3681 VSS.n3598 0.0103214
R22732 VSS.n3701 VSS.n3578 0.0103214
R22733 VSS.n3718 VSS.n3717 0.0103214
R22734 VSS.n4231 VSS.n4230 0.0103214
R22735 VSS.n4200 VSS.n4193 0.0103214
R22736 VSS.n4292 VSS.n4291 0.0103214
R22737 VSS.n4299 VSS.n4298 0.0103214
R22738 VSS.n4312 VSS.n4155 0.0103214
R22739 VSS.n4311 VSS.n4156 0.0103214
R22740 VSS.n4342 VSS.n4130 0.0103214
R22741 VSS.n4133 VSS.n4132 0.0103214
R22742 VSS.n4362 VSS.n4117 0.0103214
R22743 VSS.n4383 VSS.n4096 0.0103214
R22744 VSS.n4416 VSS.n4415 0.0103214
R22745 VSS.n4330 VSS.n4131 0.0103214
R22746 VSS.n4361 VSS.n4360 0.0103214
R22747 VSS.n4356 VSS.n4106 0.0103214
R22748 VSS.n4384 VSS.n4098 0.0103214
R22749 VSS.n4392 VSS.n4391 0.0103214
R22750 VSS.n4466 VSS.n4062 0.0103214
R22751 VSS.n4470 VSS.n4060 0.0103214
R22752 VSS.n4472 VSS.n4058 0.0103214
R22753 VSS.n4465 VSS.n4064 0.0103214
R22754 VSS.n4474 VSS.n4473 0.0103214
R22755 VSS.n4199 VSS.n4194 0.0103214
R22756 VSS.n4273 VSS.n4190 0.0103214
R22757 VSS.n4293 VSS.n4170 0.0103214
R22758 VSS.n4310 VSS.n4309 0.0103214
R22759 VSS.n4823 VSS.n4822 0.0103214
R22760 VSS.n4792 VSS.n4785 0.0103214
R22761 VSS.n4884 VSS.n4883 0.0103214
R22762 VSS.n4891 VSS.n4890 0.0103214
R22763 VSS.n4904 VSS.n4747 0.0103214
R22764 VSS.n4903 VSS.n4748 0.0103214
R22765 VSS.n4934 VSS.n4722 0.0103214
R22766 VSS.n4725 VSS.n4724 0.0103214
R22767 VSS.n4954 VSS.n4709 0.0103214
R22768 VSS.n4975 VSS.n4688 0.0103214
R22769 VSS.n5008 VSS.n5007 0.0103214
R22770 VSS.n4922 VSS.n4723 0.0103214
R22771 VSS.n4953 VSS.n4952 0.0103214
R22772 VSS.n4948 VSS.n4698 0.0103214
R22773 VSS.n4976 VSS.n4690 0.0103214
R22774 VSS.n4984 VSS.n4983 0.0103214
R22775 VSS.n5058 VSS.n4654 0.0103214
R22776 VSS.n5062 VSS.n4652 0.0103214
R22777 VSS.n5064 VSS.n4650 0.0103214
R22778 VSS.n5057 VSS.n4656 0.0103214
R22779 VSS.n5066 VSS.n5065 0.0103214
R22780 VSS.n4791 VSS.n4786 0.0103214
R22781 VSS.n4865 VSS.n4782 0.0103214
R22782 VSS.n4885 VSS.n4762 0.0103214
R22783 VSS.n4902 VSS.n4901 0.0103214
R22784 VSS.n2444 VSS.n2443 0.0103214
R22785 VSS.n2413 VSS.n2406 0.0103214
R22786 VSS.n2505 VSS.n2504 0.0103214
R22787 VSS.n2512 VSS.n2511 0.0103214
R22788 VSS.n2525 VSS.n2368 0.0103214
R22789 VSS.n2524 VSS.n2369 0.0103214
R22790 VSS.n2611 VSS.n2601 0.0103214
R22791 VSS.n5304 VSS.n5303 0.0103214
R22792 VSS.n5297 VSS.n2549 0.0103214
R22793 VSS.n2638 VSS.n2558 0.0103214
R22794 VSS.n2660 VSS.n2659 0.0103214
R22795 VSS.n2610 VSS.n2609 0.0103214
R22796 VSS.n5298 VSS.n2547 0.0103214
R22797 VSS.n5294 VSS.n2552 0.0103214
R22798 VSS.n5285 VSS.n2561 0.0103214
R22799 VSS.n2642 VSS.n2564 0.0103214
R22800 VSS.n5256 VSS.n2676 0.0103214
R22801 VSS.n5251 VSS.n2698 0.0103214
R22802 VSS.n2710 VSS.n2704 0.0103214
R22803 VSS.n5255 VSS.n5254 0.0103214
R22804 VSS.n2709 VSS.n2706 0.0103214
R22805 VSS.n2412 VSS.n2407 0.0103214
R22806 VSS.n2486 VSS.n2403 0.0103214
R22807 VSS.n2506 VSS.n2383 0.0103214
R22808 VSS.n2523 VSS.n2522 0.0103214
R22809 VSS.n5405 VSS.n5404 0.0103214
R22810 VSS.n5374 VSS.n5367 0.0103214
R22811 VSS.n5466 VSS.n5465 0.0103214
R22812 VSS.n5473 VSS.n5472 0.0103214
R22813 VSS.n5486 VSS.n5329 0.0103214
R22814 VSS.n5485 VSS.n5330 0.0103214
R22815 VSS.n5572 VSS.n5562 0.0103214
R22816 VSS.n5877 VSS.n5876 0.0103214
R22817 VSS.n5870 VSS.n5510 0.0103214
R22818 VSS.n5599 VSS.n5519 0.0103214
R22819 VSS.n5621 VSS.n5620 0.0103214
R22820 VSS.n5571 VSS.n5570 0.0103214
R22821 VSS.n5871 VSS.n5508 0.0103214
R22822 VSS.n5867 VSS.n5513 0.0103214
R22823 VSS.n5858 VSS.n5522 0.0103214
R22824 VSS.n5603 VSS.n5525 0.0103214
R22825 VSS.n5829 VSS.n5637 0.0103214
R22826 VSS.n5824 VSS.n5659 0.0103214
R22827 VSS.n5671 VSS.n5665 0.0103214
R22828 VSS.n5828 VSS.n5827 0.0103214
R22829 VSS.n5670 VSS.n5667 0.0103214
R22830 VSS.n5373 VSS.n5368 0.0103214
R22831 VSS.n5447 VSS.n5364 0.0103214
R22832 VSS.n5467 VSS.n5344 0.0103214
R22833 VSS.n5484 VSS.n5483 0.0103214
R22834 VSS.n5978 VSS.n5977 0.0103214
R22835 VSS.n5947 VSS.n5940 0.0103214
R22836 VSS.n6039 VSS.n6038 0.0103214
R22837 VSS.n6046 VSS.n6045 0.0103214
R22838 VSS.n6059 VSS.n5902 0.0103214
R22839 VSS.n6058 VSS.n5903 0.0103214
R22840 VSS.n6145 VSS.n6135 0.0103214
R22841 VSS.n6469 VSS.n6468 0.0103214
R22842 VSS.n6462 VSS.n6083 0.0103214
R22843 VSS.n6172 VSS.n6092 0.0103214
R22844 VSS.n6194 VSS.n6193 0.0103214
R22845 VSS.n6144 VSS.n6143 0.0103214
R22846 VSS.n6463 VSS.n6081 0.0103214
R22847 VSS.n6459 VSS.n6086 0.0103214
R22848 VSS.n6450 VSS.n6095 0.0103214
R22849 VSS.n6176 VSS.n6098 0.0103214
R22850 VSS.n6421 VSS.n6210 0.0103214
R22851 VSS.n6416 VSS.n6232 0.0103214
R22852 VSS.n6244 VSS.n6238 0.0103214
R22853 VSS.n6420 VSS.n6419 0.0103214
R22854 VSS.n6243 VSS.n6240 0.0103214
R22855 VSS.n5946 VSS.n5941 0.0103214
R22856 VSS.n6020 VSS.n5937 0.0103214
R22857 VSS.n6040 VSS.n5917 0.0103214
R22858 VSS.n6057 VSS.n6056 0.0103214
R22859 VSS.n7780 VSS.n7779 0.0103214
R22860 VSS.n7749 VSS.n7742 0.0103214
R22861 VSS.n7841 VSS.n7840 0.0103214
R22862 VSS.n7848 VSS.n7847 0.0103214
R22863 VSS.n7861 VSS.n7704 0.0103214
R22864 VSS.n7860 VSS.n7705 0.0103214
R22865 VSS.n7891 VSS.n7679 0.0103214
R22866 VSS.n7682 VSS.n7681 0.0103214
R22867 VSS.n7911 VSS.n7666 0.0103214
R22868 VSS.n7932 VSS.n7645 0.0103214
R22869 VSS.n7965 VSS.n7964 0.0103214
R22870 VSS.n7879 VSS.n7680 0.0103214
R22871 VSS.n7910 VSS.n7909 0.0103214
R22872 VSS.n7905 VSS.n7655 0.0103214
R22873 VSS.n7933 VSS.n7647 0.0103214
R22874 VSS.n7941 VSS.n7940 0.0103214
R22875 VSS.n8015 VSS.n7611 0.0103214
R22876 VSS.n8019 VSS.n7609 0.0103214
R22877 VSS.n8021 VSS.n7607 0.0103214
R22878 VSS.n8014 VSS.n7613 0.0103214
R22879 VSS.n8023 VSS.n8022 0.0103214
R22880 VSS.n7748 VSS.n7743 0.0103214
R22881 VSS.n7822 VSS.n7739 0.0103214
R22882 VSS.n7842 VSS.n7719 0.0103214
R22883 VSS.n7859 VSS.n7858 0.0103214
R22884 VSS.n8372 VSS.n8371 0.0103214
R22885 VSS.n8341 VSS.n8334 0.0103214
R22886 VSS.n8433 VSS.n8432 0.0103214
R22887 VSS.n8440 VSS.n8439 0.0103214
R22888 VSS.n8453 VSS.n8296 0.0103214
R22889 VSS.n8452 VSS.n8297 0.0103214
R22890 VSS.n8483 VSS.n8271 0.0103214
R22891 VSS.n8274 VSS.n8273 0.0103214
R22892 VSS.n8503 VSS.n8258 0.0103214
R22893 VSS.n8524 VSS.n8237 0.0103214
R22894 VSS.n8557 VSS.n8556 0.0103214
R22895 VSS.n8471 VSS.n8272 0.0103214
R22896 VSS.n8502 VSS.n8501 0.0103214
R22897 VSS.n8497 VSS.n8247 0.0103214
R22898 VSS.n8525 VSS.n8239 0.0103214
R22899 VSS.n8533 VSS.n8532 0.0103214
R22900 VSS.n8607 VSS.n8203 0.0103214
R22901 VSS.n8611 VSS.n8201 0.0103214
R22902 VSS.n8613 VSS.n8199 0.0103214
R22903 VSS.n8606 VSS.n8205 0.0103214
R22904 VSS.n8615 VSS.n8614 0.0103214
R22905 VSS.n8340 VSS.n8335 0.0103214
R22906 VSS.n8414 VSS.n8331 0.0103214
R22907 VSS.n8434 VSS.n8311 0.0103214
R22908 VSS.n8451 VSS.n8450 0.0103214
R22909 VSS.n8964 VSS.n8963 0.0103214
R22910 VSS.n8933 VSS.n8926 0.0103214
R22911 VSS.n9025 VSS.n9024 0.0103214
R22912 VSS.n9032 VSS.n9031 0.0103214
R22913 VSS.n9045 VSS.n8888 0.0103214
R22914 VSS.n9044 VSS.n8889 0.0103214
R22915 VSS.n9075 VSS.n8863 0.0103214
R22916 VSS.n8866 VSS.n8865 0.0103214
R22917 VSS.n9095 VSS.n8850 0.0103214
R22918 VSS.n9116 VSS.n8829 0.0103214
R22919 VSS.n9149 VSS.n9148 0.0103214
R22920 VSS.n9063 VSS.n8864 0.0103214
R22921 VSS.n9094 VSS.n9093 0.0103214
R22922 VSS.n9089 VSS.n8839 0.0103214
R22923 VSS.n9117 VSS.n8831 0.0103214
R22924 VSS.n9125 VSS.n9124 0.0103214
R22925 VSS.n9199 VSS.n8795 0.0103214
R22926 VSS.n9203 VSS.n8793 0.0103214
R22927 VSS.n9205 VSS.n8791 0.0103214
R22928 VSS.n9198 VSS.n8797 0.0103214
R22929 VSS.n9207 VSS.n9206 0.0103214
R22930 VSS.n8932 VSS.n8927 0.0103214
R22931 VSS.n9006 VSS.n8923 0.0103214
R22932 VSS.n9026 VSS.n8903 0.0103214
R22933 VSS.n9043 VSS.n9042 0.0103214
R22934 VSS.n10148 VSS.n10147 0.0103214
R22935 VSS.n10117 VSS.n10110 0.0103214
R22936 VSS.n10209 VSS.n10208 0.0103214
R22937 VSS.n10216 VSS.n10215 0.0103214
R22938 VSS.n10229 VSS.n10072 0.0103214
R22939 VSS.n10228 VSS.n10073 0.0103214
R22940 VSS.n10259 VSS.n10047 0.0103214
R22941 VSS.n10050 VSS.n10049 0.0103214
R22942 VSS.n10279 VSS.n10034 0.0103214
R22943 VSS.n10300 VSS.n10013 0.0103214
R22944 VSS.n10333 VSS.n10332 0.0103214
R22945 VSS.n10247 VSS.n10048 0.0103214
R22946 VSS.n10278 VSS.n10277 0.0103214
R22947 VSS.n10273 VSS.n10023 0.0103214
R22948 VSS.n10301 VSS.n10015 0.0103214
R22949 VSS.n10309 VSS.n10308 0.0103214
R22950 VSS.n10383 VSS.n9979 0.0103214
R22951 VSS.n10387 VSS.n9977 0.0103214
R22952 VSS.n10389 VSS.n9975 0.0103214
R22953 VSS.n10382 VSS.n9981 0.0103214
R22954 VSS.n10391 VSS.n10390 0.0103214
R22955 VSS.n10116 VSS.n10111 0.0103214
R22956 VSS.n10190 VSS.n10107 0.0103214
R22957 VSS.n10210 VSS.n10087 0.0103214
R22958 VSS.n10227 VSS.n10226 0.0103214
R22959 VSS.n10740 VSS.n10739 0.0103214
R22960 VSS.n10709 VSS.n10702 0.0103214
R22961 VSS.n10801 VSS.n10800 0.0103214
R22962 VSS.n10808 VSS.n10807 0.0103214
R22963 VSS.n10821 VSS.n10664 0.0103214
R22964 VSS.n10820 VSS.n10665 0.0103214
R22965 VSS.n10851 VSS.n10639 0.0103214
R22966 VSS.n10642 VSS.n10641 0.0103214
R22967 VSS.n10871 VSS.n10626 0.0103214
R22968 VSS.n10892 VSS.n10605 0.0103214
R22969 VSS.n10925 VSS.n10924 0.0103214
R22970 VSS.n10839 VSS.n10640 0.0103214
R22971 VSS.n10870 VSS.n10869 0.0103214
R22972 VSS.n10865 VSS.n10615 0.0103214
R22973 VSS.n10893 VSS.n10607 0.0103214
R22974 VSS.n10901 VSS.n10900 0.0103214
R22975 VSS.n10975 VSS.n10571 0.0103214
R22976 VSS.n10979 VSS.n10569 0.0103214
R22977 VSS.n10981 VSS.n10567 0.0103214
R22978 VSS.n10974 VSS.n10573 0.0103214
R22979 VSS.n10983 VSS.n10982 0.0103214
R22980 VSS.n10708 VSS.n10703 0.0103214
R22981 VSS.n10782 VSS.n10699 0.0103214
R22982 VSS.n10802 VSS.n10679 0.0103214
R22983 VSS.n10819 VSS.n10818 0.0103214
R22984 VSS.n11332 VSS.n11331 0.0103214
R22985 VSS.n11301 VSS.n11294 0.0103214
R22986 VSS.n11393 VSS.n11392 0.0103214
R22987 VSS.n11400 VSS.n11399 0.0103214
R22988 VSS.n11413 VSS.n11256 0.0103214
R22989 VSS.n11412 VSS.n11257 0.0103214
R22990 VSS.n11443 VSS.n11231 0.0103214
R22991 VSS.n11234 VSS.n11233 0.0103214
R22992 VSS.n11463 VSS.n11218 0.0103214
R22993 VSS.n11484 VSS.n11197 0.0103214
R22994 VSS.n11517 VSS.n11516 0.0103214
R22995 VSS.n11431 VSS.n11232 0.0103214
R22996 VSS.n11462 VSS.n11461 0.0103214
R22997 VSS.n11457 VSS.n11207 0.0103214
R22998 VSS.n11485 VSS.n11199 0.0103214
R22999 VSS.n11493 VSS.n11492 0.0103214
R23000 VSS.n11567 VSS.n11163 0.0103214
R23001 VSS.n11571 VSS.n11161 0.0103214
R23002 VSS.n11573 VSS.n11159 0.0103214
R23003 VSS.n11566 VSS.n11165 0.0103214
R23004 VSS.n11575 VSS.n11574 0.0103214
R23005 VSS.n11300 VSS.n11295 0.0103214
R23006 VSS.n11374 VSS.n11291 0.0103214
R23007 VSS.n11394 VSS.n11271 0.0103214
R23008 VSS.n11411 VSS.n11410 0.0103214
R23009 VSS.n11924 VSS.n11923 0.0103214
R23010 VSS.n11893 VSS.n11886 0.0103214
R23011 VSS.n11985 VSS.n11984 0.0103214
R23012 VSS.n11992 VSS.n11991 0.0103214
R23013 VSS.n12005 VSS.n11848 0.0103214
R23014 VSS.n12004 VSS.n11849 0.0103214
R23015 VSS.n12035 VSS.n11823 0.0103214
R23016 VSS.n11826 VSS.n11825 0.0103214
R23017 VSS.n12055 VSS.n11810 0.0103214
R23018 VSS.n12076 VSS.n11789 0.0103214
R23019 VSS.n12109 VSS.n12108 0.0103214
R23020 VSS.n12023 VSS.n11824 0.0103214
R23021 VSS.n12054 VSS.n12053 0.0103214
R23022 VSS.n12049 VSS.n11799 0.0103214
R23023 VSS.n12077 VSS.n11791 0.0103214
R23024 VSS.n12085 VSS.n12084 0.0103214
R23025 VSS.n12159 VSS.n11755 0.0103214
R23026 VSS.n12163 VSS.n11753 0.0103214
R23027 VSS.n12165 VSS.n11751 0.0103214
R23028 VSS.n12158 VSS.n11757 0.0103214
R23029 VSS.n12167 VSS.n12166 0.0103214
R23030 VSS.n11892 VSS.n11887 0.0103214
R23031 VSS.n11966 VSS.n11883 0.0103214
R23032 VSS.n11986 VSS.n11863 0.0103214
R23033 VSS.n12003 VSS.n12002 0.0103214
R23034 VSS.n12516 VSS.n12515 0.0103214
R23035 VSS.n12485 VSS.n12478 0.0103214
R23036 VSS.n12577 VSS.n12576 0.0103214
R23037 VSS.n12584 VSS.n12583 0.0103214
R23038 VSS.n12597 VSS.n12440 0.0103214
R23039 VSS.n12596 VSS.n12441 0.0103214
R23040 VSS.n12627 VSS.n12415 0.0103214
R23041 VSS.n12418 VSS.n12417 0.0103214
R23042 VSS.n12647 VSS.n12402 0.0103214
R23043 VSS.n12668 VSS.n12381 0.0103214
R23044 VSS.n12701 VSS.n12700 0.0103214
R23045 VSS.n12615 VSS.n12416 0.0103214
R23046 VSS.n12646 VSS.n12645 0.0103214
R23047 VSS.n12641 VSS.n12391 0.0103214
R23048 VSS.n12669 VSS.n12383 0.0103214
R23049 VSS.n12677 VSS.n12676 0.0103214
R23050 VSS.n12751 VSS.n12347 0.0103214
R23051 VSS.n12755 VSS.n12345 0.0103214
R23052 VSS.n12757 VSS.n12343 0.0103214
R23053 VSS.n12750 VSS.n12349 0.0103214
R23054 VSS.n12759 VSS.n12758 0.0103214
R23055 VSS.n12484 VSS.n12479 0.0103214
R23056 VSS.n12558 VSS.n12475 0.0103214
R23057 VSS.n12578 VSS.n12455 0.0103214
R23058 VSS.n12595 VSS.n12594 0.0103214
R23059 VSS.n13108 VSS.n13107 0.0103214
R23060 VSS.n13077 VSS.n13070 0.0103214
R23061 VSS.n13169 VSS.n13168 0.0103214
R23062 VSS.n13176 VSS.n13175 0.0103214
R23063 VSS.n13189 VSS.n13032 0.0103214
R23064 VSS.n13188 VSS.n13033 0.0103214
R23065 VSS.n13219 VSS.n13007 0.0103214
R23066 VSS.n13010 VSS.n13009 0.0103214
R23067 VSS.n13239 VSS.n12994 0.0103214
R23068 VSS.n13260 VSS.n12973 0.0103214
R23069 VSS.n13293 VSS.n13292 0.0103214
R23070 VSS.n13207 VSS.n13008 0.0103214
R23071 VSS.n13238 VSS.n13237 0.0103214
R23072 VSS.n13233 VSS.n12983 0.0103214
R23073 VSS.n13261 VSS.n12975 0.0103214
R23074 VSS.n13269 VSS.n13268 0.0103214
R23075 VSS.n13343 VSS.n12939 0.0103214
R23076 VSS.n13347 VSS.n12937 0.0103214
R23077 VSS.n13349 VSS.n12935 0.0103214
R23078 VSS.n13342 VSS.n12941 0.0103214
R23079 VSS.n13351 VSS.n13350 0.0103214
R23080 VSS.n13076 VSS.n13071 0.0103214
R23081 VSS.n13150 VSS.n13067 0.0103214
R23082 VSS.n13170 VSS.n13047 0.0103214
R23083 VSS.n13187 VSS.n13186 0.0103214
R23084 VSS.n13700 VSS.n13699 0.0103214
R23085 VSS.n13669 VSS.n13662 0.0103214
R23086 VSS.n13761 VSS.n13760 0.0103214
R23087 VSS.n13768 VSS.n13767 0.0103214
R23088 VSS.n13781 VSS.n13624 0.0103214
R23089 VSS.n13780 VSS.n13625 0.0103214
R23090 VSS.n13811 VSS.n13599 0.0103214
R23091 VSS.n13602 VSS.n13601 0.0103214
R23092 VSS.n13831 VSS.n13586 0.0103214
R23093 VSS.n13852 VSS.n13565 0.0103214
R23094 VSS.n13885 VSS.n13884 0.0103214
R23095 VSS.n13799 VSS.n13600 0.0103214
R23096 VSS.n13830 VSS.n13829 0.0103214
R23097 VSS.n13825 VSS.n13575 0.0103214
R23098 VSS.n13853 VSS.n13567 0.0103214
R23099 VSS.n13861 VSS.n13860 0.0103214
R23100 VSS.n13935 VSS.n13531 0.0103214
R23101 VSS.n13939 VSS.n13529 0.0103214
R23102 VSS.n13941 VSS.n13527 0.0103214
R23103 VSS.n13934 VSS.n13533 0.0103214
R23104 VSS.n13943 VSS.n13942 0.0103214
R23105 VSS.n13668 VSS.n13663 0.0103214
R23106 VSS.n13742 VSS.n13659 0.0103214
R23107 VSS.n13762 VSS.n13639 0.0103214
R23108 VSS.n13779 VSS.n13778 0.0103214
R23109 VSS.n14292 VSS.n14291 0.0103214
R23110 VSS.n14261 VSS.n14254 0.0103214
R23111 VSS.n14353 VSS.n14352 0.0103214
R23112 VSS.n14360 VSS.n14359 0.0103214
R23113 VSS.n14373 VSS.n14216 0.0103214
R23114 VSS.n14372 VSS.n14217 0.0103214
R23115 VSS.n14403 VSS.n14191 0.0103214
R23116 VSS.n14194 VSS.n14193 0.0103214
R23117 VSS.n14423 VSS.n14178 0.0103214
R23118 VSS.n14444 VSS.n14157 0.0103214
R23119 VSS.n14477 VSS.n14476 0.0103214
R23120 VSS.n14391 VSS.n14192 0.0103214
R23121 VSS.n14422 VSS.n14421 0.0103214
R23122 VSS.n14417 VSS.n14167 0.0103214
R23123 VSS.n14445 VSS.n14159 0.0103214
R23124 VSS.n14453 VSS.n14452 0.0103214
R23125 VSS.n14527 VSS.n14123 0.0103214
R23126 VSS.n14531 VSS.n14121 0.0103214
R23127 VSS.n14533 VSS.n14119 0.0103214
R23128 VSS.n14526 VSS.n14125 0.0103214
R23129 VSS.n14535 VSS.n14534 0.0103214
R23130 VSS.n14260 VSS.n14255 0.0103214
R23131 VSS.n14334 VSS.n14251 0.0103214
R23132 VSS.n14354 VSS.n14231 0.0103214
R23133 VSS.n14371 VSS.n14370 0.0103214
R23134 VSS.n14884 VSS.n14883 0.0103214
R23135 VSS.n14853 VSS.n14846 0.0103214
R23136 VSS.n14945 VSS.n14944 0.0103214
R23137 VSS.n14952 VSS.n14951 0.0103214
R23138 VSS.n14965 VSS.n14808 0.0103214
R23139 VSS.n14964 VSS.n14809 0.0103214
R23140 VSS.n14995 VSS.n14783 0.0103214
R23141 VSS.n14786 VSS.n14785 0.0103214
R23142 VSS.n15015 VSS.n14770 0.0103214
R23143 VSS.n15036 VSS.n14749 0.0103214
R23144 VSS.n15069 VSS.n15068 0.0103214
R23145 VSS.n14983 VSS.n14784 0.0103214
R23146 VSS.n15014 VSS.n15013 0.0103214
R23147 VSS.n15009 VSS.n14759 0.0103214
R23148 VSS.n15037 VSS.n14751 0.0103214
R23149 VSS.n15045 VSS.n15044 0.0103214
R23150 VSS.n15119 VSS.n14715 0.0103214
R23151 VSS.n15123 VSS.n14713 0.0103214
R23152 VSS.n15125 VSS.n14711 0.0103214
R23153 VSS.n15118 VSS.n14717 0.0103214
R23154 VSS.n15127 VSS.n15126 0.0103214
R23155 VSS.n14852 VSS.n14847 0.0103214
R23156 VSS.n14926 VSS.n14843 0.0103214
R23157 VSS.n14946 VSS.n14823 0.0103214
R23158 VSS.n14963 VSS.n14962 0.0103214
R23159 VSS.n15476 VSS.n15475 0.0103214
R23160 VSS.n15445 VSS.n15438 0.0103214
R23161 VSS.n15537 VSS.n15536 0.0103214
R23162 VSS.n15544 VSS.n15543 0.0103214
R23163 VSS.n15557 VSS.n15400 0.0103214
R23164 VSS.n15556 VSS.n15401 0.0103214
R23165 VSS.n15587 VSS.n15375 0.0103214
R23166 VSS.n15378 VSS.n15377 0.0103214
R23167 VSS.n15607 VSS.n15362 0.0103214
R23168 VSS.n15628 VSS.n15341 0.0103214
R23169 VSS.n15661 VSS.n15660 0.0103214
R23170 VSS.n15575 VSS.n15376 0.0103214
R23171 VSS.n15606 VSS.n15605 0.0103214
R23172 VSS.n15601 VSS.n15351 0.0103214
R23173 VSS.n15629 VSS.n15343 0.0103214
R23174 VSS.n15637 VSS.n15636 0.0103214
R23175 VSS.n15711 VSS.n15307 0.0103214
R23176 VSS.n15715 VSS.n15305 0.0103214
R23177 VSS.n15717 VSS.n15303 0.0103214
R23178 VSS.n15710 VSS.n15309 0.0103214
R23179 VSS.n15719 VSS.n15718 0.0103214
R23180 VSS.n15444 VSS.n15439 0.0103214
R23181 VSS.n15518 VSS.n15435 0.0103214
R23182 VSS.n15538 VSS.n15415 0.0103214
R23183 VSS.n15555 VSS.n15554 0.0103214
R23184 VSS.n6584 VSS.n6583 0.0103214
R23185 VSS.n6553 VSS.n6546 0.0103214
R23186 VSS.n6645 VSS.n6644 0.0103214
R23187 VSS.n6652 VSS.n6651 0.0103214
R23188 VSS.n6665 VSS.n6508 0.0103214
R23189 VSS.n6664 VSS.n6509 0.0103214
R23190 VSS.n6751 VSS.n6741 0.0103214
R23191 VSS.n15957 VSS.n15956 0.0103214
R23192 VSS.n15950 VSS.n6689 0.0103214
R23193 VSS.n6778 VSS.n6698 0.0103214
R23194 VSS.n6800 VSS.n6799 0.0103214
R23195 VSS.n6750 VSS.n6749 0.0103214
R23196 VSS.n15951 VSS.n6687 0.0103214
R23197 VSS.n15947 VSS.n6692 0.0103214
R23198 VSS.n15938 VSS.n6701 0.0103214
R23199 VSS.n6782 VSS.n6704 0.0103214
R23200 VSS.n15909 VSS.n6816 0.0103214
R23201 VSS.n15904 VSS.n6838 0.0103214
R23202 VSS.n6850 VSS.n6844 0.0103214
R23203 VSS.n15908 VSS.n15907 0.0103214
R23204 VSS.n6849 VSS.n6846 0.0103214
R23205 VSS.n6552 VSS.n6547 0.0103214
R23206 VSS.n6626 VSS.n6543 0.0103214
R23207 VSS.n6646 VSS.n6523 0.0103214
R23208 VSS.n6663 VSS.n6662 0.0103214
R23209 VSS.n7181 VSS.n7180 0.0103214
R23210 VSS.n7214 VSS.n7150 0.0103214
R23211 VSS.n7235 VSS.n7127 0.0103214
R23212 VSS.n7259 VSS.n7117 0.0103214
R23213 VSS.n7258 VSS.n7257 0.0103214
R23214 VSS.n7120 VSS.n7118 0.0103214
R23215 VSS.n7299 VSS.n7086 0.0103214
R23216 VSS.n7089 VSS.n7088 0.0103214
R23217 VSS.n7319 VSS.n7073 0.0103214
R23218 VSS.n7340 VSS.n7052 0.0103214
R23219 VSS.n7373 VSS.n7372 0.0103214
R23220 VSS.n7287 VSS.n7087 0.0103214
R23221 VSS.n7318 VSS.n7317 0.0103214
R23222 VSS.n7313 VSS.n7062 0.0103214
R23223 VSS.n7341 VSS.n7054 0.0103214
R23224 VSS.n7349 VSS.n7348 0.0103214
R23225 VSS.n7423 VSS.n7018 0.0103214
R23226 VSS.n7427 VSS.n7016 0.0103214
R23227 VSS.n7429 VSS.n7014 0.0103214
R23228 VSS.n7422 VSS.n7020 0.0103214
R23229 VSS.n7431 VSS.n7430 0.0103214
R23230 VSS.n7213 VSS.n7212 0.0103214
R23231 VSS.n7232 VSS.n7231 0.0103214
R23232 VSS.n7236 VSS.n7129 0.0103214
R23233 VSS.n7119 VSS.n7113 0.0103214
R23234 VSS.n355 VSS.n345 0.0103214
R23235 VSS.n436 VSS.n303 0.0103214
R23236 VSS.n333 VSS.n313 0.0103214
R23237 VSS.n419 VSS.n418 0.0103214
R23238 VSS.n395 VSS.n322 0.0103214
R23239 VSS.n407 VSS.n327 0.0103214
R23240 VSS.n18611 VSS.n184 0.0103214
R23241 VSS.n187 VSS.n186 0.0103214
R23242 VSS.n18631 VSS.n171 0.0103214
R23243 VSS.n18652 VSS.n150 0.0103214
R23244 VSS.n18685 VSS.n18684 0.0103214
R23245 VSS.n18599 VSS.n185 0.0103214
R23246 VSS.n18630 VSS.n18629 0.0103214
R23247 VSS.n18625 VSS.n160 0.0103214
R23248 VSS.n18653 VSS.n152 0.0103214
R23249 VSS.n18661 VSS.n18660 0.0103214
R23250 VSS.n18735 VSS.n116 0.0103214
R23251 VSS.n18739 VSS.n114 0.0103214
R23252 VSS.n18741 VSS.n112 0.0103214
R23253 VSS.n18734 VSS.n118 0.0103214
R23254 VSS.n18743 VSS.n18742 0.0103214
R23255 VSS.n437 VSS.n301 0.0103214
R23256 VSS.n314 VSS.n311 0.0103214
R23257 VSS.n424 VSS.n316 0.0103214
R23258 VSS.n408 VSS.n326 0.0103214
R23259 VSS.n574 VSS.n566 0.0103214
R23260 VSS.n871 VSS.n870 0.0103214
R23261 VSS.n864 VSS.n509 0.0103214
R23262 VSS.n601 VSS.n518 0.0103214
R23263 VSS.n623 VSS.n622 0.0103214
R23264 VSS.n573 VSS.n572 0.0103214
R23265 VSS.n865 VSS.n507 0.0103214
R23266 VSS.n861 VSS.n512 0.0103214
R23267 VSS.n852 VSS.n521 0.0103214
R23268 VSS.n605 VSS.n524 0.0103214
R23269 VSS.n823 VSS.n639 0.0103214
R23270 VSS.n818 VSS.n661 0.0103214
R23271 VSS.n673 VSS.n667 0.0103214
R23272 VSS.n822 VSS.n821 0.0103214
R23273 VSS.n672 VSS.n669 0.0103214
R23274 VSS.n1002 VSS.n467 0.0103214
R23275 VSS.n480 VSS.n477 0.0103214
R23276 VSS.n989 VSS.n482 0.0103214
R23277 VSS.n963 VSS.n889 0.0103214
R23278 VSS.n17937 VSS.n1298 0.0103214
R23279 VSS.n17932 VSS.n1320 0.0103214
R23280 VSS.n1332 VSS.n1326 0.0103214
R23281 VSS.n17936 VSS.n17935 0.0103214
R23282 VSS.n1331 VSS.n1328 0.0103214
R23283 VSS.n17191 VSS.n17190 0.00956429
R23284 VSS.n17208 VSS.n17191 0.00956429
R23285 VSS.n17783 VSS.n17782 0.00956429
R23286 VSS.n17800 VSS.n17783 0.00956429
R23287 VSS.n18503 VSS.n18352 0.00956429
R23288 VSS.n18398 VSS.n18352 0.00956429
R23289 VSS.n9833 VSS.n9832 0.00956429
R23290 VSS.n9850 VSS.n9833 0.00956429
R23291 VSS.n16776 VSS.n16775 0.00956429
R23292 VSS.n16793 VSS.n16776 0.00956429
R23293 VSS.n16183 VSS.n16182 0.00956429
R23294 VSS.n16200 VSS.n16183 0.00956429
R23295 VSS.n2151 VSS.n2150 0.00956429
R23296 VSS.n2256 VSS.n2151 0.00956429
R23297 VSS.n3324 VSS.n3323 0.00956429
R23298 VSS.n3341 VSS.n3324 0.00956429
R23299 VSS.n3916 VSS.n3915 0.00956429
R23300 VSS.n3933 VSS.n3916 0.00956429
R23301 VSS.n4508 VSS.n4507 0.00956429
R23302 VSS.n4525 VSS.n4508 0.00956429
R23303 VSS.n5100 VSS.n5099 0.00956429
R23304 VSS.n5117 VSS.n5100 0.00956429
R23305 VSS.n2747 VSS.n2746 0.00956429
R23306 VSS.n5221 VSS.n2747 0.00956429
R23307 VSS.n5708 VSS.n5707 0.00956429
R23308 VSS.n5794 VSS.n5708 0.00956429
R23309 VSS.n6281 VSS.n6280 0.00956429
R23310 VSS.n6386 VSS.n6281 0.00956429
R23311 VSS.n8057 VSS.n8056 0.00956429
R23312 VSS.n8074 VSS.n8057 0.00956429
R23313 VSS.n8649 VSS.n8648 0.00956429
R23314 VSS.n8666 VSS.n8649 0.00956429
R23315 VSS.n9241 VSS.n9240 0.00956429
R23316 VSS.n9258 VSS.n9241 0.00956429
R23317 VSS.n10425 VSS.n10424 0.00956429
R23318 VSS.n10442 VSS.n10425 0.00956429
R23319 VSS.n11017 VSS.n11016 0.00956429
R23320 VSS.n11034 VSS.n11017 0.00956429
R23321 VSS.n11609 VSS.n11608 0.00956429
R23322 VSS.n11626 VSS.n11609 0.00956429
R23323 VSS.n12201 VSS.n12200 0.00956429
R23324 VSS.n12218 VSS.n12201 0.00956429
R23325 VSS.n12793 VSS.n12792 0.00956429
R23326 VSS.n12810 VSS.n12793 0.00956429
R23327 VSS.n13385 VSS.n13384 0.00956429
R23328 VSS.n13402 VSS.n13385 0.00956429
R23329 VSS.n13977 VSS.n13976 0.00956429
R23330 VSS.n13994 VSS.n13977 0.00956429
R23331 VSS.n14569 VSS.n14568 0.00956429
R23332 VSS.n14586 VSS.n14569 0.00956429
R23333 VSS.n15161 VSS.n15160 0.00956429
R23334 VSS.n15178 VSS.n15161 0.00956429
R23335 VSS.n15753 VSS.n15752 0.00956429
R23336 VSS.n15770 VSS.n15753 0.00956429
R23337 VSS.n6887 VSS.n6886 0.00956429
R23338 VSS.n15874 VSS.n6887 0.00956429
R23339 VSS.n7465 VSS.n7464 0.00956429
R23340 VSS.n7482 VSS.n7465 0.00956429
R23341 VSS.n18777 VSS.n18776 0.00956429
R23342 VSS.n18794 VSS.n18777 0.00956429
R23343 VSS.n710 VSS.n709 0.00956429
R23344 VSS.n788 VSS.n710 0.00956429
R23345 VSS.n1369 VSS.n1368 0.00956429
R23346 VSS.n17902 VSS.n1369 0.00956429
R23347 VSS.n1227 VSS.n1226 0.00942857
R23348 VSS.n17961 VSS.n17960 0.00942857
R23349 VSS.n1277 VSS.n1276 0.00942857
R23350 VSS.n1225 VSS.n1224 0.00942857
R23351 VSS.n1238 VSS.n1167 0.00942857
R23352 VSS.n1181 VSS.n1178 0.00942857
R23353 VSS.n1278 VSS.n1204 0.00942857
R23354 VSS.n919 VSS.n909 0.00942857
R23355 VSS.n1008 VSS.n1007 0.00942857
R23356 VSS.n888 VSS.n493 0.00942857
R23357 VSS.n17017 VSS.n17016 0.00942857
R23358 VSS.n17089 VSS.n16947 0.00942857
R23359 VSS.n16950 VSS.n16948 0.00942857
R23360 VSS.n1100 VSS.n1090 0.00942857
R23361 VSS.n18034 VSS.n18033 0.00942857
R23362 VSS.n1069 VSS.n1060 0.00942857
R23363 VSS.n1099 VSS.n1098 0.00942857
R23364 VSS.n18024 VSS.n1039 0.00942857
R23365 VSS.n1129 VSS.n1052 0.00942857
R23366 VSS.n1145 VSS.n1058 0.00942857
R23367 VSS.n17182 VSS.n16903 0.00942857
R23368 VSS.n17187 VSS.n17186 0.00942857
R23369 VSS.n17198 VSS.n17196 0.00942857
R23370 VSS.n17242 VSS.n16878 0.00942857
R23371 VSS.n17256 VSS.n16871 0.00942857
R23372 VSS.n16877 VSS.n16872 0.00942857
R23373 VSS.n17015 VSS.n16998 0.00942857
R23374 VSS.n17036 VSS.n16984 0.00942857
R23375 VSS.n17063 VSS.n17062 0.00942857
R23376 VSS.n16949 VSS.n16943 0.00942857
R23377 VSS.n17609 VSS.n17608 0.00942857
R23378 VSS.n17681 VSS.n17361 0.00942857
R23379 VSS.n17364 VSS.n17362 0.00942857
R23380 VSS.n17519 VSS.n17484 0.00942857
R23381 VSS.n17488 VSS.n17487 0.00942857
R23382 VSS.n17581 VSS.n17580 0.00942857
R23383 VSS.n17507 VSS.n17485 0.00942857
R23384 VSS.n17544 VSS.n17467 0.00942857
R23385 VSS.n17452 VSS.n17442 0.00942857
R23386 VSS.n17579 VSS.n17433 0.00942857
R23387 VSS.n17774 VSS.n17317 0.00942857
R23388 VSS.n17779 VSS.n17778 0.00942857
R23389 VSS.n17790 VSS.n17788 0.00942857
R23390 VSS.n17834 VSS.n17292 0.00942857
R23391 VSS.n17848 VSS.n17285 0.00942857
R23392 VSS.n17291 VSS.n17286 0.00942857
R23393 VSS.n17607 VSS.n17412 0.00942857
R23394 VSS.n17628 VSS.n17398 0.00942857
R23395 VSS.n17655 VSS.n17654 0.00942857
R23396 VSS.n17363 VSS.n17357 0.00942857
R23397 VSS.n18096 VSS.n276 0.00942857
R23398 VSS.n280 VSS.n279 0.00942857
R23399 VSS.n18158 VSS.n18157 0.00942857
R23400 VSS.n18244 VSS.n18243 0.00942857
R23401 VSS.n18550 VSS.n18549 0.00942857
R23402 VSS.n18294 VSS.n18293 0.00942857
R23403 VSS.n18242 VSS.n18241 0.00942857
R23404 VSS.n18255 VSS.n18184 0.00942857
R23405 VSS.n18198 VSS.n18195 0.00942857
R23406 VSS.n18295 VSS.n18221 0.00942857
R23407 VSS.n18377 VSS.n18376 0.00942857
R23408 VSS.n18500 VSS.n18355 0.00942857
R23409 VSS.n18403 VSS.n18394 0.00942857
R23410 VSS.n18482 VSS.n18419 0.00942857
R23411 VSS.n18478 VSS.n18423 0.00942857
R23412 VSS.n18477 VSS.n18476 0.00942857
R23413 VSS.n18084 VSS.n277 0.00942857
R23414 VSS.n18121 VSS.n259 0.00942857
R23415 VSS.n244 VSS.n234 0.00942857
R23416 VSS.n18156 VSS.n225 0.00942857
R23417 VSS.n9569 VSS.n9534 0.00942857
R23418 VSS.n9538 VSS.n9537 0.00942857
R23419 VSS.n9631 VSS.n9630 0.00942857
R23420 VSS.n9659 VSS.n9658 0.00942857
R23421 VSS.n9731 VSS.n9411 0.00942857
R23422 VSS.n9414 VSS.n9412 0.00942857
R23423 VSS.n9657 VSS.n9462 0.00942857
R23424 VSS.n9678 VSS.n9448 0.00942857
R23425 VSS.n9705 VSS.n9704 0.00942857
R23426 VSS.n9413 VSS.n9407 0.00942857
R23427 VSS.n9824 VSS.n9367 0.00942857
R23428 VSS.n9829 VSS.n9828 0.00942857
R23429 VSS.n9840 VSS.n9838 0.00942857
R23430 VSS.n9884 VSS.n9342 0.00942857
R23431 VSS.n9899 VSS.n9336 0.00942857
R23432 VSS.n9898 VSS.n9338 0.00942857
R23433 VSS.n9557 VSS.n9535 0.00942857
R23434 VSS.n9594 VSS.n9517 0.00942857
R23435 VSS.n9502 VSS.n9492 0.00942857
R23436 VSS.n9629 VSS.n9483 0.00942857
R23437 VSS.n16505 VSS.n16472 0.00942857
R23438 VSS.n16475 VSS.n16474 0.00942857
R23439 VSS.n16575 VSS.n16423 0.00942857
R23440 VSS.n16602 VSS.n16601 0.00942857
R23441 VSS.n16674 VSS.n16353 0.00942857
R23442 VSS.n16356 VSS.n16354 0.00942857
R23443 VSS.n16600 VSS.n16404 0.00942857
R23444 VSS.n16621 VSS.n16390 0.00942857
R23445 VSS.n16648 VSS.n16647 0.00942857
R23446 VSS.n16355 VSS.n16349 0.00942857
R23447 VSS.n16767 VSS.n16309 0.00942857
R23448 VSS.n16772 VSS.n16771 0.00942857
R23449 VSS.n16783 VSS.n16781 0.00942857
R23450 VSS.n16827 VSS.n16284 0.00942857
R23451 VSS.n16842 VSS.n16278 0.00942857
R23452 VSS.n16841 VSS.n16280 0.00942857
R23453 VSS.n16493 VSS.n16473 0.00942857
R23454 VSS.n16519 VSS.n16448 0.00942857
R23455 VSS.n16555 VSS.n16554 0.00942857
R23456 VSS.n16577 VSS.n16576 0.00942857
R23457 VSS.n1670 VSS.n1637 0.00942857
R23458 VSS.n1640 VSS.n1639 0.00942857
R23459 VSS.n1740 VSS.n1588 0.00942857
R23460 VSS.n16009 VSS.n16008 0.00942857
R23461 VSS.n16081 VSS.n1525 0.00942857
R23462 VSS.n1528 VSS.n1526 0.00942857
R23463 VSS.n16007 VSS.n1576 0.00942857
R23464 VSS.n16028 VSS.n1562 0.00942857
R23465 VSS.n16055 VSS.n16054 0.00942857
R23466 VSS.n1527 VSS.n1521 0.00942857
R23467 VSS.n16174 VSS.n1481 0.00942857
R23468 VSS.n16179 VSS.n16178 0.00942857
R23469 VSS.n16190 VSS.n16188 0.00942857
R23470 VSS.n16234 VSS.n1456 0.00942857
R23471 VSS.n16249 VSS.n1450 0.00942857
R23472 VSS.n16248 VSS.n1452 0.00942857
R23473 VSS.n1658 VSS.n1638 0.00942857
R23474 VSS.n1684 VSS.n1613 0.00942857
R23475 VSS.n1720 VSS.n1719 0.00942857
R23476 VSS.n1742 VSS.n1741 0.00942857
R23477 VSS.n1861 VSS.n1826 0.00942857
R23478 VSS.n1830 VSS.n1829 0.00942857
R23479 VSS.n1923 VSS.n1922 0.00942857
R23480 VSS.n2009 VSS.n2008 0.00942857
R23481 VSS.n2315 VSS.n2314 0.00942857
R23482 VSS.n2059 VSS.n2058 0.00942857
R23483 VSS.n2007 VSS.n2006 0.00942857
R23484 VSS.n2020 VSS.n1949 0.00942857
R23485 VSS.n1963 VSS.n1960 0.00942857
R23486 VSS.n2060 VSS.n1986 0.00942857
R23487 VSS.n2142 VSS.n2133 0.00942857
R23488 VSS.n2147 VSS.n2146 0.00942857
R23489 VSS.n2181 VSS.n2180 0.00942857
R23490 VSS.n2171 VSS.n2163 0.00942857
R23491 VSS.n2234 VSS.n2172 0.00942857
R23492 VSS.n2209 VSS.n2170 0.00942857
R23493 VSS.n1849 VSS.n1827 0.00942857
R23494 VSS.n1886 VSS.n1809 0.00942857
R23495 VSS.n1794 VSS.n1784 0.00942857
R23496 VSS.n1921 VSS.n1775 0.00942857
R23497 VSS.n3060 VSS.n3025 0.00942857
R23498 VSS.n3029 VSS.n3028 0.00942857
R23499 VSS.n3122 VSS.n3121 0.00942857
R23500 VSS.n3150 VSS.n3149 0.00942857
R23501 VSS.n3222 VSS.n2902 0.00942857
R23502 VSS.n2905 VSS.n2903 0.00942857
R23503 VSS.n3148 VSS.n2953 0.00942857
R23504 VSS.n3169 VSS.n2939 0.00942857
R23505 VSS.n3196 VSS.n3195 0.00942857
R23506 VSS.n2904 VSS.n2898 0.00942857
R23507 VSS.n3315 VSS.n2858 0.00942857
R23508 VSS.n3320 VSS.n3319 0.00942857
R23509 VSS.n3331 VSS.n3329 0.00942857
R23510 VSS.n3375 VSS.n2833 0.00942857
R23511 VSS.n3390 VSS.n2827 0.00942857
R23512 VSS.n3389 VSS.n2829 0.00942857
R23513 VSS.n3048 VSS.n3026 0.00942857
R23514 VSS.n3085 VSS.n3008 0.00942857
R23515 VSS.n2993 VSS.n2983 0.00942857
R23516 VSS.n3120 VSS.n2974 0.00942857
R23517 VSS.n3652 VSS.n3617 0.00942857
R23518 VSS.n3621 VSS.n3620 0.00942857
R23519 VSS.n3714 VSS.n3713 0.00942857
R23520 VSS.n3742 VSS.n3741 0.00942857
R23521 VSS.n3814 VSS.n3494 0.00942857
R23522 VSS.n3497 VSS.n3495 0.00942857
R23523 VSS.n3740 VSS.n3545 0.00942857
R23524 VSS.n3761 VSS.n3531 0.00942857
R23525 VSS.n3788 VSS.n3787 0.00942857
R23526 VSS.n3496 VSS.n3490 0.00942857
R23527 VSS.n3907 VSS.n3450 0.00942857
R23528 VSS.n3912 VSS.n3911 0.00942857
R23529 VSS.n3923 VSS.n3921 0.00942857
R23530 VSS.n3967 VSS.n3425 0.00942857
R23531 VSS.n3982 VSS.n3419 0.00942857
R23532 VSS.n3981 VSS.n3421 0.00942857
R23533 VSS.n3640 VSS.n3618 0.00942857
R23534 VSS.n3677 VSS.n3600 0.00942857
R23535 VSS.n3585 VSS.n3575 0.00942857
R23536 VSS.n3712 VSS.n3566 0.00942857
R23537 VSS.n4244 VSS.n4209 0.00942857
R23538 VSS.n4213 VSS.n4212 0.00942857
R23539 VSS.n4306 VSS.n4305 0.00942857
R23540 VSS.n4334 VSS.n4333 0.00942857
R23541 VSS.n4406 VSS.n4086 0.00942857
R23542 VSS.n4089 VSS.n4087 0.00942857
R23543 VSS.n4332 VSS.n4137 0.00942857
R23544 VSS.n4353 VSS.n4123 0.00942857
R23545 VSS.n4380 VSS.n4379 0.00942857
R23546 VSS.n4088 VSS.n4082 0.00942857
R23547 VSS.n4499 VSS.n4042 0.00942857
R23548 VSS.n4504 VSS.n4503 0.00942857
R23549 VSS.n4515 VSS.n4513 0.00942857
R23550 VSS.n4559 VSS.n4017 0.00942857
R23551 VSS.n4574 VSS.n4011 0.00942857
R23552 VSS.n4573 VSS.n4013 0.00942857
R23553 VSS.n4232 VSS.n4210 0.00942857
R23554 VSS.n4269 VSS.n4192 0.00942857
R23555 VSS.n4177 VSS.n4167 0.00942857
R23556 VSS.n4304 VSS.n4158 0.00942857
R23557 VSS.n4836 VSS.n4801 0.00942857
R23558 VSS.n4805 VSS.n4804 0.00942857
R23559 VSS.n4898 VSS.n4897 0.00942857
R23560 VSS.n4926 VSS.n4925 0.00942857
R23561 VSS.n4998 VSS.n4678 0.00942857
R23562 VSS.n4681 VSS.n4679 0.00942857
R23563 VSS.n4924 VSS.n4729 0.00942857
R23564 VSS.n4945 VSS.n4715 0.00942857
R23565 VSS.n4972 VSS.n4971 0.00942857
R23566 VSS.n4680 VSS.n4674 0.00942857
R23567 VSS.n5091 VSS.n4634 0.00942857
R23568 VSS.n5096 VSS.n5095 0.00942857
R23569 VSS.n5107 VSS.n5105 0.00942857
R23570 VSS.n5151 VSS.n4609 0.00942857
R23571 VSS.n5166 VSS.n4603 0.00942857
R23572 VSS.n5165 VSS.n4605 0.00942857
R23573 VSS.n4824 VSS.n4802 0.00942857
R23574 VSS.n4861 VSS.n4784 0.00942857
R23575 VSS.n4769 VSS.n4759 0.00942857
R23576 VSS.n4896 VSS.n4750 0.00942857
R23577 VSS.n2457 VSS.n2422 0.00942857
R23578 VSS.n2426 VSS.n2425 0.00942857
R23579 VSS.n2519 VSS.n2518 0.00942857
R23580 VSS.n2605 VSS.n2604 0.00942857
R23581 VSS.n5280 VSS.n5279 0.00942857
R23582 VSS.n2655 VSS.n2654 0.00942857
R23583 VSS.n2603 VSS.n2602 0.00942857
R23584 VSS.n2616 VSS.n2545 0.00942857
R23585 VSS.n2559 VSS.n2556 0.00942857
R23586 VSS.n2656 VSS.n2582 0.00942857
R23587 VSS.n2738 VSS.n2729 0.00942857
R23588 VSS.n2743 VSS.n2742 0.00942857
R23589 VSS.n2777 VSS.n2776 0.00942857
R23590 VSS.n2767 VSS.n2759 0.00942857
R23591 VSS.n5199 VSS.n2768 0.00942857
R23592 VSS.n2805 VSS.n2766 0.00942857
R23593 VSS.n2445 VSS.n2423 0.00942857
R23594 VSS.n2482 VSS.n2405 0.00942857
R23595 VSS.n2390 VSS.n2380 0.00942857
R23596 VSS.n2517 VSS.n2371 0.00942857
R23597 VSS.n5418 VSS.n5383 0.00942857
R23598 VSS.n5387 VSS.n5386 0.00942857
R23599 VSS.n5480 VSS.n5479 0.00942857
R23600 VSS.n5566 VSS.n5565 0.00942857
R23601 VSS.n5853 VSS.n5852 0.00942857
R23602 VSS.n5616 VSS.n5615 0.00942857
R23603 VSS.n5564 VSS.n5563 0.00942857
R23604 VSS.n5577 VSS.n5506 0.00942857
R23605 VSS.n5520 VSS.n5517 0.00942857
R23606 VSS.n5617 VSS.n5543 0.00942857
R23607 VSS.n5699 VSS.n5690 0.00942857
R23608 VSS.n5704 VSS.n5703 0.00942857
R23609 VSS.n5751 VSS.n5750 0.00942857
R23610 VSS.n5728 VSS.n5720 0.00942857
R23611 VSS.n5772 VSS.n5741 0.00942857
R23612 VSS.n5740 VSS.n5727 0.00942857
R23613 VSS.n5406 VSS.n5384 0.00942857
R23614 VSS.n5443 VSS.n5366 0.00942857
R23615 VSS.n5351 VSS.n5341 0.00942857
R23616 VSS.n5478 VSS.n5332 0.00942857
R23617 VSS.n5991 VSS.n5956 0.00942857
R23618 VSS.n5960 VSS.n5959 0.00942857
R23619 VSS.n6053 VSS.n6052 0.00942857
R23620 VSS.n6139 VSS.n6138 0.00942857
R23621 VSS.n6445 VSS.n6444 0.00942857
R23622 VSS.n6189 VSS.n6188 0.00942857
R23623 VSS.n6137 VSS.n6136 0.00942857
R23624 VSS.n6150 VSS.n6079 0.00942857
R23625 VSS.n6093 VSS.n6090 0.00942857
R23626 VSS.n6190 VSS.n6116 0.00942857
R23627 VSS.n6272 VSS.n6263 0.00942857
R23628 VSS.n6277 VSS.n6276 0.00942857
R23629 VSS.n6311 VSS.n6310 0.00942857
R23630 VSS.n6301 VSS.n6293 0.00942857
R23631 VSS.n6364 VSS.n6302 0.00942857
R23632 VSS.n6339 VSS.n6300 0.00942857
R23633 VSS.n5979 VSS.n5957 0.00942857
R23634 VSS.n6016 VSS.n5939 0.00942857
R23635 VSS.n5924 VSS.n5914 0.00942857
R23636 VSS.n6051 VSS.n5905 0.00942857
R23637 VSS.n7793 VSS.n7758 0.00942857
R23638 VSS.n7762 VSS.n7761 0.00942857
R23639 VSS.n7855 VSS.n7854 0.00942857
R23640 VSS.n7883 VSS.n7882 0.00942857
R23641 VSS.n7955 VSS.n7635 0.00942857
R23642 VSS.n7638 VSS.n7636 0.00942857
R23643 VSS.n7881 VSS.n7686 0.00942857
R23644 VSS.n7902 VSS.n7672 0.00942857
R23645 VSS.n7929 VSS.n7928 0.00942857
R23646 VSS.n7637 VSS.n7631 0.00942857
R23647 VSS.n8048 VSS.n7591 0.00942857
R23648 VSS.n8053 VSS.n8052 0.00942857
R23649 VSS.n8064 VSS.n8062 0.00942857
R23650 VSS.n8108 VSS.n7566 0.00942857
R23651 VSS.n8123 VSS.n7560 0.00942857
R23652 VSS.n8122 VSS.n7562 0.00942857
R23653 VSS.n7781 VSS.n7759 0.00942857
R23654 VSS.n7818 VSS.n7741 0.00942857
R23655 VSS.n7726 VSS.n7716 0.00942857
R23656 VSS.n7853 VSS.n7707 0.00942857
R23657 VSS.n8385 VSS.n8350 0.00942857
R23658 VSS.n8354 VSS.n8353 0.00942857
R23659 VSS.n8447 VSS.n8446 0.00942857
R23660 VSS.n8475 VSS.n8474 0.00942857
R23661 VSS.n8547 VSS.n8227 0.00942857
R23662 VSS.n8230 VSS.n8228 0.00942857
R23663 VSS.n8473 VSS.n8278 0.00942857
R23664 VSS.n8494 VSS.n8264 0.00942857
R23665 VSS.n8521 VSS.n8520 0.00942857
R23666 VSS.n8229 VSS.n8223 0.00942857
R23667 VSS.n8640 VSS.n8183 0.00942857
R23668 VSS.n8645 VSS.n8644 0.00942857
R23669 VSS.n8656 VSS.n8654 0.00942857
R23670 VSS.n8700 VSS.n8158 0.00942857
R23671 VSS.n8715 VSS.n8152 0.00942857
R23672 VSS.n8714 VSS.n8154 0.00942857
R23673 VSS.n8373 VSS.n8351 0.00942857
R23674 VSS.n8410 VSS.n8333 0.00942857
R23675 VSS.n8318 VSS.n8308 0.00942857
R23676 VSS.n8445 VSS.n8299 0.00942857
R23677 VSS.n8977 VSS.n8942 0.00942857
R23678 VSS.n8946 VSS.n8945 0.00942857
R23679 VSS.n9039 VSS.n9038 0.00942857
R23680 VSS.n9067 VSS.n9066 0.00942857
R23681 VSS.n9139 VSS.n8819 0.00942857
R23682 VSS.n8822 VSS.n8820 0.00942857
R23683 VSS.n9065 VSS.n8870 0.00942857
R23684 VSS.n9086 VSS.n8856 0.00942857
R23685 VSS.n9113 VSS.n9112 0.00942857
R23686 VSS.n8821 VSS.n8815 0.00942857
R23687 VSS.n9232 VSS.n8775 0.00942857
R23688 VSS.n9237 VSS.n9236 0.00942857
R23689 VSS.n9248 VSS.n9246 0.00942857
R23690 VSS.n9292 VSS.n8750 0.00942857
R23691 VSS.n9307 VSS.n8744 0.00942857
R23692 VSS.n9306 VSS.n8746 0.00942857
R23693 VSS.n8965 VSS.n8943 0.00942857
R23694 VSS.n9002 VSS.n8925 0.00942857
R23695 VSS.n8910 VSS.n8900 0.00942857
R23696 VSS.n9037 VSS.n8891 0.00942857
R23697 VSS.n10161 VSS.n10126 0.00942857
R23698 VSS.n10130 VSS.n10129 0.00942857
R23699 VSS.n10223 VSS.n10222 0.00942857
R23700 VSS.n10251 VSS.n10250 0.00942857
R23701 VSS.n10323 VSS.n10003 0.00942857
R23702 VSS.n10006 VSS.n10004 0.00942857
R23703 VSS.n10249 VSS.n10054 0.00942857
R23704 VSS.n10270 VSS.n10040 0.00942857
R23705 VSS.n10297 VSS.n10296 0.00942857
R23706 VSS.n10005 VSS.n9999 0.00942857
R23707 VSS.n10416 VSS.n9959 0.00942857
R23708 VSS.n10421 VSS.n10420 0.00942857
R23709 VSS.n10432 VSS.n10430 0.00942857
R23710 VSS.n10476 VSS.n9934 0.00942857
R23711 VSS.n10491 VSS.n9928 0.00942857
R23712 VSS.n10490 VSS.n9930 0.00942857
R23713 VSS.n10149 VSS.n10127 0.00942857
R23714 VSS.n10186 VSS.n10109 0.00942857
R23715 VSS.n10094 VSS.n10084 0.00942857
R23716 VSS.n10221 VSS.n10075 0.00942857
R23717 VSS.n10753 VSS.n10718 0.00942857
R23718 VSS.n10722 VSS.n10721 0.00942857
R23719 VSS.n10815 VSS.n10814 0.00942857
R23720 VSS.n10843 VSS.n10842 0.00942857
R23721 VSS.n10915 VSS.n10595 0.00942857
R23722 VSS.n10598 VSS.n10596 0.00942857
R23723 VSS.n10841 VSS.n10646 0.00942857
R23724 VSS.n10862 VSS.n10632 0.00942857
R23725 VSS.n10889 VSS.n10888 0.00942857
R23726 VSS.n10597 VSS.n10591 0.00942857
R23727 VSS.n11008 VSS.n10551 0.00942857
R23728 VSS.n11013 VSS.n11012 0.00942857
R23729 VSS.n11024 VSS.n11022 0.00942857
R23730 VSS.n11068 VSS.n10526 0.00942857
R23731 VSS.n11083 VSS.n10520 0.00942857
R23732 VSS.n11082 VSS.n10522 0.00942857
R23733 VSS.n10741 VSS.n10719 0.00942857
R23734 VSS.n10778 VSS.n10701 0.00942857
R23735 VSS.n10686 VSS.n10676 0.00942857
R23736 VSS.n10813 VSS.n10667 0.00942857
R23737 VSS.n11345 VSS.n11310 0.00942857
R23738 VSS.n11314 VSS.n11313 0.00942857
R23739 VSS.n11407 VSS.n11406 0.00942857
R23740 VSS.n11435 VSS.n11434 0.00942857
R23741 VSS.n11507 VSS.n11187 0.00942857
R23742 VSS.n11190 VSS.n11188 0.00942857
R23743 VSS.n11433 VSS.n11238 0.00942857
R23744 VSS.n11454 VSS.n11224 0.00942857
R23745 VSS.n11481 VSS.n11480 0.00942857
R23746 VSS.n11189 VSS.n11183 0.00942857
R23747 VSS.n11600 VSS.n11143 0.00942857
R23748 VSS.n11605 VSS.n11604 0.00942857
R23749 VSS.n11616 VSS.n11614 0.00942857
R23750 VSS.n11660 VSS.n11118 0.00942857
R23751 VSS.n11675 VSS.n11112 0.00942857
R23752 VSS.n11674 VSS.n11114 0.00942857
R23753 VSS.n11333 VSS.n11311 0.00942857
R23754 VSS.n11370 VSS.n11293 0.00942857
R23755 VSS.n11278 VSS.n11268 0.00942857
R23756 VSS.n11405 VSS.n11259 0.00942857
R23757 VSS.n11937 VSS.n11902 0.00942857
R23758 VSS.n11906 VSS.n11905 0.00942857
R23759 VSS.n11999 VSS.n11998 0.00942857
R23760 VSS.n12027 VSS.n12026 0.00942857
R23761 VSS.n12099 VSS.n11779 0.00942857
R23762 VSS.n11782 VSS.n11780 0.00942857
R23763 VSS.n12025 VSS.n11830 0.00942857
R23764 VSS.n12046 VSS.n11816 0.00942857
R23765 VSS.n12073 VSS.n12072 0.00942857
R23766 VSS.n11781 VSS.n11775 0.00942857
R23767 VSS.n12192 VSS.n11735 0.00942857
R23768 VSS.n12197 VSS.n12196 0.00942857
R23769 VSS.n12208 VSS.n12206 0.00942857
R23770 VSS.n12252 VSS.n11710 0.00942857
R23771 VSS.n12267 VSS.n11704 0.00942857
R23772 VSS.n12266 VSS.n11706 0.00942857
R23773 VSS.n11925 VSS.n11903 0.00942857
R23774 VSS.n11962 VSS.n11885 0.00942857
R23775 VSS.n11870 VSS.n11860 0.00942857
R23776 VSS.n11997 VSS.n11851 0.00942857
R23777 VSS.n12529 VSS.n12494 0.00942857
R23778 VSS.n12498 VSS.n12497 0.00942857
R23779 VSS.n12591 VSS.n12590 0.00942857
R23780 VSS.n12619 VSS.n12618 0.00942857
R23781 VSS.n12691 VSS.n12371 0.00942857
R23782 VSS.n12374 VSS.n12372 0.00942857
R23783 VSS.n12617 VSS.n12422 0.00942857
R23784 VSS.n12638 VSS.n12408 0.00942857
R23785 VSS.n12665 VSS.n12664 0.00942857
R23786 VSS.n12373 VSS.n12367 0.00942857
R23787 VSS.n12784 VSS.n12327 0.00942857
R23788 VSS.n12789 VSS.n12788 0.00942857
R23789 VSS.n12800 VSS.n12798 0.00942857
R23790 VSS.n12844 VSS.n12302 0.00942857
R23791 VSS.n12859 VSS.n12296 0.00942857
R23792 VSS.n12858 VSS.n12298 0.00942857
R23793 VSS.n12517 VSS.n12495 0.00942857
R23794 VSS.n12554 VSS.n12477 0.00942857
R23795 VSS.n12462 VSS.n12452 0.00942857
R23796 VSS.n12589 VSS.n12443 0.00942857
R23797 VSS.n13121 VSS.n13086 0.00942857
R23798 VSS.n13090 VSS.n13089 0.00942857
R23799 VSS.n13183 VSS.n13182 0.00942857
R23800 VSS.n13211 VSS.n13210 0.00942857
R23801 VSS.n13283 VSS.n12963 0.00942857
R23802 VSS.n12966 VSS.n12964 0.00942857
R23803 VSS.n13209 VSS.n13014 0.00942857
R23804 VSS.n13230 VSS.n13000 0.00942857
R23805 VSS.n13257 VSS.n13256 0.00942857
R23806 VSS.n12965 VSS.n12959 0.00942857
R23807 VSS.n13376 VSS.n12919 0.00942857
R23808 VSS.n13381 VSS.n13380 0.00942857
R23809 VSS.n13392 VSS.n13390 0.00942857
R23810 VSS.n13436 VSS.n12894 0.00942857
R23811 VSS.n13451 VSS.n12888 0.00942857
R23812 VSS.n13450 VSS.n12890 0.00942857
R23813 VSS.n13109 VSS.n13087 0.00942857
R23814 VSS.n13146 VSS.n13069 0.00942857
R23815 VSS.n13054 VSS.n13044 0.00942857
R23816 VSS.n13181 VSS.n13035 0.00942857
R23817 VSS.n13713 VSS.n13678 0.00942857
R23818 VSS.n13682 VSS.n13681 0.00942857
R23819 VSS.n13775 VSS.n13774 0.00942857
R23820 VSS.n13803 VSS.n13802 0.00942857
R23821 VSS.n13875 VSS.n13555 0.00942857
R23822 VSS.n13558 VSS.n13556 0.00942857
R23823 VSS.n13801 VSS.n13606 0.00942857
R23824 VSS.n13822 VSS.n13592 0.00942857
R23825 VSS.n13849 VSS.n13848 0.00942857
R23826 VSS.n13557 VSS.n13551 0.00942857
R23827 VSS.n13968 VSS.n13511 0.00942857
R23828 VSS.n13973 VSS.n13972 0.00942857
R23829 VSS.n13984 VSS.n13982 0.00942857
R23830 VSS.n14028 VSS.n13486 0.00942857
R23831 VSS.n14043 VSS.n13480 0.00942857
R23832 VSS.n14042 VSS.n13482 0.00942857
R23833 VSS.n13701 VSS.n13679 0.00942857
R23834 VSS.n13738 VSS.n13661 0.00942857
R23835 VSS.n13646 VSS.n13636 0.00942857
R23836 VSS.n13773 VSS.n13627 0.00942857
R23837 VSS.n14305 VSS.n14270 0.00942857
R23838 VSS.n14274 VSS.n14273 0.00942857
R23839 VSS.n14367 VSS.n14366 0.00942857
R23840 VSS.n14395 VSS.n14394 0.00942857
R23841 VSS.n14467 VSS.n14147 0.00942857
R23842 VSS.n14150 VSS.n14148 0.00942857
R23843 VSS.n14393 VSS.n14198 0.00942857
R23844 VSS.n14414 VSS.n14184 0.00942857
R23845 VSS.n14441 VSS.n14440 0.00942857
R23846 VSS.n14149 VSS.n14143 0.00942857
R23847 VSS.n14560 VSS.n14103 0.00942857
R23848 VSS.n14565 VSS.n14564 0.00942857
R23849 VSS.n14576 VSS.n14574 0.00942857
R23850 VSS.n14620 VSS.n14078 0.00942857
R23851 VSS.n14635 VSS.n14072 0.00942857
R23852 VSS.n14634 VSS.n14074 0.00942857
R23853 VSS.n14293 VSS.n14271 0.00942857
R23854 VSS.n14330 VSS.n14253 0.00942857
R23855 VSS.n14238 VSS.n14228 0.00942857
R23856 VSS.n14365 VSS.n14219 0.00942857
R23857 VSS.n14897 VSS.n14862 0.00942857
R23858 VSS.n14866 VSS.n14865 0.00942857
R23859 VSS.n14959 VSS.n14958 0.00942857
R23860 VSS.n14987 VSS.n14986 0.00942857
R23861 VSS.n15059 VSS.n14739 0.00942857
R23862 VSS.n14742 VSS.n14740 0.00942857
R23863 VSS.n14985 VSS.n14790 0.00942857
R23864 VSS.n15006 VSS.n14776 0.00942857
R23865 VSS.n15033 VSS.n15032 0.00942857
R23866 VSS.n14741 VSS.n14735 0.00942857
R23867 VSS.n15152 VSS.n14695 0.00942857
R23868 VSS.n15157 VSS.n15156 0.00942857
R23869 VSS.n15168 VSS.n15166 0.00942857
R23870 VSS.n15212 VSS.n14670 0.00942857
R23871 VSS.n15227 VSS.n14664 0.00942857
R23872 VSS.n15226 VSS.n14666 0.00942857
R23873 VSS.n14885 VSS.n14863 0.00942857
R23874 VSS.n14922 VSS.n14845 0.00942857
R23875 VSS.n14830 VSS.n14820 0.00942857
R23876 VSS.n14957 VSS.n14811 0.00942857
R23877 VSS.n15489 VSS.n15454 0.00942857
R23878 VSS.n15458 VSS.n15457 0.00942857
R23879 VSS.n15551 VSS.n15550 0.00942857
R23880 VSS.n15579 VSS.n15578 0.00942857
R23881 VSS.n15651 VSS.n15331 0.00942857
R23882 VSS.n15334 VSS.n15332 0.00942857
R23883 VSS.n15577 VSS.n15382 0.00942857
R23884 VSS.n15598 VSS.n15368 0.00942857
R23885 VSS.n15625 VSS.n15624 0.00942857
R23886 VSS.n15333 VSS.n15327 0.00942857
R23887 VSS.n15744 VSS.n15287 0.00942857
R23888 VSS.n15749 VSS.n15748 0.00942857
R23889 VSS.n15760 VSS.n15758 0.00942857
R23890 VSS.n15804 VSS.n15262 0.00942857
R23891 VSS.n15819 VSS.n15256 0.00942857
R23892 VSS.n15818 VSS.n15258 0.00942857
R23893 VSS.n15477 VSS.n15455 0.00942857
R23894 VSS.n15514 VSS.n15437 0.00942857
R23895 VSS.n15422 VSS.n15412 0.00942857
R23896 VSS.n15549 VSS.n15403 0.00942857
R23897 VSS.n6597 VSS.n6562 0.00942857
R23898 VSS.n6566 VSS.n6565 0.00942857
R23899 VSS.n6659 VSS.n6658 0.00942857
R23900 VSS.n6745 VSS.n6744 0.00942857
R23901 VSS.n15933 VSS.n15932 0.00942857
R23902 VSS.n6795 VSS.n6794 0.00942857
R23903 VSS.n6743 VSS.n6742 0.00942857
R23904 VSS.n6756 VSS.n6685 0.00942857
R23905 VSS.n6699 VSS.n6696 0.00942857
R23906 VSS.n6796 VSS.n6722 0.00942857
R23907 VSS.n6878 VSS.n6869 0.00942857
R23908 VSS.n6883 VSS.n6882 0.00942857
R23909 VSS.n6917 VSS.n6916 0.00942857
R23910 VSS.n6907 VSS.n6899 0.00942857
R23911 VSS.n15852 VSS.n6908 0.00942857
R23912 VSS.n6945 VSS.n6906 0.00942857
R23913 VSS.n6585 VSS.n6563 0.00942857
R23914 VSS.n6622 VSS.n6545 0.00942857
R23915 VSS.n6530 VSS.n6520 0.00942857
R23916 VSS.n6657 VSS.n6511 0.00942857
R23917 VSS.n7194 VSS.n7161 0.00942857
R23918 VSS.n7164 VSS.n7163 0.00942857
R23919 VSS.n7264 VSS.n7112 0.00942857
R23920 VSS.n7291 VSS.n7290 0.00942857
R23921 VSS.n7363 VSS.n7042 0.00942857
R23922 VSS.n7045 VSS.n7043 0.00942857
R23923 VSS.n7289 VSS.n7093 0.00942857
R23924 VSS.n7310 VSS.n7079 0.00942857
R23925 VSS.n7337 VSS.n7336 0.00942857
R23926 VSS.n7044 VSS.n7038 0.00942857
R23927 VSS.n7456 VSS.n6998 0.00942857
R23928 VSS.n7461 VSS.n7460 0.00942857
R23929 VSS.n7472 VSS.n7470 0.00942857
R23930 VSS.n7516 VSS.n6973 0.00942857
R23931 VSS.n7531 VSS.n6967 0.00942857
R23932 VSS.n7530 VSS.n6969 0.00942857
R23933 VSS.n7182 VSS.n7162 0.00942857
R23934 VSS.n7208 VSS.n7137 0.00942857
R23935 VSS.n7244 VSS.n7243 0.00942857
R23936 VSS.n7266 VSS.n7265 0.00942857
R23937 VSS.n354 VSS.n346 0.00942857
R23938 VSS.n443 VSS.n442 0.00942857
R23939 VSS.n412 VSS.n411 0.00942857
R23940 VSS.n18603 VSS.n18602 0.00942857
R23941 VSS.n18675 VSS.n140 0.00942857
R23942 VSS.n143 VSS.n141 0.00942857
R23943 VSS.n18601 VSS.n191 0.00942857
R23944 VSS.n18622 VSS.n177 0.00942857
R23945 VSS.n18649 VSS.n18648 0.00942857
R23946 VSS.n142 VSS.n136 0.00942857
R23947 VSS.n18768 VSS.n96 0.00942857
R23948 VSS.n18773 VSS.n18772 0.00942857
R23949 VSS.n18784 VSS.n18782 0.00942857
R23950 VSS.n18828 VSS.n71 0.00942857
R23951 VSS.n18843 VSS.n65 0.00942857
R23952 VSS.n18842 VSS.n67 0.00942857
R23953 VSS.n353 VSS.n352 0.00942857
R23954 VSS.n433 VSS.n306 0.00942857
R23955 VSS.n390 VSS.n319 0.00942857
R23956 VSS.n413 VSS.n324 0.00942857
R23957 VSS.n568 VSS.n498 0.00942857
R23958 VSS.n847 VSS.n846 0.00942857
R23959 VSS.n618 VSS.n617 0.00942857
R23960 VSS.n567 VSS.n499 0.00942857
R23961 VSS.n579 VSS.n505 0.00942857
R23962 VSS.n519 VSS.n516 0.00942857
R23963 VSS.n619 VSS.n542 0.00942857
R23964 VSS.n701 VSS.n692 0.00942857
R23965 VSS.n706 VSS.n705 0.00942857
R23966 VSS.n749 VSS.n748 0.00942857
R23967 VSS.n730 VSS.n722 0.00942857
R23968 VSS.n766 VSS.n742 0.00942857
R23969 VSS.n741 VSS.n729 0.00942857
R23970 VSS.n918 VSS.n917 0.00942857
R23971 VSS.n998 VSS.n472 0.00942857
R23972 VSS.n948 VSS.n485 0.00942857
R23973 VSS.n964 VSS.n491 0.00942857
R23974 VSS.n1360 VSS.n1351 0.00942857
R23975 VSS.n1365 VSS.n1364 0.00942857
R23976 VSS.n1399 VSS.n1398 0.00942857
R23977 VSS.n1389 VSS.n1381 0.00942857
R23978 VSS.n17880 VSS.n1390 0.00942857
R23979 VSS.n1427 VSS.n1388 0.00942857
R23980 VSS.n1203 VSS.n1194 0.00853571
R23981 VSS.n1279 VSS.n1192 0.00853571
R23982 VSS.n1196 VSS.n1193 0.00853571
R23983 VSS.n913 VSS.n912 0.00853571
R23984 VSS.n924 VSS.n923 0.00853571
R23985 VSS.n17094 VSS.n16942 0.00853571
R23986 VSS.n1094 VSS.n1093 0.00853571
R23987 VSS.n1105 VSS.n1104 0.00853571
R23988 VSS.n18040 VSS.n18039 0.00853571
R23989 VSS.n1092 VSS.n1091 0.00853571
R23990 VSS.n1102 VSS.n1034 0.00853571
R23991 VSS.n17172 VSS.n17171 0.00853571
R23992 VSS.n17211 VSS.n16898 0.00853571
R23993 VSS.n17224 VSS.n17223 0.00853571
R23994 VSS.n17136 VSS.n16931 0.00853571
R23995 VSS.n17143 VSS.n16928 0.00853571
R23996 VSS.n17173 VSS.n16906 0.00853571
R23997 VSS.n17178 VSS.n17177 0.00853571
R23998 VSS.n17225 VSS.n16888 0.00853571
R23999 VSS.n17225 VSS.n16889 0.00853571
R24000 VSS.n17252 VSS.n16874 0.00853571
R24001 VSS.n17248 VSS.n16874 0.00853571
R24002 VSS.n17270 VSS.n16861 0.00853571
R24003 VSS.n17096 VSS.n17095 0.00853571
R24004 VSS.n17132 VSS.n16933 0.00853571
R24005 VSS.n17686 VSS.n17356 0.00853571
R24006 VSS.n17511 VSS.n17510 0.00853571
R24007 VSS.n17534 VSS.n17473 0.00853571
R24008 VSS.n17503 VSS.n17491 0.00853571
R24009 VSS.n17509 VSS.n17492 0.00853571
R24010 VSS.n17474 VSS.n17472 0.00853571
R24011 VSS.n17764 VSS.n17763 0.00853571
R24012 VSS.n17803 VSS.n17312 0.00853571
R24013 VSS.n17816 VSS.n17815 0.00853571
R24014 VSS.n17728 VSS.n17345 0.00853571
R24015 VSS.n17735 VSS.n17342 0.00853571
R24016 VSS.n17765 VSS.n17320 0.00853571
R24017 VSS.n17770 VSS.n17769 0.00853571
R24018 VSS.n17817 VSS.n17302 0.00853571
R24019 VSS.n17817 VSS.n17303 0.00853571
R24020 VSS.n17844 VSS.n17288 0.00853571
R24021 VSS.n17840 VSS.n17288 0.00853571
R24022 VSS.n17862 VSS.n17275 0.00853571
R24023 VSS.n17688 VSS.n17687 0.00853571
R24024 VSS.n17724 VSS.n17347 0.00853571
R24025 VSS.n18088 VSS.n18087 0.00853571
R24026 VSS.n18111 VSS.n265 0.00853571
R24027 VSS.n18220 VSS.n18211 0.00853571
R24028 VSS.n18296 VSS.n18209 0.00853571
R24029 VSS.n18213 VSS.n18210 0.00853571
R24030 VSS.n18508 VSS.n18342 0.00853571
R24031 VSS.n18402 VSS.n18401 0.00853571
R24032 VSS.n18488 VSS.n18389 0.00853571
R24033 VSS.n18330 VSS.n18326 0.00853571
R24034 VSS.n18335 VSS.n18319 0.00853571
R24035 VSS.n18349 VSS.n18348 0.00853571
R24036 VSS.n18505 VSS.n18346 0.00853571
R24037 VSS.n18487 VSS.n18390 0.00853571
R24038 VSS.n18487 VSS.n18391 0.00853571
R24039 VSS.n18471 VSS.n18427 0.00853571
R24040 VSS.n18431 VSS.n18427 0.00853571
R24041 VSS.n18467 VSS.n18466 0.00853571
R24042 VSS.n18080 VSS.n283 0.00853571
R24043 VSS.n18086 VSS.n284 0.00853571
R24044 VSS.n266 VSS.n264 0.00853571
R24045 VSS.n9561 VSS.n9560 0.00853571
R24046 VSS.n9584 VSS.n9523 0.00853571
R24047 VSS.n9736 VSS.n9406 0.00853571
R24048 VSS.n9738 VSS.n9737 0.00853571
R24049 VSS.n9774 VSS.n9397 0.00853571
R24050 VSS.n9814 VSS.n9813 0.00853571
R24051 VSS.n9853 VSS.n9362 0.00853571
R24052 VSS.n9866 VSS.n9865 0.00853571
R24053 VSS.n9778 VSS.n9395 0.00853571
R24054 VSS.n9785 VSS.n9392 0.00853571
R24055 VSS.n9815 VSS.n9370 0.00853571
R24056 VSS.n9820 VSS.n9819 0.00853571
R24057 VSS.n9867 VSS.n9352 0.00853571
R24058 VSS.n9867 VSS.n9353 0.00853571
R24059 VSS.n9890 VSS.n9339 0.00853571
R24060 VSS.n9891 VSS.n9890 0.00853571
R24061 VSS.n9913 VSS.n9326 0.00853571
R24062 VSS.n9553 VSS.n9541 0.00853571
R24063 VSS.n9559 VSS.n9542 0.00853571
R24064 VSS.n9524 VSS.n9522 0.00853571
R24065 VSS.n16497 VSS.n16496 0.00853571
R24066 VSS.n16515 VSS.n16514 0.00853571
R24067 VSS.n16679 VSS.n16348 0.00853571
R24068 VSS.n16681 VSS.n16680 0.00853571
R24069 VSS.n16717 VSS.n16339 0.00853571
R24070 VSS.n16757 VSS.n16756 0.00853571
R24071 VSS.n16796 VSS.n16304 0.00853571
R24072 VSS.n16809 VSS.n16808 0.00853571
R24073 VSS.n16721 VSS.n16337 0.00853571
R24074 VSS.n16728 VSS.n16334 0.00853571
R24075 VSS.n16758 VSS.n16312 0.00853571
R24076 VSS.n16763 VSS.n16762 0.00853571
R24077 VSS.n16810 VSS.n16294 0.00853571
R24078 VSS.n16810 VSS.n16295 0.00853571
R24079 VSS.n16833 VSS.n16281 0.00853571
R24080 VSS.n16834 VSS.n16833 0.00853571
R24081 VSS.n16856 VSS.n16268 0.00853571
R24082 VSS.n16489 VSS.n16478 0.00853571
R24083 VSS.n16495 VSS.n16479 0.00853571
R24084 VSS.n16524 VSS.n16462 0.00853571
R24085 VSS.n1662 VSS.n1661 0.00853571
R24086 VSS.n1680 VSS.n1679 0.00853571
R24087 VSS.n16086 VSS.n1520 0.00853571
R24088 VSS.n16088 VSS.n16087 0.00853571
R24089 VSS.n16124 VSS.n1511 0.00853571
R24090 VSS.n16164 VSS.n16163 0.00853571
R24091 VSS.n16203 VSS.n1476 0.00853571
R24092 VSS.n16216 VSS.n16215 0.00853571
R24093 VSS.n16128 VSS.n1509 0.00853571
R24094 VSS.n16135 VSS.n1506 0.00853571
R24095 VSS.n16165 VSS.n1484 0.00853571
R24096 VSS.n16170 VSS.n16169 0.00853571
R24097 VSS.n16217 VSS.n1466 0.00853571
R24098 VSS.n16217 VSS.n1467 0.00853571
R24099 VSS.n16240 VSS.n1453 0.00853571
R24100 VSS.n16241 VSS.n16240 0.00853571
R24101 VSS.n16263 VSS.n1440 0.00853571
R24102 VSS.n1654 VSS.n1643 0.00853571
R24103 VSS.n1660 VSS.n1644 0.00853571
R24104 VSS.n1689 VSS.n1627 0.00853571
R24105 VSS.n1853 VSS.n1852 0.00853571
R24106 VSS.n1876 VSS.n1815 0.00853571
R24107 VSS.n1985 VSS.n1976 0.00853571
R24108 VSS.n2061 VSS.n1974 0.00853571
R24109 VSS.n1978 VSS.n1975 0.00853571
R24110 VSS.n2271 VSS.n2270 0.00853571
R24111 VSS.n2259 VSS.n2128 0.00853571
R24112 VSS.n2247 VSS.n2156 0.00853571
R24113 VSS.n2094 VSS.n2090 0.00853571
R24114 VSS.n2099 VSS.n2084 0.00853571
R24115 VSS.n2272 VSS.n2111 0.00853571
R24116 VSS.n2138 VSS.n2137 0.00853571
R24117 VSS.n2166 VSS.n2160 0.00853571
R24118 VSS.n2246 VSS.n2160 0.00853571
R24119 VSS.n2217 VSS.n2215 0.00853571
R24120 VSS.n2217 VSS.n2216 0.00853571
R24121 VSS.n2222 VSS.n2202 0.00853571
R24122 VSS.n1845 VSS.n1833 0.00853571
R24123 VSS.n1851 VSS.n1834 0.00853571
R24124 VSS.n1816 VSS.n1814 0.00853571
R24125 VSS.n3052 VSS.n3051 0.00853571
R24126 VSS.n3075 VSS.n3014 0.00853571
R24127 VSS.n3227 VSS.n2897 0.00853571
R24128 VSS.n3229 VSS.n3228 0.00853571
R24129 VSS.n3265 VSS.n2888 0.00853571
R24130 VSS.n3305 VSS.n3304 0.00853571
R24131 VSS.n3344 VSS.n2853 0.00853571
R24132 VSS.n3357 VSS.n3356 0.00853571
R24133 VSS.n3269 VSS.n2886 0.00853571
R24134 VSS.n3276 VSS.n2883 0.00853571
R24135 VSS.n3306 VSS.n2861 0.00853571
R24136 VSS.n3311 VSS.n3310 0.00853571
R24137 VSS.n3358 VSS.n2843 0.00853571
R24138 VSS.n3358 VSS.n2844 0.00853571
R24139 VSS.n3381 VSS.n2830 0.00853571
R24140 VSS.n3382 VSS.n3381 0.00853571
R24141 VSS.n3404 VSS.n2817 0.00853571
R24142 VSS.n3044 VSS.n3032 0.00853571
R24143 VSS.n3050 VSS.n3033 0.00853571
R24144 VSS.n3015 VSS.n3013 0.00853571
R24145 VSS.n3644 VSS.n3643 0.00853571
R24146 VSS.n3667 VSS.n3606 0.00853571
R24147 VSS.n3819 VSS.n3489 0.00853571
R24148 VSS.n3821 VSS.n3820 0.00853571
R24149 VSS.n3857 VSS.n3480 0.00853571
R24150 VSS.n3897 VSS.n3896 0.00853571
R24151 VSS.n3936 VSS.n3445 0.00853571
R24152 VSS.n3949 VSS.n3948 0.00853571
R24153 VSS.n3861 VSS.n3478 0.00853571
R24154 VSS.n3868 VSS.n3475 0.00853571
R24155 VSS.n3898 VSS.n3453 0.00853571
R24156 VSS.n3903 VSS.n3902 0.00853571
R24157 VSS.n3950 VSS.n3435 0.00853571
R24158 VSS.n3950 VSS.n3436 0.00853571
R24159 VSS.n3973 VSS.n3422 0.00853571
R24160 VSS.n3974 VSS.n3973 0.00853571
R24161 VSS.n3996 VSS.n3409 0.00853571
R24162 VSS.n3636 VSS.n3624 0.00853571
R24163 VSS.n3642 VSS.n3625 0.00853571
R24164 VSS.n3607 VSS.n3605 0.00853571
R24165 VSS.n4236 VSS.n4235 0.00853571
R24166 VSS.n4259 VSS.n4198 0.00853571
R24167 VSS.n4411 VSS.n4081 0.00853571
R24168 VSS.n4413 VSS.n4412 0.00853571
R24169 VSS.n4449 VSS.n4072 0.00853571
R24170 VSS.n4489 VSS.n4488 0.00853571
R24171 VSS.n4528 VSS.n4037 0.00853571
R24172 VSS.n4541 VSS.n4540 0.00853571
R24173 VSS.n4453 VSS.n4070 0.00853571
R24174 VSS.n4460 VSS.n4067 0.00853571
R24175 VSS.n4490 VSS.n4045 0.00853571
R24176 VSS.n4495 VSS.n4494 0.00853571
R24177 VSS.n4542 VSS.n4027 0.00853571
R24178 VSS.n4542 VSS.n4028 0.00853571
R24179 VSS.n4565 VSS.n4014 0.00853571
R24180 VSS.n4566 VSS.n4565 0.00853571
R24181 VSS.n4588 VSS.n4001 0.00853571
R24182 VSS.n4228 VSS.n4216 0.00853571
R24183 VSS.n4234 VSS.n4217 0.00853571
R24184 VSS.n4199 VSS.n4197 0.00853571
R24185 VSS.n4828 VSS.n4827 0.00853571
R24186 VSS.n4851 VSS.n4790 0.00853571
R24187 VSS.n5003 VSS.n4673 0.00853571
R24188 VSS.n5005 VSS.n5004 0.00853571
R24189 VSS.n5041 VSS.n4664 0.00853571
R24190 VSS.n5081 VSS.n5080 0.00853571
R24191 VSS.n5120 VSS.n4629 0.00853571
R24192 VSS.n5133 VSS.n5132 0.00853571
R24193 VSS.n5045 VSS.n4662 0.00853571
R24194 VSS.n5052 VSS.n4659 0.00853571
R24195 VSS.n5082 VSS.n4637 0.00853571
R24196 VSS.n5087 VSS.n5086 0.00853571
R24197 VSS.n5134 VSS.n4619 0.00853571
R24198 VSS.n5134 VSS.n4620 0.00853571
R24199 VSS.n5157 VSS.n4606 0.00853571
R24200 VSS.n5158 VSS.n5157 0.00853571
R24201 VSS.n5180 VSS.n4593 0.00853571
R24202 VSS.n4820 VSS.n4808 0.00853571
R24203 VSS.n4826 VSS.n4809 0.00853571
R24204 VSS.n4791 VSS.n4789 0.00853571
R24205 VSS.n2449 VSS.n2448 0.00853571
R24206 VSS.n2472 VSS.n2411 0.00853571
R24207 VSS.n2581 VSS.n2572 0.00853571
R24208 VSS.n2657 VSS.n2570 0.00853571
R24209 VSS.n2574 VSS.n2571 0.00853571
R24210 VSS.n5236 VSS.n5235 0.00853571
R24211 VSS.n5224 VSS.n2724 0.00853571
R24212 VSS.n5212 VSS.n2752 0.00853571
R24213 VSS.n2690 VSS.n2686 0.00853571
R24214 VSS.n2695 VSS.n2680 0.00853571
R24215 VSS.n5237 VSS.n2707 0.00853571
R24216 VSS.n2734 VSS.n2733 0.00853571
R24217 VSS.n2762 VSS.n2756 0.00853571
R24218 VSS.n5211 VSS.n2756 0.00853571
R24219 VSS.n2813 VSS.n2811 0.00853571
R24220 VSS.n2813 VSS.n2812 0.00853571
R24221 VSS.n5187 VSS.n2798 0.00853571
R24222 VSS.n2441 VSS.n2429 0.00853571
R24223 VSS.n2447 VSS.n2430 0.00853571
R24224 VSS.n2412 VSS.n2410 0.00853571
R24225 VSS.n5410 VSS.n5409 0.00853571
R24226 VSS.n5433 VSS.n5372 0.00853571
R24227 VSS.n5542 VSS.n5533 0.00853571
R24228 VSS.n5618 VSS.n5531 0.00853571
R24229 VSS.n5535 VSS.n5532 0.00853571
R24230 VSS.n5809 VSS.n5808 0.00853571
R24231 VSS.n5797 VSS.n5685 0.00853571
R24232 VSS.n5785 VSS.n5713 0.00853571
R24233 VSS.n5651 VSS.n5647 0.00853571
R24234 VSS.n5656 VSS.n5641 0.00853571
R24235 VSS.n5810 VSS.n5668 0.00853571
R24236 VSS.n5695 VSS.n5694 0.00853571
R24237 VSS.n5723 VSS.n5717 0.00853571
R24238 VSS.n5784 VSS.n5717 0.00853571
R24239 VSS.n5732 VSS.n5730 0.00853571
R24240 VSS.n5733 VSS.n5732 0.00853571
R24241 VSS.n18886 VSS.n2 0.00853571
R24242 VSS.n5402 VSS.n5390 0.00853571
R24243 VSS.n5408 VSS.n5391 0.00853571
R24244 VSS.n5373 VSS.n5371 0.00853571
R24245 VSS.n5983 VSS.n5982 0.00853571
R24246 VSS.n6006 VSS.n5945 0.00853571
R24247 VSS.n6115 VSS.n6106 0.00853571
R24248 VSS.n6191 VSS.n6104 0.00853571
R24249 VSS.n6108 VSS.n6105 0.00853571
R24250 VSS.n6401 VSS.n6400 0.00853571
R24251 VSS.n6389 VSS.n6258 0.00853571
R24252 VSS.n6377 VSS.n6286 0.00853571
R24253 VSS.n6224 VSS.n6220 0.00853571
R24254 VSS.n6229 VSS.n6214 0.00853571
R24255 VSS.n6402 VSS.n6241 0.00853571
R24256 VSS.n6268 VSS.n6267 0.00853571
R24257 VSS.n6296 VSS.n6290 0.00853571
R24258 VSS.n6376 VSS.n6290 0.00853571
R24259 VSS.n6347 VSS.n6345 0.00853571
R24260 VSS.n6347 VSS.n6346 0.00853571
R24261 VSS.n6352 VSS.n6332 0.00853571
R24262 VSS.n5975 VSS.n5963 0.00853571
R24263 VSS.n5981 VSS.n5964 0.00853571
R24264 VSS.n5946 VSS.n5944 0.00853571
R24265 VSS.n7785 VSS.n7784 0.00853571
R24266 VSS.n7808 VSS.n7747 0.00853571
R24267 VSS.n7960 VSS.n7630 0.00853571
R24268 VSS.n7962 VSS.n7961 0.00853571
R24269 VSS.n7998 VSS.n7621 0.00853571
R24270 VSS.n8038 VSS.n8037 0.00853571
R24271 VSS.n8077 VSS.n7586 0.00853571
R24272 VSS.n8090 VSS.n8089 0.00853571
R24273 VSS.n8002 VSS.n7619 0.00853571
R24274 VSS.n8009 VSS.n7616 0.00853571
R24275 VSS.n8039 VSS.n7594 0.00853571
R24276 VSS.n8044 VSS.n8043 0.00853571
R24277 VSS.n8091 VSS.n7576 0.00853571
R24278 VSS.n8091 VSS.n7577 0.00853571
R24279 VSS.n8114 VSS.n7563 0.00853571
R24280 VSS.n8115 VSS.n8114 0.00853571
R24281 VSS.n8137 VSS.n7550 0.00853571
R24282 VSS.n7777 VSS.n7765 0.00853571
R24283 VSS.n7783 VSS.n7766 0.00853571
R24284 VSS.n7748 VSS.n7746 0.00853571
R24285 VSS.n8377 VSS.n8376 0.00853571
R24286 VSS.n8400 VSS.n8339 0.00853571
R24287 VSS.n8552 VSS.n8222 0.00853571
R24288 VSS.n8554 VSS.n8553 0.00853571
R24289 VSS.n8590 VSS.n8213 0.00853571
R24290 VSS.n8630 VSS.n8629 0.00853571
R24291 VSS.n8669 VSS.n8178 0.00853571
R24292 VSS.n8682 VSS.n8681 0.00853571
R24293 VSS.n8594 VSS.n8211 0.00853571
R24294 VSS.n8601 VSS.n8208 0.00853571
R24295 VSS.n8631 VSS.n8186 0.00853571
R24296 VSS.n8636 VSS.n8635 0.00853571
R24297 VSS.n8683 VSS.n8168 0.00853571
R24298 VSS.n8683 VSS.n8169 0.00853571
R24299 VSS.n8706 VSS.n8155 0.00853571
R24300 VSS.n8707 VSS.n8706 0.00853571
R24301 VSS.n8729 VSS.n8142 0.00853571
R24302 VSS.n8369 VSS.n8357 0.00853571
R24303 VSS.n8375 VSS.n8358 0.00853571
R24304 VSS.n8340 VSS.n8338 0.00853571
R24305 VSS.n8969 VSS.n8968 0.00853571
R24306 VSS.n8992 VSS.n8931 0.00853571
R24307 VSS.n9144 VSS.n8814 0.00853571
R24308 VSS.n9146 VSS.n9145 0.00853571
R24309 VSS.n9182 VSS.n8805 0.00853571
R24310 VSS.n9222 VSS.n9221 0.00853571
R24311 VSS.n9261 VSS.n8770 0.00853571
R24312 VSS.n9274 VSS.n9273 0.00853571
R24313 VSS.n9186 VSS.n8803 0.00853571
R24314 VSS.n9193 VSS.n8800 0.00853571
R24315 VSS.n9223 VSS.n8778 0.00853571
R24316 VSS.n9228 VSS.n9227 0.00853571
R24317 VSS.n9275 VSS.n8760 0.00853571
R24318 VSS.n9275 VSS.n8761 0.00853571
R24319 VSS.n9298 VSS.n8747 0.00853571
R24320 VSS.n9299 VSS.n9298 0.00853571
R24321 VSS.n9321 VSS.n8734 0.00853571
R24322 VSS.n8961 VSS.n8949 0.00853571
R24323 VSS.n8967 VSS.n8950 0.00853571
R24324 VSS.n8932 VSS.n8930 0.00853571
R24325 VSS.n10153 VSS.n10152 0.00853571
R24326 VSS.n10176 VSS.n10115 0.00853571
R24327 VSS.n10328 VSS.n9998 0.00853571
R24328 VSS.n10330 VSS.n10329 0.00853571
R24329 VSS.n10366 VSS.n9989 0.00853571
R24330 VSS.n10406 VSS.n10405 0.00853571
R24331 VSS.n10445 VSS.n9954 0.00853571
R24332 VSS.n10458 VSS.n10457 0.00853571
R24333 VSS.n10370 VSS.n9987 0.00853571
R24334 VSS.n10377 VSS.n9984 0.00853571
R24335 VSS.n10407 VSS.n9962 0.00853571
R24336 VSS.n10412 VSS.n10411 0.00853571
R24337 VSS.n10459 VSS.n9944 0.00853571
R24338 VSS.n10459 VSS.n9945 0.00853571
R24339 VSS.n10482 VSS.n9931 0.00853571
R24340 VSS.n10483 VSS.n10482 0.00853571
R24341 VSS.n10505 VSS.n9918 0.00853571
R24342 VSS.n10145 VSS.n10133 0.00853571
R24343 VSS.n10151 VSS.n10134 0.00853571
R24344 VSS.n10116 VSS.n10114 0.00853571
R24345 VSS.n10745 VSS.n10744 0.00853571
R24346 VSS.n10768 VSS.n10707 0.00853571
R24347 VSS.n10920 VSS.n10590 0.00853571
R24348 VSS.n10922 VSS.n10921 0.00853571
R24349 VSS.n10958 VSS.n10581 0.00853571
R24350 VSS.n10998 VSS.n10997 0.00853571
R24351 VSS.n11037 VSS.n10546 0.00853571
R24352 VSS.n11050 VSS.n11049 0.00853571
R24353 VSS.n10962 VSS.n10579 0.00853571
R24354 VSS.n10969 VSS.n10576 0.00853571
R24355 VSS.n10999 VSS.n10554 0.00853571
R24356 VSS.n11004 VSS.n11003 0.00853571
R24357 VSS.n11051 VSS.n10536 0.00853571
R24358 VSS.n11051 VSS.n10537 0.00853571
R24359 VSS.n11074 VSS.n10523 0.00853571
R24360 VSS.n11075 VSS.n11074 0.00853571
R24361 VSS.n11097 VSS.n10510 0.00853571
R24362 VSS.n10737 VSS.n10725 0.00853571
R24363 VSS.n10743 VSS.n10726 0.00853571
R24364 VSS.n10708 VSS.n10706 0.00853571
R24365 VSS.n11337 VSS.n11336 0.00853571
R24366 VSS.n11360 VSS.n11299 0.00853571
R24367 VSS.n11512 VSS.n11182 0.00853571
R24368 VSS.n11514 VSS.n11513 0.00853571
R24369 VSS.n11550 VSS.n11173 0.00853571
R24370 VSS.n11590 VSS.n11589 0.00853571
R24371 VSS.n11629 VSS.n11138 0.00853571
R24372 VSS.n11642 VSS.n11641 0.00853571
R24373 VSS.n11554 VSS.n11171 0.00853571
R24374 VSS.n11561 VSS.n11168 0.00853571
R24375 VSS.n11591 VSS.n11146 0.00853571
R24376 VSS.n11596 VSS.n11595 0.00853571
R24377 VSS.n11643 VSS.n11128 0.00853571
R24378 VSS.n11643 VSS.n11129 0.00853571
R24379 VSS.n11666 VSS.n11115 0.00853571
R24380 VSS.n11667 VSS.n11666 0.00853571
R24381 VSS.n11689 VSS.n11102 0.00853571
R24382 VSS.n11329 VSS.n11317 0.00853571
R24383 VSS.n11335 VSS.n11318 0.00853571
R24384 VSS.n11300 VSS.n11298 0.00853571
R24385 VSS.n11929 VSS.n11928 0.00853571
R24386 VSS.n11952 VSS.n11891 0.00853571
R24387 VSS.n12104 VSS.n11774 0.00853571
R24388 VSS.n12106 VSS.n12105 0.00853571
R24389 VSS.n12142 VSS.n11765 0.00853571
R24390 VSS.n12182 VSS.n12181 0.00853571
R24391 VSS.n12221 VSS.n11730 0.00853571
R24392 VSS.n12234 VSS.n12233 0.00853571
R24393 VSS.n12146 VSS.n11763 0.00853571
R24394 VSS.n12153 VSS.n11760 0.00853571
R24395 VSS.n12183 VSS.n11738 0.00853571
R24396 VSS.n12188 VSS.n12187 0.00853571
R24397 VSS.n12235 VSS.n11720 0.00853571
R24398 VSS.n12235 VSS.n11721 0.00853571
R24399 VSS.n12258 VSS.n11707 0.00853571
R24400 VSS.n12259 VSS.n12258 0.00853571
R24401 VSS.n12281 VSS.n11694 0.00853571
R24402 VSS.n11921 VSS.n11909 0.00853571
R24403 VSS.n11927 VSS.n11910 0.00853571
R24404 VSS.n11892 VSS.n11890 0.00853571
R24405 VSS.n12521 VSS.n12520 0.00853571
R24406 VSS.n12544 VSS.n12483 0.00853571
R24407 VSS.n12696 VSS.n12366 0.00853571
R24408 VSS.n12698 VSS.n12697 0.00853571
R24409 VSS.n12734 VSS.n12357 0.00853571
R24410 VSS.n12774 VSS.n12773 0.00853571
R24411 VSS.n12813 VSS.n12322 0.00853571
R24412 VSS.n12826 VSS.n12825 0.00853571
R24413 VSS.n12738 VSS.n12355 0.00853571
R24414 VSS.n12745 VSS.n12352 0.00853571
R24415 VSS.n12775 VSS.n12330 0.00853571
R24416 VSS.n12780 VSS.n12779 0.00853571
R24417 VSS.n12827 VSS.n12312 0.00853571
R24418 VSS.n12827 VSS.n12313 0.00853571
R24419 VSS.n12850 VSS.n12299 0.00853571
R24420 VSS.n12851 VSS.n12850 0.00853571
R24421 VSS.n12873 VSS.n12286 0.00853571
R24422 VSS.n12513 VSS.n12501 0.00853571
R24423 VSS.n12519 VSS.n12502 0.00853571
R24424 VSS.n12484 VSS.n12482 0.00853571
R24425 VSS.n13113 VSS.n13112 0.00853571
R24426 VSS.n13136 VSS.n13075 0.00853571
R24427 VSS.n13288 VSS.n12958 0.00853571
R24428 VSS.n13290 VSS.n13289 0.00853571
R24429 VSS.n13326 VSS.n12949 0.00853571
R24430 VSS.n13366 VSS.n13365 0.00853571
R24431 VSS.n13405 VSS.n12914 0.00853571
R24432 VSS.n13418 VSS.n13417 0.00853571
R24433 VSS.n13330 VSS.n12947 0.00853571
R24434 VSS.n13337 VSS.n12944 0.00853571
R24435 VSS.n13367 VSS.n12922 0.00853571
R24436 VSS.n13372 VSS.n13371 0.00853571
R24437 VSS.n13419 VSS.n12904 0.00853571
R24438 VSS.n13419 VSS.n12905 0.00853571
R24439 VSS.n13442 VSS.n12891 0.00853571
R24440 VSS.n13443 VSS.n13442 0.00853571
R24441 VSS.n13465 VSS.n12878 0.00853571
R24442 VSS.n13105 VSS.n13093 0.00853571
R24443 VSS.n13111 VSS.n13094 0.00853571
R24444 VSS.n13076 VSS.n13074 0.00853571
R24445 VSS.n13705 VSS.n13704 0.00853571
R24446 VSS.n13728 VSS.n13667 0.00853571
R24447 VSS.n13880 VSS.n13550 0.00853571
R24448 VSS.n13882 VSS.n13881 0.00853571
R24449 VSS.n13918 VSS.n13541 0.00853571
R24450 VSS.n13958 VSS.n13957 0.00853571
R24451 VSS.n13997 VSS.n13506 0.00853571
R24452 VSS.n14010 VSS.n14009 0.00853571
R24453 VSS.n13922 VSS.n13539 0.00853571
R24454 VSS.n13929 VSS.n13536 0.00853571
R24455 VSS.n13959 VSS.n13514 0.00853571
R24456 VSS.n13964 VSS.n13963 0.00853571
R24457 VSS.n14011 VSS.n13496 0.00853571
R24458 VSS.n14011 VSS.n13497 0.00853571
R24459 VSS.n14034 VSS.n13483 0.00853571
R24460 VSS.n14035 VSS.n14034 0.00853571
R24461 VSS.n14057 VSS.n13470 0.00853571
R24462 VSS.n13697 VSS.n13685 0.00853571
R24463 VSS.n13703 VSS.n13686 0.00853571
R24464 VSS.n13668 VSS.n13666 0.00853571
R24465 VSS.n14297 VSS.n14296 0.00853571
R24466 VSS.n14320 VSS.n14259 0.00853571
R24467 VSS.n14472 VSS.n14142 0.00853571
R24468 VSS.n14474 VSS.n14473 0.00853571
R24469 VSS.n14510 VSS.n14133 0.00853571
R24470 VSS.n14550 VSS.n14549 0.00853571
R24471 VSS.n14589 VSS.n14098 0.00853571
R24472 VSS.n14602 VSS.n14601 0.00853571
R24473 VSS.n14514 VSS.n14131 0.00853571
R24474 VSS.n14521 VSS.n14128 0.00853571
R24475 VSS.n14551 VSS.n14106 0.00853571
R24476 VSS.n14556 VSS.n14555 0.00853571
R24477 VSS.n14603 VSS.n14088 0.00853571
R24478 VSS.n14603 VSS.n14089 0.00853571
R24479 VSS.n14626 VSS.n14075 0.00853571
R24480 VSS.n14627 VSS.n14626 0.00853571
R24481 VSS.n14649 VSS.n14062 0.00853571
R24482 VSS.n14289 VSS.n14277 0.00853571
R24483 VSS.n14295 VSS.n14278 0.00853571
R24484 VSS.n14260 VSS.n14258 0.00853571
R24485 VSS.n14889 VSS.n14888 0.00853571
R24486 VSS.n14912 VSS.n14851 0.00853571
R24487 VSS.n15064 VSS.n14734 0.00853571
R24488 VSS.n15066 VSS.n15065 0.00853571
R24489 VSS.n15102 VSS.n14725 0.00853571
R24490 VSS.n15142 VSS.n15141 0.00853571
R24491 VSS.n15181 VSS.n14690 0.00853571
R24492 VSS.n15194 VSS.n15193 0.00853571
R24493 VSS.n15106 VSS.n14723 0.00853571
R24494 VSS.n15113 VSS.n14720 0.00853571
R24495 VSS.n15143 VSS.n14698 0.00853571
R24496 VSS.n15148 VSS.n15147 0.00853571
R24497 VSS.n15195 VSS.n14680 0.00853571
R24498 VSS.n15195 VSS.n14681 0.00853571
R24499 VSS.n15218 VSS.n14667 0.00853571
R24500 VSS.n15219 VSS.n15218 0.00853571
R24501 VSS.n15241 VSS.n14654 0.00853571
R24502 VSS.n14881 VSS.n14869 0.00853571
R24503 VSS.n14887 VSS.n14870 0.00853571
R24504 VSS.n14852 VSS.n14850 0.00853571
R24505 VSS.n15481 VSS.n15480 0.00853571
R24506 VSS.n15504 VSS.n15443 0.00853571
R24507 VSS.n15656 VSS.n15326 0.00853571
R24508 VSS.n15658 VSS.n15657 0.00853571
R24509 VSS.n15694 VSS.n15317 0.00853571
R24510 VSS.n15734 VSS.n15733 0.00853571
R24511 VSS.n15773 VSS.n15282 0.00853571
R24512 VSS.n15786 VSS.n15785 0.00853571
R24513 VSS.n15698 VSS.n15315 0.00853571
R24514 VSS.n15705 VSS.n15312 0.00853571
R24515 VSS.n15735 VSS.n15290 0.00853571
R24516 VSS.n15740 VSS.n15739 0.00853571
R24517 VSS.n15787 VSS.n15272 0.00853571
R24518 VSS.n15787 VSS.n15273 0.00853571
R24519 VSS.n15810 VSS.n15259 0.00853571
R24520 VSS.n15811 VSS.n15810 0.00853571
R24521 VSS.n15833 VSS.n15246 0.00853571
R24522 VSS.n15473 VSS.n15461 0.00853571
R24523 VSS.n15479 VSS.n15462 0.00853571
R24524 VSS.n15444 VSS.n15442 0.00853571
R24525 VSS.n6589 VSS.n6588 0.00853571
R24526 VSS.n6612 VSS.n6551 0.00853571
R24527 VSS.n6721 VSS.n6712 0.00853571
R24528 VSS.n6797 VSS.n6710 0.00853571
R24529 VSS.n6714 VSS.n6711 0.00853571
R24530 VSS.n15889 VSS.n15888 0.00853571
R24531 VSS.n15877 VSS.n6864 0.00853571
R24532 VSS.n15865 VSS.n6892 0.00853571
R24533 VSS.n6830 VSS.n6826 0.00853571
R24534 VSS.n6835 VSS.n6820 0.00853571
R24535 VSS.n15890 VSS.n6847 0.00853571
R24536 VSS.n6874 VSS.n6873 0.00853571
R24537 VSS.n6902 VSS.n6896 0.00853571
R24538 VSS.n15864 VSS.n6896 0.00853571
R24539 VSS.n6953 VSS.n6951 0.00853571
R24540 VSS.n6953 VSS.n6952 0.00853571
R24541 VSS.n15840 VSS.n6938 0.00853571
R24542 VSS.n6581 VSS.n6569 0.00853571
R24543 VSS.n6587 VSS.n6570 0.00853571
R24544 VSS.n6552 VSS.n6550 0.00853571
R24545 VSS.n7186 VSS.n7185 0.00853571
R24546 VSS.n7204 VSS.n7203 0.00853571
R24547 VSS.n7368 VSS.n7037 0.00853571
R24548 VSS.n7370 VSS.n7369 0.00853571
R24549 VSS.n7406 VSS.n7028 0.00853571
R24550 VSS.n7446 VSS.n7445 0.00853571
R24551 VSS.n7485 VSS.n6993 0.00853571
R24552 VSS.n7498 VSS.n7497 0.00853571
R24553 VSS.n7410 VSS.n7026 0.00853571
R24554 VSS.n7417 VSS.n7023 0.00853571
R24555 VSS.n7447 VSS.n7001 0.00853571
R24556 VSS.n7452 VSS.n7451 0.00853571
R24557 VSS.n7499 VSS.n6983 0.00853571
R24558 VSS.n7499 VSS.n6984 0.00853571
R24559 VSS.n7522 VSS.n6970 0.00853571
R24560 VSS.n7523 VSS.n7522 0.00853571
R24561 VSS.n7545 VSS.n6957 0.00853571
R24562 VSS.n7178 VSS.n7167 0.00853571
R24563 VSS.n7184 VSS.n7168 0.00853571
R24564 VSS.n7213 VSS.n7151 0.00853571
R24565 VSS.n349 VSS.n348 0.00853571
R24566 VSS.n367 VSS.n366 0.00853571
R24567 VSS.n18680 VSS.n135 0.00853571
R24568 VSS.n18682 VSS.n18681 0.00853571
R24569 VSS.n18718 VSS.n126 0.00853571
R24570 VSS.n18758 VSS.n18757 0.00853571
R24571 VSS.n18797 VSS.n91 0.00853571
R24572 VSS.n18810 VSS.n18809 0.00853571
R24573 VSS.n18722 VSS.n124 0.00853571
R24574 VSS.n18729 VSS.n121 0.00853571
R24575 VSS.n18759 VSS.n99 0.00853571
R24576 VSS.n18764 VSS.n18763 0.00853571
R24577 VSS.n18811 VSS.n81 0.00853571
R24578 VSS.n18811 VSS.n82 0.00853571
R24579 VSS.n18834 VSS.n68 0.00853571
R24580 VSS.n18835 VSS.n18834 0.00853571
R24581 VSS.n18857 VSS.n55 0.00853571
R24582 VSS.n449 VSS.n448 0.00853571
R24583 VSS.n350 VSS.n347 0.00853571
R24584 VSS.n368 VSS.n301 0.00853571
R24585 VSS.n541 VSS.n532 0.00853571
R24586 VSS.n620 VSS.n530 0.00853571
R24587 VSS.n534 VSS.n531 0.00853571
R24588 VSS.n803 VSS.n802 0.00853571
R24589 VSS.n791 VSS.n687 0.00853571
R24590 VSS.n779 VSS.n715 0.00853571
R24591 VSS.n653 VSS.n649 0.00853571
R24592 VSS.n658 VSS.n643 0.00853571
R24593 VSS.n804 VSS.n670 0.00853571
R24594 VSS.n697 VSS.n696 0.00853571
R24595 VSS.n725 VSS.n719 0.00853571
R24596 VSS.n778 VSS.n719 0.00853571
R24597 VSS.n735 VSS.n734 0.00853571
R24598 VSS.n734 VSS.n732 0.00853571
R24599 VSS.n18863 VSS.n51 0.00853571
R24600 VSS.n1014 VSS.n1013 0.00853571
R24601 VSS.n911 VSS.n910 0.00853571
R24602 VSS.n921 VSS.n467 0.00853571
R24603 VSS.n17917 VSS.n17916 0.00853571
R24604 VSS.n17905 VSS.n1346 0.00853571
R24605 VSS.n17893 VSS.n1374 0.00853571
R24606 VSS.n1312 VSS.n1308 0.00853571
R24607 VSS.n1317 VSS.n1302 0.00853571
R24608 VSS.n17918 VSS.n1329 0.00853571
R24609 VSS.n1356 VSS.n1355 0.00853571
R24610 VSS.n1384 VSS.n1378 0.00853571
R24611 VSS.n17892 VSS.n1378 0.00853571
R24612 VSS.n1435 VSS.n1433 0.00853571
R24613 VSS.n1435 VSS.n1434 0.00853571
R24614 VSS.n17868 VSS.n1420 0.00853571
R24615 VSS.n18038 VSS.n1025 0.00822143
R24616 VSS.n18030 VSS.n1027 0.00822143
R24617 VSS.n18013 VSS.n1051 0.00822143
R24618 VSS.n17007 VSS.n1057 0.00822143
R24619 VSS.n17008 VSS.n16996 0.00822143
R24620 VSS.n17038 VSS.n16982 0.00822143
R24621 VSS.n17069 VSS.n16944 0.00822143
R24622 VSS.n17133 VSS.n16932 0.00822143
R24623 VSS.n17502 VSS.n17490 0.00822143
R24624 VSS.n17537 VSS.n17470 0.00822143
R24625 VSS.n17570 VSS.n17439 0.00822143
R24626 VSS.n17599 VSS.n17421 0.00822143
R24627 VSS.n17600 VSS.n17410 0.00822143
R24628 VSS.n17630 VSS.n17396 0.00822143
R24629 VSS.n17661 VSS.n17358 0.00822143
R24630 VSS.n17725 VSS.n17346 0.00822143
R24631 VSS.n18079 VSS.n282 0.00822143
R24632 VSS.n18114 VSS.n262 0.00822143
R24633 VSS.n18147 VSS.n231 0.00822143
R24634 VSS.n18176 VSS.n213 0.00822143
R24635 VSS.n18578 VSS.n18177 0.00822143
R24636 VSS.n18570 VSS.n18179 0.00822143
R24637 VSS.n18553 VSS.n18202 0.00822143
R24638 VSS.n18327 VSS.n18208 0.00822143
R24639 VSS.n9650 VSS.n9460 0.00822143
R24640 VSS.n9680 VSS.n9446 0.00822143
R24641 VSS.n9711 VSS.n9408 0.00822143
R24642 VSS.n9775 VSS.n9396 0.00822143
R24643 VSS.n16488 VSS.n16477 0.00822143
R24644 VSS.n16518 VSS.n16465 0.00822143
R24645 VSS.n16549 VSS.n16425 0.00822143
R24646 VSS.n16592 VSS.n16413 0.00822143
R24647 VSS.n16593 VSS.n16402 0.00822143
R24648 VSS.n16623 VSS.n16388 0.00822143
R24649 VSS.n16654 VSS.n16350 0.00822143
R24650 VSS.n16718 VSS.n16338 0.00822143
R24651 VSS.n1653 VSS.n1642 0.00822143
R24652 VSS.n1683 VSS.n1630 0.00822143
R24653 VSS.n1714 VSS.n1590 0.00822143
R24654 VSS.n15999 VSS.n1578 0.00822143
R24655 VSS.n16000 VSS.n1574 0.00822143
R24656 VSS.n16030 VSS.n1560 0.00822143
R24657 VSS.n16061 VSS.n1522 0.00822143
R24658 VSS.n16125 VSS.n1510 0.00822143
R24659 VSS.n1844 VSS.n1832 0.00822143
R24660 VSS.n1879 VSS.n1812 0.00822143
R24661 VSS.n1912 VSS.n1781 0.00822143
R24662 VSS.n1941 VSS.n1763 0.00822143
R24663 VSS.n2343 VSS.n1942 0.00822143
R24664 VSS.n2335 VSS.n1944 0.00822143
R24665 VSS.n2318 VSS.n1967 0.00822143
R24666 VSS.n2091 VSS.n1973 0.00822143
R24667 VSS.n3043 VSS.n3031 0.00822143
R24668 VSS.n3078 VSS.n3011 0.00822143
R24669 VSS.n3111 VSS.n2980 0.00822143
R24670 VSS.n3140 VSS.n2962 0.00822143
R24671 VSS.n3141 VSS.n2951 0.00822143
R24672 VSS.n3171 VSS.n2937 0.00822143
R24673 VSS.n3202 VSS.n2899 0.00822143
R24674 VSS.n3266 VSS.n2887 0.00822143
R24675 VSS.n3635 VSS.n3623 0.00822143
R24676 VSS.n3670 VSS.n3603 0.00822143
R24677 VSS.n3703 VSS.n3572 0.00822143
R24678 VSS.n3732 VSS.n3554 0.00822143
R24679 VSS.n3733 VSS.n3543 0.00822143
R24680 VSS.n3763 VSS.n3529 0.00822143
R24681 VSS.n3794 VSS.n3491 0.00822143
R24682 VSS.n3858 VSS.n3479 0.00822143
R24683 VSS.n4227 VSS.n4215 0.00822143
R24684 VSS.n4262 VSS.n4195 0.00822143
R24685 VSS.n4295 VSS.n4164 0.00822143
R24686 VSS.n4324 VSS.n4146 0.00822143
R24687 VSS.n4325 VSS.n4135 0.00822143
R24688 VSS.n4355 VSS.n4121 0.00822143
R24689 VSS.n4386 VSS.n4083 0.00822143
R24690 VSS.n4450 VSS.n4071 0.00822143
R24691 VSS.n4819 VSS.n4807 0.00822143
R24692 VSS.n4854 VSS.n4787 0.00822143
R24693 VSS.n4887 VSS.n4756 0.00822143
R24694 VSS.n4916 VSS.n4738 0.00822143
R24695 VSS.n4917 VSS.n4727 0.00822143
R24696 VSS.n4947 VSS.n4713 0.00822143
R24697 VSS.n4978 VSS.n4675 0.00822143
R24698 VSS.n5042 VSS.n4663 0.00822143
R24699 VSS.n2440 VSS.n2428 0.00822143
R24700 VSS.n2475 VSS.n2408 0.00822143
R24701 VSS.n2508 VSS.n2377 0.00822143
R24702 VSS.n2537 VSS.n2359 0.00822143
R24703 VSS.n5308 VSS.n2538 0.00822143
R24704 VSS.n5300 VSS.n2540 0.00822143
R24705 VSS.n5283 VSS.n2563 0.00822143
R24706 VSS.n2687 VSS.n2569 0.00822143
R24707 VSS.n5401 VSS.n5389 0.00822143
R24708 VSS.n5436 VSS.n5369 0.00822143
R24709 VSS.n5469 VSS.n5338 0.00822143
R24710 VSS.n5498 VSS.n5320 0.00822143
R24711 VSS.n5881 VSS.n5499 0.00822143
R24712 VSS.n5873 VSS.n5501 0.00822143
R24713 VSS.n5856 VSS.n5524 0.00822143
R24714 VSS.n5648 VSS.n5530 0.00822143
R24715 VSS.n5974 VSS.n5962 0.00822143
R24716 VSS.n6009 VSS.n5942 0.00822143
R24717 VSS.n6042 VSS.n5911 0.00822143
R24718 VSS.n6071 VSS.n5893 0.00822143
R24719 VSS.n6473 VSS.n6072 0.00822143
R24720 VSS.n6465 VSS.n6074 0.00822143
R24721 VSS.n6448 VSS.n6097 0.00822143
R24722 VSS.n6221 VSS.n6103 0.00822143
R24723 VSS.n7776 VSS.n7764 0.00822143
R24724 VSS.n7811 VSS.n7744 0.00822143
R24725 VSS.n7844 VSS.n7713 0.00822143
R24726 VSS.n7873 VSS.n7695 0.00822143
R24727 VSS.n7874 VSS.n7684 0.00822143
R24728 VSS.n7904 VSS.n7670 0.00822143
R24729 VSS.n7935 VSS.n7632 0.00822143
R24730 VSS.n7999 VSS.n7620 0.00822143
R24731 VSS.n8368 VSS.n8356 0.00822143
R24732 VSS.n8403 VSS.n8336 0.00822143
R24733 VSS.n8436 VSS.n8305 0.00822143
R24734 VSS.n8465 VSS.n8287 0.00822143
R24735 VSS.n8466 VSS.n8276 0.00822143
R24736 VSS.n8496 VSS.n8262 0.00822143
R24737 VSS.n8527 VSS.n8224 0.00822143
R24738 VSS.n8591 VSS.n8212 0.00822143
R24739 VSS.n8960 VSS.n8948 0.00822143
R24740 VSS.n8995 VSS.n8928 0.00822143
R24741 VSS.n9028 VSS.n8897 0.00822143
R24742 VSS.n9057 VSS.n8879 0.00822143
R24743 VSS.n9058 VSS.n8868 0.00822143
R24744 VSS.n9088 VSS.n8854 0.00822143
R24745 VSS.n9119 VSS.n8816 0.00822143
R24746 VSS.n9183 VSS.n8804 0.00822143
R24747 VSS.n10144 VSS.n10132 0.00822143
R24748 VSS.n10179 VSS.n10112 0.00822143
R24749 VSS.n10212 VSS.n10081 0.00822143
R24750 VSS.n10241 VSS.n10063 0.00822143
R24751 VSS.n10242 VSS.n10052 0.00822143
R24752 VSS.n10272 VSS.n10038 0.00822143
R24753 VSS.n10303 VSS.n10000 0.00822143
R24754 VSS.n10367 VSS.n9988 0.00822143
R24755 VSS.n10736 VSS.n10724 0.00822143
R24756 VSS.n10771 VSS.n10704 0.00822143
R24757 VSS.n10804 VSS.n10673 0.00822143
R24758 VSS.n10833 VSS.n10655 0.00822143
R24759 VSS.n10834 VSS.n10644 0.00822143
R24760 VSS.n10864 VSS.n10630 0.00822143
R24761 VSS.n10895 VSS.n10592 0.00822143
R24762 VSS.n10959 VSS.n10580 0.00822143
R24763 VSS.n11328 VSS.n11316 0.00822143
R24764 VSS.n11363 VSS.n11296 0.00822143
R24765 VSS.n11396 VSS.n11265 0.00822143
R24766 VSS.n11425 VSS.n11247 0.00822143
R24767 VSS.n11426 VSS.n11236 0.00822143
R24768 VSS.n11456 VSS.n11222 0.00822143
R24769 VSS.n11487 VSS.n11184 0.00822143
R24770 VSS.n11551 VSS.n11172 0.00822143
R24771 VSS.n11920 VSS.n11908 0.00822143
R24772 VSS.n11955 VSS.n11888 0.00822143
R24773 VSS.n11988 VSS.n11857 0.00822143
R24774 VSS.n12017 VSS.n11839 0.00822143
R24775 VSS.n12018 VSS.n11828 0.00822143
R24776 VSS.n12048 VSS.n11814 0.00822143
R24777 VSS.n12079 VSS.n11776 0.00822143
R24778 VSS.n12143 VSS.n11764 0.00822143
R24779 VSS.n12512 VSS.n12500 0.00822143
R24780 VSS.n12547 VSS.n12480 0.00822143
R24781 VSS.n12580 VSS.n12449 0.00822143
R24782 VSS.n12609 VSS.n12431 0.00822143
R24783 VSS.n12610 VSS.n12420 0.00822143
R24784 VSS.n12640 VSS.n12406 0.00822143
R24785 VSS.n12671 VSS.n12368 0.00822143
R24786 VSS.n12735 VSS.n12356 0.00822143
R24787 VSS.n13104 VSS.n13092 0.00822143
R24788 VSS.n13139 VSS.n13072 0.00822143
R24789 VSS.n13172 VSS.n13041 0.00822143
R24790 VSS.n13201 VSS.n13023 0.00822143
R24791 VSS.n13202 VSS.n13012 0.00822143
R24792 VSS.n13232 VSS.n12998 0.00822143
R24793 VSS.n13263 VSS.n12960 0.00822143
R24794 VSS.n13327 VSS.n12948 0.00822143
R24795 VSS.n13696 VSS.n13684 0.00822143
R24796 VSS.n13731 VSS.n13664 0.00822143
R24797 VSS.n13764 VSS.n13633 0.00822143
R24798 VSS.n13793 VSS.n13615 0.00822143
R24799 VSS.n13794 VSS.n13604 0.00822143
R24800 VSS.n13824 VSS.n13590 0.00822143
R24801 VSS.n13855 VSS.n13552 0.00822143
R24802 VSS.n13919 VSS.n13540 0.00822143
R24803 VSS.n14288 VSS.n14276 0.00822143
R24804 VSS.n14323 VSS.n14256 0.00822143
R24805 VSS.n14356 VSS.n14225 0.00822143
R24806 VSS.n14385 VSS.n14207 0.00822143
R24807 VSS.n14386 VSS.n14196 0.00822143
R24808 VSS.n14416 VSS.n14182 0.00822143
R24809 VSS.n14447 VSS.n14144 0.00822143
R24810 VSS.n14511 VSS.n14132 0.00822143
R24811 VSS.n14880 VSS.n14868 0.00822143
R24812 VSS.n14915 VSS.n14848 0.00822143
R24813 VSS.n14948 VSS.n14817 0.00822143
R24814 VSS.n14977 VSS.n14799 0.00822143
R24815 VSS.n14978 VSS.n14788 0.00822143
R24816 VSS.n15008 VSS.n14774 0.00822143
R24817 VSS.n15039 VSS.n14736 0.00822143
R24818 VSS.n15103 VSS.n14724 0.00822143
R24819 VSS.n15472 VSS.n15460 0.00822143
R24820 VSS.n15507 VSS.n15440 0.00822143
R24821 VSS.n15540 VSS.n15409 0.00822143
R24822 VSS.n15569 VSS.n15391 0.00822143
R24823 VSS.n15570 VSS.n15380 0.00822143
R24824 VSS.n15600 VSS.n15366 0.00822143
R24825 VSS.n15631 VSS.n15328 0.00822143
R24826 VSS.n15695 VSS.n15316 0.00822143
R24827 VSS.n6580 VSS.n6568 0.00822143
R24828 VSS.n6615 VSS.n6548 0.00822143
R24829 VSS.n6648 VSS.n6517 0.00822143
R24830 VSS.n6677 VSS.n6499 0.00822143
R24831 VSS.n15961 VSS.n6678 0.00822143
R24832 VSS.n15953 VSS.n6680 0.00822143
R24833 VSS.n15936 VSS.n6703 0.00822143
R24834 VSS.n6827 VSS.n6709 0.00822143
R24835 VSS.n7177 VSS.n7166 0.00822143
R24836 VSS.n7207 VSS.n7154 0.00822143
R24837 VSS.n7238 VSS.n7114 0.00822143
R24838 VSS.n7281 VSS.n7102 0.00822143
R24839 VSS.n7282 VSS.n7091 0.00822143
R24840 VSS.n7312 VSS.n7077 0.00822143
R24841 VSS.n7343 VSS.n7039 0.00822143
R24842 VSS.n7407 VSS.n7027 0.00822143
R24843 VSS.n447 VSS.n292 0.00822143
R24844 VSS.n439 VSS.n294 0.00822143
R24845 VSS.n422 VSS.n318 0.00822143
R24846 VSS.n18593 VSS.n193 0.00822143
R24847 VSS.n18594 VSS.n189 0.00822143
R24848 VSS.n18624 VSS.n175 0.00822143
R24849 VSS.n18655 VSS.n137 0.00822143
R24850 VSS.n18719 VSS.n125 0.00822143
R24851 VSS.n1012 VSS.n458 0.00822143
R24852 VSS.n1004 VSS.n460 0.00822143
R24853 VSS.n987 VSS.n484 0.00822143
R24854 VSS.n880 VSS.n490 0.00822143
R24855 VSS.n879 VSS.n495 0.00822143
R24856 VSS.n867 VSS.n500 0.00822143
R24857 VSS.n850 VSS.n523 0.00822143
R24858 VSS.n650 VSS.n529 0.00822143
R24859 VSS.n17989 VSS.n1160 0.00822143
R24860 VSS.n17981 VSS.n1162 0.00822143
R24861 VSS.n17964 VSS.n1185 0.00822143
R24862 VSS.n1309 VSS.n1191 0.00822143
R24863 VSS.n9552 VSS.n9540 0.00816667
R24864 VSS.n9587 VSS.n9520 0.00816667
R24865 VSS.n9620 VSS.n9489 0.00816667
R24866 VSS.n9649 VSS.n9471 0.00816667
R24867 VSS.n1240 VSS.n1239 0.00764286
R24868 VSS.n1263 VSS.n1262 0.00764286
R24869 VSS.n17991 VSS.n17990 0.00764286
R24870 VSS.n17982 VSS.n1167 0.00764286
R24871 VSS.n1237 VSS.n1169 0.00764286
R24872 VSS.n1174 VSS.n1173 0.00764286
R24873 VSS.n1182 VSS.n1181 0.00764286
R24874 VSS.n1265 VSS.n1183 0.00764286
R24875 VSS.n950 VSS.n947 0.00764286
R24876 VSS.n17034 VSS.n16986 0.00764286
R24877 VSS.n17072 VSS.n16958 0.00764286
R24878 VSS.n1131 VSS.n1128 0.00764286
R24879 VSS.n1039 VSS.n1038 0.00764286
R24880 VSS.n1048 VSS.n1047 0.00764286
R24881 VSS.n1130 VSS.n1129 0.00764286
R24882 VSS.n18012 VSS.n1052 0.00764286
R24883 VSS.n1062 VSS.n1059 0.00764286
R24884 VSS.n17142 VSS.n17141 0.00764286
R24885 VSS.n17140 VSS.n16923 0.00764286
R24886 VSS.n17172 VSS.n16909 0.00764286
R24887 VSS.n17224 VSS.n16890 0.00764286
R24888 VSS.n17256 VSS.n17255 0.00764286
R24889 VSS.n17255 VSS.n16873 0.00764286
R24890 VSS.n17137 VSS.n17136 0.00764286
R24891 VSS.n17137 VSS.n16928 0.00764286
R24892 VSS.n17143 VSS.n16929 0.00764286
R24893 VSS.n17139 VSS.n16925 0.00764286
R24894 VSS.n17158 VSS.n17157 0.00764286
R24895 VSS.n17173 VSS.n16908 0.00764286
R24896 VSS.n17195 VSS.n17194 0.00764286
R24897 VSS.n17231 VSS.n16886 0.00764286
R24898 VSS.n17254 VSS.n16872 0.00764286
R24899 VSS.n17254 VSS.n17253 0.00764286
R24900 VSS.n17009 VSS.n16997 0.00764286
R24901 VSS.n17037 VSS.n17036 0.00764286
R24902 VSS.n17044 VSS.n16979 0.00764286
R24903 VSS.n17040 VSS.n17039 0.00764286
R24904 VSS.n17062 VSS.n16965 0.00764286
R24905 VSS.n17076 VSS.n16959 0.00764286
R24906 VSS.n17626 VSS.n17400 0.00764286
R24907 VSS.n17664 VSS.n17372 0.00764286
R24908 VSS.n17453 VSS.n17447 0.00764286
R24909 VSS.n17540 VSS.n17467 0.00764286
R24910 VSS.n17548 VSS.n17547 0.00764286
R24911 VSS.n17452 VSS.n17451 0.00764286
R24912 VSS.n17571 VSS.n17442 0.00764286
R24913 VSS.n17598 VSS.n17422 0.00764286
R24914 VSS.n17734 VSS.n17733 0.00764286
R24915 VSS.n17732 VSS.n17337 0.00764286
R24916 VSS.n17764 VSS.n17323 0.00764286
R24917 VSS.n17816 VSS.n17304 0.00764286
R24918 VSS.n17848 VSS.n17847 0.00764286
R24919 VSS.n17847 VSS.n17287 0.00764286
R24920 VSS.n17729 VSS.n17728 0.00764286
R24921 VSS.n17729 VSS.n17342 0.00764286
R24922 VSS.n17735 VSS.n17343 0.00764286
R24923 VSS.n17731 VSS.n17339 0.00764286
R24924 VSS.n17750 VSS.n17749 0.00764286
R24925 VSS.n17765 VSS.n17322 0.00764286
R24926 VSS.n17787 VSS.n17786 0.00764286
R24927 VSS.n17823 VSS.n17300 0.00764286
R24928 VSS.n17846 VSS.n17286 0.00764286
R24929 VSS.n17846 VSS.n17845 0.00764286
R24930 VSS.n17601 VSS.n17411 0.00764286
R24931 VSS.n17629 VSS.n17628 0.00764286
R24932 VSS.n17636 VSS.n17393 0.00764286
R24933 VSS.n17632 VSS.n17631 0.00764286
R24934 VSS.n17654 VSS.n17379 0.00764286
R24935 VSS.n17668 VSS.n17373 0.00764286
R24936 VSS.n245 VSS.n239 0.00764286
R24937 VSS.n18257 VSS.n18256 0.00764286
R24938 VSS.n18280 VSS.n18279 0.00764286
R24939 VSS.n18580 VSS.n18579 0.00764286
R24940 VSS.n18571 VSS.n18184 0.00764286
R24941 VSS.n18254 VSS.n18186 0.00764286
R24942 VSS.n18191 VSS.n18190 0.00764286
R24943 VSS.n18199 VSS.n18198 0.00764286
R24944 VSS.n18282 VSS.n18200 0.00764286
R24945 VSS.n18334 VSS.n18333 0.00764286
R24946 VSS.n18526 VSS.n18314 0.00764286
R24947 VSS.n18512 VSS.n18342 0.00764286
R24948 VSS.n18489 VSS.n18488 0.00764286
R24949 VSS.n18474 VSS.n18423 0.00764286
R24950 VSS.n18474 VSS.n18473 0.00764286
R24951 VSS.n18331 VSS.n18330 0.00764286
R24952 VSS.n18331 VSS.n18319 0.00764286
R24953 VSS.n18335 VSS.n18321 0.00764286
R24954 VSS.n18320 VSS.n18315 0.00764286
R24955 VSS.n18515 VSS.n18514 0.00764286
R24956 VSS.n18348 VSS.n18341 0.00764286
R24957 VSS.n18412 VSS.n18411 0.00764286
R24958 VSS.n18445 VSS.n18444 0.00764286
R24959 VSS.n18476 VSS.n18475 0.00764286
R24960 VSS.n18475 VSS.n18425 0.00764286
R24961 VSS.n18117 VSS.n259 0.00764286
R24962 VSS.n18125 VSS.n18124 0.00764286
R24963 VSS.n244 VSS.n243 0.00764286
R24964 VSS.n18148 VSS.n234 0.00764286
R24965 VSS.n18175 VSS.n214 0.00764286
R24966 VSS.n9503 VSS.n9497 0.00764286
R24967 VSS.n9676 VSS.n9450 0.00764286
R24968 VSS.n9714 VSS.n9422 0.00764286
R24969 VSS.n9651 VSS.n9461 0.00764286
R24970 VSS.n9679 VSS.n9678 0.00764286
R24971 VSS.n9686 VSS.n9443 0.00764286
R24972 VSS.n9682 VSS.n9681 0.00764286
R24973 VSS.n9704 VSS.n9429 0.00764286
R24974 VSS.n9718 VSS.n9423 0.00764286
R24975 VSS.n9784 VSS.n9783 0.00764286
R24976 VSS.n9782 VSS.n9387 0.00764286
R24977 VSS.n9814 VSS.n9373 0.00764286
R24978 VSS.n9866 VSS.n9354 0.00764286
R24979 VSS.n9899 VSS.n9337 0.00764286
R24980 VSS.n9895 VSS.n9337 0.00764286
R24981 VSS.n9779 VSS.n9778 0.00764286
R24982 VSS.n9779 VSS.n9392 0.00764286
R24983 VSS.n9785 VSS.n9393 0.00764286
R24984 VSS.n9781 VSS.n9389 0.00764286
R24985 VSS.n9800 VSS.n9799 0.00764286
R24986 VSS.n9815 VSS.n9372 0.00764286
R24987 VSS.n9837 VSS.n9836 0.00764286
R24988 VSS.n9873 VSS.n9350 0.00764286
R24989 VSS.n9898 VSS.n9897 0.00764286
R24990 VSS.n9897 VSS.n9896 0.00764286
R24991 VSS.n9590 VSS.n9517 0.00764286
R24992 VSS.n9598 VSS.n9597 0.00764286
R24993 VSS.n9502 VSS.n9501 0.00764286
R24994 VSS.n9621 VSS.n9492 0.00764286
R24995 VSS.n9648 VSS.n9472 0.00764286
R24996 VSS.n16557 VSS.n16439 0.00764286
R24997 VSS.n16619 VSS.n16392 0.00764286
R24998 VSS.n16657 VSS.n16364 0.00764286
R24999 VSS.n16594 VSS.n16403 0.00764286
R25000 VSS.n16622 VSS.n16621 0.00764286
R25001 VSS.n16629 VSS.n16385 0.00764286
R25002 VSS.n16625 VSS.n16624 0.00764286
R25003 VSS.n16647 VSS.n16371 0.00764286
R25004 VSS.n16661 VSS.n16365 0.00764286
R25005 VSS.n16727 VSS.n16726 0.00764286
R25006 VSS.n16725 VSS.n16329 0.00764286
R25007 VSS.n16757 VSS.n16315 0.00764286
R25008 VSS.n16809 VSS.n16296 0.00764286
R25009 VSS.n16842 VSS.n16279 0.00764286
R25010 VSS.n16838 VSS.n16279 0.00764286
R25011 VSS.n16722 VSS.n16721 0.00764286
R25012 VSS.n16722 VSS.n16334 0.00764286
R25013 VSS.n16728 VSS.n16335 0.00764286
R25014 VSS.n16724 VSS.n16331 0.00764286
R25015 VSS.n16743 VSS.n16742 0.00764286
R25016 VSS.n16758 VSS.n16314 0.00764286
R25017 VSS.n16780 VSS.n16779 0.00764286
R25018 VSS.n16816 VSS.n16292 0.00764286
R25019 VSS.n16841 VSS.n16840 0.00764286
R25020 VSS.n16840 VSS.n16839 0.00764286
R25021 VSS.n16520 VSS.n16519 0.00764286
R25022 VSS.n16542 VSS.n16446 0.00764286
R25023 VSS.n16556 VSS.n16555 0.00764286
R25024 VSS.n16554 VSS.n16550 0.00764286
R25025 VSS.n16591 VSS.n16414 0.00764286
R25026 VSS.n1722 VSS.n1604 0.00764286
R25027 VSS.n16026 VSS.n1564 0.00764286
R25028 VSS.n16064 VSS.n1536 0.00764286
R25029 VSS.n16001 VSS.n1575 0.00764286
R25030 VSS.n16029 VSS.n16028 0.00764286
R25031 VSS.n16036 VSS.n1557 0.00764286
R25032 VSS.n16032 VSS.n16031 0.00764286
R25033 VSS.n16054 VSS.n1543 0.00764286
R25034 VSS.n16068 VSS.n1537 0.00764286
R25035 VSS.n16134 VSS.n16133 0.00764286
R25036 VSS.n16132 VSS.n1501 0.00764286
R25037 VSS.n16164 VSS.n1487 0.00764286
R25038 VSS.n16216 VSS.n1468 0.00764286
R25039 VSS.n16249 VSS.n1451 0.00764286
R25040 VSS.n16245 VSS.n1451 0.00764286
R25041 VSS.n16129 VSS.n16128 0.00764286
R25042 VSS.n16129 VSS.n1506 0.00764286
R25043 VSS.n16135 VSS.n1507 0.00764286
R25044 VSS.n16131 VSS.n1503 0.00764286
R25045 VSS.n16150 VSS.n16149 0.00764286
R25046 VSS.n16165 VSS.n1486 0.00764286
R25047 VSS.n16187 VSS.n16186 0.00764286
R25048 VSS.n16223 VSS.n1464 0.00764286
R25049 VSS.n16248 VSS.n16247 0.00764286
R25050 VSS.n16247 VSS.n16246 0.00764286
R25051 VSS.n1685 VSS.n1684 0.00764286
R25052 VSS.n1707 VSS.n1611 0.00764286
R25053 VSS.n1721 VSS.n1720 0.00764286
R25054 VSS.n1719 VSS.n1715 0.00764286
R25055 VSS.n15998 VSS.n1579 0.00764286
R25056 VSS.n1795 VSS.n1789 0.00764286
R25057 VSS.n2022 VSS.n2021 0.00764286
R25058 VSS.n2045 VSS.n2044 0.00764286
R25059 VSS.n2345 VSS.n2344 0.00764286
R25060 VSS.n2336 VSS.n1949 0.00764286
R25061 VSS.n2019 VSS.n1951 0.00764286
R25062 VSS.n1956 VSS.n1955 0.00764286
R25063 VSS.n1964 VSS.n1963 0.00764286
R25064 VSS.n2047 VSS.n1965 0.00764286
R25065 VSS.n2098 VSS.n2097 0.00764286
R25066 VSS.n2291 VSS.n2079 0.00764286
R25067 VSS.n2271 VSS.n2109 0.00764286
R25068 VSS.n2251 VSS.n2156 0.00764286
R25069 VSS.n2211 VSS.n2172 0.00764286
R25070 VSS.n2212 VSS.n2211 0.00764286
R25071 VSS.n2095 VSS.n2094 0.00764286
R25072 VSS.n2095 VSS.n2084 0.00764286
R25073 VSS.n2099 VSS.n2085 0.00764286
R25074 VSS.n2290 VSS.n2081 0.00764286
R25075 VSS.n2274 VSS.n2110 0.00764286
R25076 VSS.n2273 VSS.n2272 0.00764286
R25077 VSS.n2165 VSS.n2154 0.00764286
R25078 VSS.n2245 VSS.n2244 0.00764286
R25079 VSS.n2210 VSS.n2209 0.00764286
R25080 VSS.n2210 VSS.n2208 0.00764286
R25081 VSS.n1882 VSS.n1809 0.00764286
R25082 VSS.n1890 VSS.n1889 0.00764286
R25083 VSS.n1794 VSS.n1793 0.00764286
R25084 VSS.n1913 VSS.n1784 0.00764286
R25085 VSS.n1940 VSS.n1764 0.00764286
R25086 VSS.n2994 VSS.n2988 0.00764286
R25087 VSS.n3167 VSS.n2941 0.00764286
R25088 VSS.n3205 VSS.n2913 0.00764286
R25089 VSS.n3142 VSS.n2952 0.00764286
R25090 VSS.n3170 VSS.n3169 0.00764286
R25091 VSS.n3177 VSS.n2934 0.00764286
R25092 VSS.n3173 VSS.n3172 0.00764286
R25093 VSS.n3195 VSS.n2920 0.00764286
R25094 VSS.n3209 VSS.n2914 0.00764286
R25095 VSS.n3275 VSS.n3274 0.00764286
R25096 VSS.n3273 VSS.n2878 0.00764286
R25097 VSS.n3305 VSS.n2864 0.00764286
R25098 VSS.n3357 VSS.n2845 0.00764286
R25099 VSS.n3390 VSS.n2828 0.00764286
R25100 VSS.n3386 VSS.n2828 0.00764286
R25101 VSS.n3270 VSS.n3269 0.00764286
R25102 VSS.n3270 VSS.n2883 0.00764286
R25103 VSS.n3276 VSS.n2884 0.00764286
R25104 VSS.n3272 VSS.n2880 0.00764286
R25105 VSS.n3291 VSS.n3290 0.00764286
R25106 VSS.n3306 VSS.n2863 0.00764286
R25107 VSS.n3328 VSS.n3327 0.00764286
R25108 VSS.n3364 VSS.n2841 0.00764286
R25109 VSS.n3389 VSS.n3388 0.00764286
R25110 VSS.n3388 VSS.n3387 0.00764286
R25111 VSS.n3081 VSS.n3008 0.00764286
R25112 VSS.n3089 VSS.n3088 0.00764286
R25113 VSS.n2993 VSS.n2992 0.00764286
R25114 VSS.n3112 VSS.n2983 0.00764286
R25115 VSS.n3139 VSS.n2963 0.00764286
R25116 VSS.n3586 VSS.n3580 0.00764286
R25117 VSS.n3759 VSS.n3533 0.00764286
R25118 VSS.n3797 VSS.n3505 0.00764286
R25119 VSS.n3734 VSS.n3544 0.00764286
R25120 VSS.n3762 VSS.n3761 0.00764286
R25121 VSS.n3769 VSS.n3526 0.00764286
R25122 VSS.n3765 VSS.n3764 0.00764286
R25123 VSS.n3787 VSS.n3512 0.00764286
R25124 VSS.n3801 VSS.n3506 0.00764286
R25125 VSS.n3867 VSS.n3866 0.00764286
R25126 VSS.n3865 VSS.n3470 0.00764286
R25127 VSS.n3897 VSS.n3456 0.00764286
R25128 VSS.n3949 VSS.n3437 0.00764286
R25129 VSS.n3982 VSS.n3420 0.00764286
R25130 VSS.n3978 VSS.n3420 0.00764286
R25131 VSS.n3862 VSS.n3861 0.00764286
R25132 VSS.n3862 VSS.n3475 0.00764286
R25133 VSS.n3868 VSS.n3476 0.00764286
R25134 VSS.n3864 VSS.n3472 0.00764286
R25135 VSS.n3883 VSS.n3882 0.00764286
R25136 VSS.n3898 VSS.n3455 0.00764286
R25137 VSS.n3920 VSS.n3919 0.00764286
R25138 VSS.n3956 VSS.n3433 0.00764286
R25139 VSS.n3981 VSS.n3980 0.00764286
R25140 VSS.n3980 VSS.n3979 0.00764286
R25141 VSS.n3673 VSS.n3600 0.00764286
R25142 VSS.n3681 VSS.n3680 0.00764286
R25143 VSS.n3585 VSS.n3584 0.00764286
R25144 VSS.n3704 VSS.n3575 0.00764286
R25145 VSS.n3731 VSS.n3555 0.00764286
R25146 VSS.n4178 VSS.n4172 0.00764286
R25147 VSS.n4351 VSS.n4125 0.00764286
R25148 VSS.n4389 VSS.n4097 0.00764286
R25149 VSS.n4326 VSS.n4136 0.00764286
R25150 VSS.n4354 VSS.n4353 0.00764286
R25151 VSS.n4361 VSS.n4118 0.00764286
R25152 VSS.n4357 VSS.n4356 0.00764286
R25153 VSS.n4379 VSS.n4104 0.00764286
R25154 VSS.n4393 VSS.n4098 0.00764286
R25155 VSS.n4459 VSS.n4458 0.00764286
R25156 VSS.n4457 VSS.n4062 0.00764286
R25157 VSS.n4489 VSS.n4048 0.00764286
R25158 VSS.n4541 VSS.n4029 0.00764286
R25159 VSS.n4574 VSS.n4012 0.00764286
R25160 VSS.n4570 VSS.n4012 0.00764286
R25161 VSS.n4454 VSS.n4453 0.00764286
R25162 VSS.n4454 VSS.n4067 0.00764286
R25163 VSS.n4460 VSS.n4068 0.00764286
R25164 VSS.n4456 VSS.n4064 0.00764286
R25165 VSS.n4475 VSS.n4474 0.00764286
R25166 VSS.n4490 VSS.n4047 0.00764286
R25167 VSS.n4512 VSS.n4511 0.00764286
R25168 VSS.n4548 VSS.n4025 0.00764286
R25169 VSS.n4573 VSS.n4572 0.00764286
R25170 VSS.n4572 VSS.n4571 0.00764286
R25171 VSS.n4265 VSS.n4192 0.00764286
R25172 VSS.n4273 VSS.n4272 0.00764286
R25173 VSS.n4177 VSS.n4176 0.00764286
R25174 VSS.n4296 VSS.n4167 0.00764286
R25175 VSS.n4323 VSS.n4147 0.00764286
R25176 VSS.n4770 VSS.n4764 0.00764286
R25177 VSS.n4943 VSS.n4717 0.00764286
R25178 VSS.n4981 VSS.n4689 0.00764286
R25179 VSS.n4918 VSS.n4728 0.00764286
R25180 VSS.n4946 VSS.n4945 0.00764286
R25181 VSS.n4953 VSS.n4710 0.00764286
R25182 VSS.n4949 VSS.n4948 0.00764286
R25183 VSS.n4971 VSS.n4696 0.00764286
R25184 VSS.n4985 VSS.n4690 0.00764286
R25185 VSS.n5051 VSS.n5050 0.00764286
R25186 VSS.n5049 VSS.n4654 0.00764286
R25187 VSS.n5081 VSS.n4640 0.00764286
R25188 VSS.n5133 VSS.n4621 0.00764286
R25189 VSS.n5166 VSS.n4604 0.00764286
R25190 VSS.n5162 VSS.n4604 0.00764286
R25191 VSS.n5046 VSS.n5045 0.00764286
R25192 VSS.n5046 VSS.n4659 0.00764286
R25193 VSS.n5052 VSS.n4660 0.00764286
R25194 VSS.n5048 VSS.n4656 0.00764286
R25195 VSS.n5067 VSS.n5066 0.00764286
R25196 VSS.n5082 VSS.n4639 0.00764286
R25197 VSS.n5104 VSS.n5103 0.00764286
R25198 VSS.n5140 VSS.n4617 0.00764286
R25199 VSS.n5165 VSS.n5164 0.00764286
R25200 VSS.n5164 VSS.n5163 0.00764286
R25201 VSS.n4857 VSS.n4784 0.00764286
R25202 VSS.n4865 VSS.n4864 0.00764286
R25203 VSS.n4769 VSS.n4768 0.00764286
R25204 VSS.n4888 VSS.n4759 0.00764286
R25205 VSS.n4915 VSS.n4739 0.00764286
R25206 VSS.n2391 VSS.n2385 0.00764286
R25207 VSS.n2618 VSS.n2617 0.00764286
R25208 VSS.n2641 VSS.n2640 0.00764286
R25209 VSS.n5310 VSS.n5309 0.00764286
R25210 VSS.n5301 VSS.n2545 0.00764286
R25211 VSS.n2615 VSS.n2547 0.00764286
R25212 VSS.n2552 VSS.n2551 0.00764286
R25213 VSS.n2560 VSS.n2559 0.00764286
R25214 VSS.n2643 VSS.n2561 0.00764286
R25215 VSS.n2694 VSS.n2693 0.00764286
R25216 VSS.n5256 VSS.n2675 0.00764286
R25217 VSS.n5236 VSS.n2705 0.00764286
R25218 VSS.n5216 VSS.n2752 0.00764286
R25219 VSS.n2807 VSS.n2768 0.00764286
R25220 VSS.n2808 VSS.n2807 0.00764286
R25221 VSS.n2691 VSS.n2690 0.00764286
R25222 VSS.n2691 VSS.n2680 0.00764286
R25223 VSS.n2695 VSS.n2681 0.00764286
R25224 VSS.n5255 VSS.n2677 0.00764286
R25225 VSS.n5239 VSS.n2706 0.00764286
R25226 VSS.n5238 VSS.n5237 0.00764286
R25227 VSS.n2761 VSS.n2750 0.00764286
R25228 VSS.n5210 VSS.n5209 0.00764286
R25229 VSS.n2806 VSS.n2805 0.00764286
R25230 VSS.n2806 VSS.n2804 0.00764286
R25231 VSS.n2478 VSS.n2405 0.00764286
R25232 VSS.n2486 VSS.n2485 0.00764286
R25233 VSS.n2390 VSS.n2389 0.00764286
R25234 VSS.n2509 VSS.n2380 0.00764286
R25235 VSS.n2536 VSS.n2360 0.00764286
R25236 VSS.n5352 VSS.n5346 0.00764286
R25237 VSS.n5579 VSS.n5578 0.00764286
R25238 VSS.n5602 VSS.n5601 0.00764286
R25239 VSS.n5883 VSS.n5882 0.00764286
R25240 VSS.n5874 VSS.n5506 0.00764286
R25241 VSS.n5576 VSS.n5508 0.00764286
R25242 VSS.n5513 VSS.n5512 0.00764286
R25243 VSS.n5521 VSS.n5520 0.00764286
R25244 VSS.n5604 VSS.n5522 0.00764286
R25245 VSS.n5655 VSS.n5654 0.00764286
R25246 VSS.n5829 VSS.n5636 0.00764286
R25247 VSS.n5809 VSS.n5666 0.00764286
R25248 VSS.n5789 VSS.n5713 0.00764286
R25249 VSS.n5741 VSS.n5729 0.00764286
R25250 VSS.n5737 VSS.n5729 0.00764286
R25251 VSS.n5652 VSS.n5651 0.00764286
R25252 VSS.n5652 VSS.n5641 0.00764286
R25253 VSS.n5656 VSS.n5642 0.00764286
R25254 VSS.n5828 VSS.n5638 0.00764286
R25255 VSS.n5812 VSS.n5667 0.00764286
R25256 VSS.n5811 VSS.n5810 0.00764286
R25257 VSS.n5722 VSS.n5711 0.00764286
R25258 VSS.n5783 VSS.n5782 0.00764286
R25259 VSS.n5740 VSS.n5739 0.00764286
R25260 VSS.n5739 VSS.n5738 0.00764286
R25261 VSS.n5439 VSS.n5366 0.00764286
R25262 VSS.n5447 VSS.n5446 0.00764286
R25263 VSS.n5351 VSS.n5350 0.00764286
R25264 VSS.n5470 VSS.n5341 0.00764286
R25265 VSS.n5497 VSS.n5321 0.00764286
R25266 VSS.n5925 VSS.n5919 0.00764286
R25267 VSS.n6152 VSS.n6151 0.00764286
R25268 VSS.n6175 VSS.n6174 0.00764286
R25269 VSS.n6475 VSS.n6474 0.00764286
R25270 VSS.n6466 VSS.n6079 0.00764286
R25271 VSS.n6149 VSS.n6081 0.00764286
R25272 VSS.n6086 VSS.n6085 0.00764286
R25273 VSS.n6094 VSS.n6093 0.00764286
R25274 VSS.n6177 VSS.n6095 0.00764286
R25275 VSS.n6228 VSS.n6227 0.00764286
R25276 VSS.n6421 VSS.n6209 0.00764286
R25277 VSS.n6401 VSS.n6239 0.00764286
R25278 VSS.n6381 VSS.n6286 0.00764286
R25279 VSS.n6341 VSS.n6302 0.00764286
R25280 VSS.n6342 VSS.n6341 0.00764286
R25281 VSS.n6225 VSS.n6224 0.00764286
R25282 VSS.n6225 VSS.n6214 0.00764286
R25283 VSS.n6229 VSS.n6215 0.00764286
R25284 VSS.n6420 VSS.n6211 0.00764286
R25285 VSS.n6404 VSS.n6240 0.00764286
R25286 VSS.n6403 VSS.n6402 0.00764286
R25287 VSS.n6295 VSS.n6284 0.00764286
R25288 VSS.n6375 VSS.n6374 0.00764286
R25289 VSS.n6340 VSS.n6339 0.00764286
R25290 VSS.n6340 VSS.n6338 0.00764286
R25291 VSS.n6012 VSS.n5939 0.00764286
R25292 VSS.n6020 VSS.n6019 0.00764286
R25293 VSS.n5924 VSS.n5923 0.00764286
R25294 VSS.n6043 VSS.n5914 0.00764286
R25295 VSS.n6070 VSS.n5894 0.00764286
R25296 VSS.n7727 VSS.n7721 0.00764286
R25297 VSS.n7900 VSS.n7674 0.00764286
R25298 VSS.n7938 VSS.n7646 0.00764286
R25299 VSS.n7875 VSS.n7685 0.00764286
R25300 VSS.n7903 VSS.n7902 0.00764286
R25301 VSS.n7910 VSS.n7667 0.00764286
R25302 VSS.n7906 VSS.n7905 0.00764286
R25303 VSS.n7928 VSS.n7653 0.00764286
R25304 VSS.n7942 VSS.n7647 0.00764286
R25305 VSS.n8008 VSS.n8007 0.00764286
R25306 VSS.n8006 VSS.n7611 0.00764286
R25307 VSS.n8038 VSS.n7597 0.00764286
R25308 VSS.n8090 VSS.n7578 0.00764286
R25309 VSS.n8123 VSS.n7561 0.00764286
R25310 VSS.n8119 VSS.n7561 0.00764286
R25311 VSS.n8003 VSS.n8002 0.00764286
R25312 VSS.n8003 VSS.n7616 0.00764286
R25313 VSS.n8009 VSS.n7617 0.00764286
R25314 VSS.n8005 VSS.n7613 0.00764286
R25315 VSS.n8024 VSS.n8023 0.00764286
R25316 VSS.n8039 VSS.n7596 0.00764286
R25317 VSS.n8061 VSS.n8060 0.00764286
R25318 VSS.n8097 VSS.n7574 0.00764286
R25319 VSS.n8122 VSS.n8121 0.00764286
R25320 VSS.n8121 VSS.n8120 0.00764286
R25321 VSS.n7814 VSS.n7741 0.00764286
R25322 VSS.n7822 VSS.n7821 0.00764286
R25323 VSS.n7726 VSS.n7725 0.00764286
R25324 VSS.n7845 VSS.n7716 0.00764286
R25325 VSS.n7872 VSS.n7696 0.00764286
R25326 VSS.n8319 VSS.n8313 0.00764286
R25327 VSS.n8492 VSS.n8266 0.00764286
R25328 VSS.n8530 VSS.n8238 0.00764286
R25329 VSS.n8467 VSS.n8277 0.00764286
R25330 VSS.n8495 VSS.n8494 0.00764286
R25331 VSS.n8502 VSS.n8259 0.00764286
R25332 VSS.n8498 VSS.n8497 0.00764286
R25333 VSS.n8520 VSS.n8245 0.00764286
R25334 VSS.n8534 VSS.n8239 0.00764286
R25335 VSS.n8600 VSS.n8599 0.00764286
R25336 VSS.n8598 VSS.n8203 0.00764286
R25337 VSS.n8630 VSS.n8189 0.00764286
R25338 VSS.n8682 VSS.n8170 0.00764286
R25339 VSS.n8715 VSS.n8153 0.00764286
R25340 VSS.n8711 VSS.n8153 0.00764286
R25341 VSS.n8595 VSS.n8594 0.00764286
R25342 VSS.n8595 VSS.n8208 0.00764286
R25343 VSS.n8601 VSS.n8209 0.00764286
R25344 VSS.n8597 VSS.n8205 0.00764286
R25345 VSS.n8616 VSS.n8615 0.00764286
R25346 VSS.n8631 VSS.n8188 0.00764286
R25347 VSS.n8653 VSS.n8652 0.00764286
R25348 VSS.n8689 VSS.n8166 0.00764286
R25349 VSS.n8714 VSS.n8713 0.00764286
R25350 VSS.n8713 VSS.n8712 0.00764286
R25351 VSS.n8406 VSS.n8333 0.00764286
R25352 VSS.n8414 VSS.n8413 0.00764286
R25353 VSS.n8318 VSS.n8317 0.00764286
R25354 VSS.n8437 VSS.n8308 0.00764286
R25355 VSS.n8464 VSS.n8288 0.00764286
R25356 VSS.n8911 VSS.n8905 0.00764286
R25357 VSS.n9084 VSS.n8858 0.00764286
R25358 VSS.n9122 VSS.n8830 0.00764286
R25359 VSS.n9059 VSS.n8869 0.00764286
R25360 VSS.n9087 VSS.n9086 0.00764286
R25361 VSS.n9094 VSS.n8851 0.00764286
R25362 VSS.n9090 VSS.n9089 0.00764286
R25363 VSS.n9112 VSS.n8837 0.00764286
R25364 VSS.n9126 VSS.n8831 0.00764286
R25365 VSS.n9192 VSS.n9191 0.00764286
R25366 VSS.n9190 VSS.n8795 0.00764286
R25367 VSS.n9222 VSS.n8781 0.00764286
R25368 VSS.n9274 VSS.n8762 0.00764286
R25369 VSS.n9307 VSS.n8745 0.00764286
R25370 VSS.n9303 VSS.n8745 0.00764286
R25371 VSS.n9187 VSS.n9186 0.00764286
R25372 VSS.n9187 VSS.n8800 0.00764286
R25373 VSS.n9193 VSS.n8801 0.00764286
R25374 VSS.n9189 VSS.n8797 0.00764286
R25375 VSS.n9208 VSS.n9207 0.00764286
R25376 VSS.n9223 VSS.n8780 0.00764286
R25377 VSS.n9245 VSS.n9244 0.00764286
R25378 VSS.n9281 VSS.n8758 0.00764286
R25379 VSS.n9306 VSS.n9305 0.00764286
R25380 VSS.n9305 VSS.n9304 0.00764286
R25381 VSS.n8998 VSS.n8925 0.00764286
R25382 VSS.n9006 VSS.n9005 0.00764286
R25383 VSS.n8910 VSS.n8909 0.00764286
R25384 VSS.n9029 VSS.n8900 0.00764286
R25385 VSS.n9056 VSS.n8880 0.00764286
R25386 VSS.n10095 VSS.n10089 0.00764286
R25387 VSS.n10268 VSS.n10042 0.00764286
R25388 VSS.n10306 VSS.n10014 0.00764286
R25389 VSS.n10243 VSS.n10053 0.00764286
R25390 VSS.n10271 VSS.n10270 0.00764286
R25391 VSS.n10278 VSS.n10035 0.00764286
R25392 VSS.n10274 VSS.n10273 0.00764286
R25393 VSS.n10296 VSS.n10021 0.00764286
R25394 VSS.n10310 VSS.n10015 0.00764286
R25395 VSS.n10376 VSS.n10375 0.00764286
R25396 VSS.n10374 VSS.n9979 0.00764286
R25397 VSS.n10406 VSS.n9965 0.00764286
R25398 VSS.n10458 VSS.n9946 0.00764286
R25399 VSS.n10491 VSS.n9929 0.00764286
R25400 VSS.n10487 VSS.n9929 0.00764286
R25401 VSS.n10371 VSS.n10370 0.00764286
R25402 VSS.n10371 VSS.n9984 0.00764286
R25403 VSS.n10377 VSS.n9985 0.00764286
R25404 VSS.n10373 VSS.n9981 0.00764286
R25405 VSS.n10392 VSS.n10391 0.00764286
R25406 VSS.n10407 VSS.n9964 0.00764286
R25407 VSS.n10429 VSS.n10428 0.00764286
R25408 VSS.n10465 VSS.n9942 0.00764286
R25409 VSS.n10490 VSS.n10489 0.00764286
R25410 VSS.n10489 VSS.n10488 0.00764286
R25411 VSS.n10182 VSS.n10109 0.00764286
R25412 VSS.n10190 VSS.n10189 0.00764286
R25413 VSS.n10094 VSS.n10093 0.00764286
R25414 VSS.n10213 VSS.n10084 0.00764286
R25415 VSS.n10240 VSS.n10064 0.00764286
R25416 VSS.n10687 VSS.n10681 0.00764286
R25417 VSS.n10860 VSS.n10634 0.00764286
R25418 VSS.n10898 VSS.n10606 0.00764286
R25419 VSS.n10835 VSS.n10645 0.00764286
R25420 VSS.n10863 VSS.n10862 0.00764286
R25421 VSS.n10870 VSS.n10627 0.00764286
R25422 VSS.n10866 VSS.n10865 0.00764286
R25423 VSS.n10888 VSS.n10613 0.00764286
R25424 VSS.n10902 VSS.n10607 0.00764286
R25425 VSS.n10968 VSS.n10967 0.00764286
R25426 VSS.n10966 VSS.n10571 0.00764286
R25427 VSS.n10998 VSS.n10557 0.00764286
R25428 VSS.n11050 VSS.n10538 0.00764286
R25429 VSS.n11083 VSS.n10521 0.00764286
R25430 VSS.n11079 VSS.n10521 0.00764286
R25431 VSS.n10963 VSS.n10962 0.00764286
R25432 VSS.n10963 VSS.n10576 0.00764286
R25433 VSS.n10969 VSS.n10577 0.00764286
R25434 VSS.n10965 VSS.n10573 0.00764286
R25435 VSS.n10984 VSS.n10983 0.00764286
R25436 VSS.n10999 VSS.n10556 0.00764286
R25437 VSS.n11021 VSS.n11020 0.00764286
R25438 VSS.n11057 VSS.n10534 0.00764286
R25439 VSS.n11082 VSS.n11081 0.00764286
R25440 VSS.n11081 VSS.n11080 0.00764286
R25441 VSS.n10774 VSS.n10701 0.00764286
R25442 VSS.n10782 VSS.n10781 0.00764286
R25443 VSS.n10686 VSS.n10685 0.00764286
R25444 VSS.n10805 VSS.n10676 0.00764286
R25445 VSS.n10832 VSS.n10656 0.00764286
R25446 VSS.n11279 VSS.n11273 0.00764286
R25447 VSS.n11452 VSS.n11226 0.00764286
R25448 VSS.n11490 VSS.n11198 0.00764286
R25449 VSS.n11427 VSS.n11237 0.00764286
R25450 VSS.n11455 VSS.n11454 0.00764286
R25451 VSS.n11462 VSS.n11219 0.00764286
R25452 VSS.n11458 VSS.n11457 0.00764286
R25453 VSS.n11480 VSS.n11205 0.00764286
R25454 VSS.n11494 VSS.n11199 0.00764286
R25455 VSS.n11560 VSS.n11559 0.00764286
R25456 VSS.n11558 VSS.n11163 0.00764286
R25457 VSS.n11590 VSS.n11149 0.00764286
R25458 VSS.n11642 VSS.n11130 0.00764286
R25459 VSS.n11675 VSS.n11113 0.00764286
R25460 VSS.n11671 VSS.n11113 0.00764286
R25461 VSS.n11555 VSS.n11554 0.00764286
R25462 VSS.n11555 VSS.n11168 0.00764286
R25463 VSS.n11561 VSS.n11169 0.00764286
R25464 VSS.n11557 VSS.n11165 0.00764286
R25465 VSS.n11576 VSS.n11575 0.00764286
R25466 VSS.n11591 VSS.n11148 0.00764286
R25467 VSS.n11613 VSS.n11612 0.00764286
R25468 VSS.n11649 VSS.n11126 0.00764286
R25469 VSS.n11674 VSS.n11673 0.00764286
R25470 VSS.n11673 VSS.n11672 0.00764286
R25471 VSS.n11366 VSS.n11293 0.00764286
R25472 VSS.n11374 VSS.n11373 0.00764286
R25473 VSS.n11278 VSS.n11277 0.00764286
R25474 VSS.n11397 VSS.n11268 0.00764286
R25475 VSS.n11424 VSS.n11248 0.00764286
R25476 VSS.n11871 VSS.n11865 0.00764286
R25477 VSS.n12044 VSS.n11818 0.00764286
R25478 VSS.n12082 VSS.n11790 0.00764286
R25479 VSS.n12019 VSS.n11829 0.00764286
R25480 VSS.n12047 VSS.n12046 0.00764286
R25481 VSS.n12054 VSS.n11811 0.00764286
R25482 VSS.n12050 VSS.n12049 0.00764286
R25483 VSS.n12072 VSS.n11797 0.00764286
R25484 VSS.n12086 VSS.n11791 0.00764286
R25485 VSS.n12152 VSS.n12151 0.00764286
R25486 VSS.n12150 VSS.n11755 0.00764286
R25487 VSS.n12182 VSS.n11741 0.00764286
R25488 VSS.n12234 VSS.n11722 0.00764286
R25489 VSS.n12267 VSS.n11705 0.00764286
R25490 VSS.n12263 VSS.n11705 0.00764286
R25491 VSS.n12147 VSS.n12146 0.00764286
R25492 VSS.n12147 VSS.n11760 0.00764286
R25493 VSS.n12153 VSS.n11761 0.00764286
R25494 VSS.n12149 VSS.n11757 0.00764286
R25495 VSS.n12168 VSS.n12167 0.00764286
R25496 VSS.n12183 VSS.n11740 0.00764286
R25497 VSS.n12205 VSS.n12204 0.00764286
R25498 VSS.n12241 VSS.n11718 0.00764286
R25499 VSS.n12266 VSS.n12265 0.00764286
R25500 VSS.n12265 VSS.n12264 0.00764286
R25501 VSS.n11958 VSS.n11885 0.00764286
R25502 VSS.n11966 VSS.n11965 0.00764286
R25503 VSS.n11870 VSS.n11869 0.00764286
R25504 VSS.n11989 VSS.n11860 0.00764286
R25505 VSS.n12016 VSS.n11840 0.00764286
R25506 VSS.n12463 VSS.n12457 0.00764286
R25507 VSS.n12636 VSS.n12410 0.00764286
R25508 VSS.n12674 VSS.n12382 0.00764286
R25509 VSS.n12611 VSS.n12421 0.00764286
R25510 VSS.n12639 VSS.n12638 0.00764286
R25511 VSS.n12646 VSS.n12403 0.00764286
R25512 VSS.n12642 VSS.n12641 0.00764286
R25513 VSS.n12664 VSS.n12389 0.00764286
R25514 VSS.n12678 VSS.n12383 0.00764286
R25515 VSS.n12744 VSS.n12743 0.00764286
R25516 VSS.n12742 VSS.n12347 0.00764286
R25517 VSS.n12774 VSS.n12333 0.00764286
R25518 VSS.n12826 VSS.n12314 0.00764286
R25519 VSS.n12859 VSS.n12297 0.00764286
R25520 VSS.n12855 VSS.n12297 0.00764286
R25521 VSS.n12739 VSS.n12738 0.00764286
R25522 VSS.n12739 VSS.n12352 0.00764286
R25523 VSS.n12745 VSS.n12353 0.00764286
R25524 VSS.n12741 VSS.n12349 0.00764286
R25525 VSS.n12760 VSS.n12759 0.00764286
R25526 VSS.n12775 VSS.n12332 0.00764286
R25527 VSS.n12797 VSS.n12796 0.00764286
R25528 VSS.n12833 VSS.n12310 0.00764286
R25529 VSS.n12858 VSS.n12857 0.00764286
R25530 VSS.n12857 VSS.n12856 0.00764286
R25531 VSS.n12550 VSS.n12477 0.00764286
R25532 VSS.n12558 VSS.n12557 0.00764286
R25533 VSS.n12462 VSS.n12461 0.00764286
R25534 VSS.n12581 VSS.n12452 0.00764286
R25535 VSS.n12608 VSS.n12432 0.00764286
R25536 VSS.n13055 VSS.n13049 0.00764286
R25537 VSS.n13228 VSS.n13002 0.00764286
R25538 VSS.n13266 VSS.n12974 0.00764286
R25539 VSS.n13203 VSS.n13013 0.00764286
R25540 VSS.n13231 VSS.n13230 0.00764286
R25541 VSS.n13238 VSS.n12995 0.00764286
R25542 VSS.n13234 VSS.n13233 0.00764286
R25543 VSS.n13256 VSS.n12981 0.00764286
R25544 VSS.n13270 VSS.n12975 0.00764286
R25545 VSS.n13336 VSS.n13335 0.00764286
R25546 VSS.n13334 VSS.n12939 0.00764286
R25547 VSS.n13366 VSS.n12925 0.00764286
R25548 VSS.n13418 VSS.n12906 0.00764286
R25549 VSS.n13451 VSS.n12889 0.00764286
R25550 VSS.n13447 VSS.n12889 0.00764286
R25551 VSS.n13331 VSS.n13330 0.00764286
R25552 VSS.n13331 VSS.n12944 0.00764286
R25553 VSS.n13337 VSS.n12945 0.00764286
R25554 VSS.n13333 VSS.n12941 0.00764286
R25555 VSS.n13352 VSS.n13351 0.00764286
R25556 VSS.n13367 VSS.n12924 0.00764286
R25557 VSS.n13389 VSS.n13388 0.00764286
R25558 VSS.n13425 VSS.n12902 0.00764286
R25559 VSS.n13450 VSS.n13449 0.00764286
R25560 VSS.n13449 VSS.n13448 0.00764286
R25561 VSS.n13142 VSS.n13069 0.00764286
R25562 VSS.n13150 VSS.n13149 0.00764286
R25563 VSS.n13054 VSS.n13053 0.00764286
R25564 VSS.n13173 VSS.n13044 0.00764286
R25565 VSS.n13200 VSS.n13024 0.00764286
R25566 VSS.n13647 VSS.n13641 0.00764286
R25567 VSS.n13820 VSS.n13594 0.00764286
R25568 VSS.n13858 VSS.n13566 0.00764286
R25569 VSS.n13795 VSS.n13605 0.00764286
R25570 VSS.n13823 VSS.n13822 0.00764286
R25571 VSS.n13830 VSS.n13587 0.00764286
R25572 VSS.n13826 VSS.n13825 0.00764286
R25573 VSS.n13848 VSS.n13573 0.00764286
R25574 VSS.n13862 VSS.n13567 0.00764286
R25575 VSS.n13928 VSS.n13927 0.00764286
R25576 VSS.n13926 VSS.n13531 0.00764286
R25577 VSS.n13958 VSS.n13517 0.00764286
R25578 VSS.n14010 VSS.n13498 0.00764286
R25579 VSS.n14043 VSS.n13481 0.00764286
R25580 VSS.n14039 VSS.n13481 0.00764286
R25581 VSS.n13923 VSS.n13922 0.00764286
R25582 VSS.n13923 VSS.n13536 0.00764286
R25583 VSS.n13929 VSS.n13537 0.00764286
R25584 VSS.n13925 VSS.n13533 0.00764286
R25585 VSS.n13944 VSS.n13943 0.00764286
R25586 VSS.n13959 VSS.n13516 0.00764286
R25587 VSS.n13981 VSS.n13980 0.00764286
R25588 VSS.n14017 VSS.n13494 0.00764286
R25589 VSS.n14042 VSS.n14041 0.00764286
R25590 VSS.n14041 VSS.n14040 0.00764286
R25591 VSS.n13734 VSS.n13661 0.00764286
R25592 VSS.n13742 VSS.n13741 0.00764286
R25593 VSS.n13646 VSS.n13645 0.00764286
R25594 VSS.n13765 VSS.n13636 0.00764286
R25595 VSS.n13792 VSS.n13616 0.00764286
R25596 VSS.n14239 VSS.n14233 0.00764286
R25597 VSS.n14412 VSS.n14186 0.00764286
R25598 VSS.n14450 VSS.n14158 0.00764286
R25599 VSS.n14387 VSS.n14197 0.00764286
R25600 VSS.n14415 VSS.n14414 0.00764286
R25601 VSS.n14422 VSS.n14179 0.00764286
R25602 VSS.n14418 VSS.n14417 0.00764286
R25603 VSS.n14440 VSS.n14165 0.00764286
R25604 VSS.n14454 VSS.n14159 0.00764286
R25605 VSS.n14520 VSS.n14519 0.00764286
R25606 VSS.n14518 VSS.n14123 0.00764286
R25607 VSS.n14550 VSS.n14109 0.00764286
R25608 VSS.n14602 VSS.n14090 0.00764286
R25609 VSS.n14635 VSS.n14073 0.00764286
R25610 VSS.n14631 VSS.n14073 0.00764286
R25611 VSS.n14515 VSS.n14514 0.00764286
R25612 VSS.n14515 VSS.n14128 0.00764286
R25613 VSS.n14521 VSS.n14129 0.00764286
R25614 VSS.n14517 VSS.n14125 0.00764286
R25615 VSS.n14536 VSS.n14535 0.00764286
R25616 VSS.n14551 VSS.n14108 0.00764286
R25617 VSS.n14573 VSS.n14572 0.00764286
R25618 VSS.n14609 VSS.n14086 0.00764286
R25619 VSS.n14634 VSS.n14633 0.00764286
R25620 VSS.n14633 VSS.n14632 0.00764286
R25621 VSS.n14326 VSS.n14253 0.00764286
R25622 VSS.n14334 VSS.n14333 0.00764286
R25623 VSS.n14238 VSS.n14237 0.00764286
R25624 VSS.n14357 VSS.n14228 0.00764286
R25625 VSS.n14384 VSS.n14208 0.00764286
R25626 VSS.n14831 VSS.n14825 0.00764286
R25627 VSS.n15004 VSS.n14778 0.00764286
R25628 VSS.n15042 VSS.n14750 0.00764286
R25629 VSS.n14979 VSS.n14789 0.00764286
R25630 VSS.n15007 VSS.n15006 0.00764286
R25631 VSS.n15014 VSS.n14771 0.00764286
R25632 VSS.n15010 VSS.n15009 0.00764286
R25633 VSS.n15032 VSS.n14757 0.00764286
R25634 VSS.n15046 VSS.n14751 0.00764286
R25635 VSS.n15112 VSS.n15111 0.00764286
R25636 VSS.n15110 VSS.n14715 0.00764286
R25637 VSS.n15142 VSS.n14701 0.00764286
R25638 VSS.n15194 VSS.n14682 0.00764286
R25639 VSS.n15227 VSS.n14665 0.00764286
R25640 VSS.n15223 VSS.n14665 0.00764286
R25641 VSS.n15107 VSS.n15106 0.00764286
R25642 VSS.n15107 VSS.n14720 0.00764286
R25643 VSS.n15113 VSS.n14721 0.00764286
R25644 VSS.n15109 VSS.n14717 0.00764286
R25645 VSS.n15128 VSS.n15127 0.00764286
R25646 VSS.n15143 VSS.n14700 0.00764286
R25647 VSS.n15165 VSS.n15164 0.00764286
R25648 VSS.n15201 VSS.n14678 0.00764286
R25649 VSS.n15226 VSS.n15225 0.00764286
R25650 VSS.n15225 VSS.n15224 0.00764286
R25651 VSS.n14918 VSS.n14845 0.00764286
R25652 VSS.n14926 VSS.n14925 0.00764286
R25653 VSS.n14830 VSS.n14829 0.00764286
R25654 VSS.n14949 VSS.n14820 0.00764286
R25655 VSS.n14976 VSS.n14800 0.00764286
R25656 VSS.n15423 VSS.n15417 0.00764286
R25657 VSS.n15596 VSS.n15370 0.00764286
R25658 VSS.n15634 VSS.n15342 0.00764286
R25659 VSS.n15571 VSS.n15381 0.00764286
R25660 VSS.n15599 VSS.n15598 0.00764286
R25661 VSS.n15606 VSS.n15363 0.00764286
R25662 VSS.n15602 VSS.n15601 0.00764286
R25663 VSS.n15624 VSS.n15349 0.00764286
R25664 VSS.n15638 VSS.n15343 0.00764286
R25665 VSS.n15704 VSS.n15703 0.00764286
R25666 VSS.n15702 VSS.n15307 0.00764286
R25667 VSS.n15734 VSS.n15293 0.00764286
R25668 VSS.n15786 VSS.n15274 0.00764286
R25669 VSS.n15819 VSS.n15257 0.00764286
R25670 VSS.n15815 VSS.n15257 0.00764286
R25671 VSS.n15699 VSS.n15698 0.00764286
R25672 VSS.n15699 VSS.n15312 0.00764286
R25673 VSS.n15705 VSS.n15313 0.00764286
R25674 VSS.n15701 VSS.n15309 0.00764286
R25675 VSS.n15720 VSS.n15719 0.00764286
R25676 VSS.n15735 VSS.n15292 0.00764286
R25677 VSS.n15757 VSS.n15756 0.00764286
R25678 VSS.n15793 VSS.n15270 0.00764286
R25679 VSS.n15818 VSS.n15817 0.00764286
R25680 VSS.n15817 VSS.n15816 0.00764286
R25681 VSS.n15510 VSS.n15437 0.00764286
R25682 VSS.n15518 VSS.n15517 0.00764286
R25683 VSS.n15422 VSS.n15421 0.00764286
R25684 VSS.n15541 VSS.n15412 0.00764286
R25685 VSS.n15568 VSS.n15392 0.00764286
R25686 VSS.n6531 VSS.n6525 0.00764286
R25687 VSS.n6758 VSS.n6757 0.00764286
R25688 VSS.n6781 VSS.n6780 0.00764286
R25689 VSS.n15963 VSS.n15962 0.00764286
R25690 VSS.n15954 VSS.n6685 0.00764286
R25691 VSS.n6755 VSS.n6687 0.00764286
R25692 VSS.n6692 VSS.n6691 0.00764286
R25693 VSS.n6700 VSS.n6699 0.00764286
R25694 VSS.n6783 VSS.n6701 0.00764286
R25695 VSS.n6834 VSS.n6833 0.00764286
R25696 VSS.n15909 VSS.n6815 0.00764286
R25697 VSS.n15889 VSS.n6845 0.00764286
R25698 VSS.n15869 VSS.n6892 0.00764286
R25699 VSS.n6947 VSS.n6908 0.00764286
R25700 VSS.n6948 VSS.n6947 0.00764286
R25701 VSS.n6831 VSS.n6830 0.00764286
R25702 VSS.n6831 VSS.n6820 0.00764286
R25703 VSS.n6835 VSS.n6821 0.00764286
R25704 VSS.n15908 VSS.n6817 0.00764286
R25705 VSS.n15892 VSS.n6846 0.00764286
R25706 VSS.n15891 VSS.n15890 0.00764286
R25707 VSS.n6901 VSS.n6890 0.00764286
R25708 VSS.n15863 VSS.n15862 0.00764286
R25709 VSS.n6946 VSS.n6945 0.00764286
R25710 VSS.n6946 VSS.n6944 0.00764286
R25711 VSS.n6618 VSS.n6545 0.00764286
R25712 VSS.n6626 VSS.n6625 0.00764286
R25713 VSS.n6530 VSS.n6529 0.00764286
R25714 VSS.n6649 VSS.n6520 0.00764286
R25715 VSS.n6676 VSS.n6500 0.00764286
R25716 VSS.n7246 VSS.n7128 0.00764286
R25717 VSS.n7308 VSS.n7081 0.00764286
R25718 VSS.n7346 VSS.n7053 0.00764286
R25719 VSS.n7283 VSS.n7092 0.00764286
R25720 VSS.n7311 VSS.n7310 0.00764286
R25721 VSS.n7318 VSS.n7074 0.00764286
R25722 VSS.n7314 VSS.n7313 0.00764286
R25723 VSS.n7336 VSS.n7060 0.00764286
R25724 VSS.n7350 VSS.n7054 0.00764286
R25725 VSS.n7416 VSS.n7415 0.00764286
R25726 VSS.n7414 VSS.n7018 0.00764286
R25727 VSS.n7446 VSS.n7004 0.00764286
R25728 VSS.n7498 VSS.n6985 0.00764286
R25729 VSS.n7531 VSS.n6968 0.00764286
R25730 VSS.n7527 VSS.n6968 0.00764286
R25731 VSS.n7411 VSS.n7410 0.00764286
R25732 VSS.n7411 VSS.n7023 0.00764286
R25733 VSS.n7417 VSS.n7024 0.00764286
R25734 VSS.n7413 VSS.n7020 0.00764286
R25735 VSS.n7432 VSS.n7431 0.00764286
R25736 VSS.n7447 VSS.n7003 0.00764286
R25737 VSS.n7469 VSS.n7468 0.00764286
R25738 VSS.n7505 VSS.n6981 0.00764286
R25739 VSS.n7530 VSS.n7529 0.00764286
R25740 VSS.n7529 VSS.n7528 0.00764286
R25741 VSS.n7209 VSS.n7208 0.00764286
R25742 VSS.n7231 VSS.n7135 0.00764286
R25743 VSS.n7245 VSS.n7244 0.00764286
R25744 VSS.n7243 VSS.n7239 0.00764286
R25745 VSS.n7280 VSS.n7103 0.00764286
R25746 VSS.n391 VSS.n388 0.00764286
R25747 VSS.n18620 VSS.n179 0.00764286
R25748 VSS.n18658 VSS.n151 0.00764286
R25749 VSS.n18595 VSS.n190 0.00764286
R25750 VSS.n18623 VSS.n18622 0.00764286
R25751 VSS.n18630 VSS.n172 0.00764286
R25752 VSS.n18626 VSS.n18625 0.00764286
R25753 VSS.n18648 VSS.n158 0.00764286
R25754 VSS.n18662 VSS.n152 0.00764286
R25755 VSS.n18728 VSS.n18727 0.00764286
R25756 VSS.n18726 VSS.n116 0.00764286
R25757 VSS.n18758 VSS.n102 0.00764286
R25758 VSS.n18810 VSS.n83 0.00764286
R25759 VSS.n18843 VSS.n66 0.00764286
R25760 VSS.n18839 VSS.n66 0.00764286
R25761 VSS.n18723 VSS.n18722 0.00764286
R25762 VSS.n18723 VSS.n121 0.00764286
R25763 VSS.n18729 VSS.n122 0.00764286
R25764 VSS.n18725 VSS.n118 0.00764286
R25765 VSS.n18744 VSS.n18743 0.00764286
R25766 VSS.n18759 VSS.n101 0.00764286
R25767 VSS.n18781 VSS.n18780 0.00764286
R25768 VSS.n18817 VSS.n79 0.00764286
R25769 VSS.n18842 VSS.n18841 0.00764286
R25770 VSS.n18841 VSS.n18840 0.00764286
R25771 VSS.n306 VSS.n305 0.00764286
R25772 VSS.n315 VSS.n314 0.00764286
R25773 VSS.n390 VSS.n389 0.00764286
R25774 VSS.n421 VSS.n319 0.00764286
R25775 VSS.n18592 VSS.n194 0.00764286
R25776 VSS.n581 VSS.n580 0.00764286
R25777 VSS.n604 VSS.n603 0.00764286
R25778 VSS.n878 VSS.n496 0.00764286
R25779 VSS.n868 VSS.n505 0.00764286
R25780 VSS.n578 VSS.n507 0.00764286
R25781 VSS.n512 VSS.n511 0.00764286
R25782 VSS.n520 VSS.n519 0.00764286
R25783 VSS.n606 VSS.n521 0.00764286
R25784 VSS.n657 VSS.n656 0.00764286
R25785 VSS.n823 VSS.n638 0.00764286
R25786 VSS.n803 VSS.n668 0.00764286
R25787 VSS.n783 VSS.n715 0.00764286
R25788 VSS.n742 VSS.n731 0.00764286
R25789 VSS.n738 VSS.n731 0.00764286
R25790 VSS.n654 VSS.n653 0.00764286
R25791 VSS.n654 VSS.n643 0.00764286
R25792 VSS.n658 VSS.n644 0.00764286
R25793 VSS.n822 VSS.n640 0.00764286
R25794 VSS.n806 VSS.n669 0.00764286
R25795 VSS.n805 VSS.n804 0.00764286
R25796 VSS.n724 VSS.n713 0.00764286
R25797 VSS.n777 VSS.n776 0.00764286
R25798 VSS.n741 VSS.n740 0.00764286
R25799 VSS.n740 VSS.n739 0.00764286
R25800 VSS.n472 VSS.n471 0.00764286
R25801 VSS.n481 VSS.n480 0.00764286
R25802 VSS.n949 VSS.n948 0.00764286
R25803 VSS.n986 VSS.n485 0.00764286
R25804 VSS.n881 VSS.n492 0.00764286
R25805 VSS.n1316 VSS.n1315 0.00764286
R25806 VSS.n17937 VSS.n1297 0.00764286
R25807 VSS.n17917 VSS.n1327 0.00764286
R25808 VSS.n17897 VSS.n1374 0.00764286
R25809 VSS.n1429 VSS.n1390 0.00764286
R25810 VSS.n1430 VSS.n1429 0.00764286
R25811 VSS.n1313 VSS.n1312 0.00764286
R25812 VSS.n1313 VSS.n1302 0.00764286
R25813 VSS.n1317 VSS.n1303 0.00764286
R25814 VSS.n17936 VSS.n1299 0.00764286
R25815 VSS.n17920 VSS.n1328 0.00764286
R25816 VSS.n17919 VSS.n17918 0.00764286
R25817 VSS.n1383 VSS.n1372 0.00764286
R25818 VSS.n17891 VSS.n17890 0.00764286
R25819 VSS.n1428 VSS.n1427 0.00764286
R25820 VSS.n1428 VSS.n1426 0.00764286
R25821 VSS.n1239 VSS.n1236 0.00675
R25822 VSS.n17978 VSS.n17977 0.00675
R25823 VSS.n1266 VSS.n1263 0.00675
R25824 VSS.n1238 VSS.n1237 0.00675
R25825 VSS.n17979 VSS.n1170 0.00675
R25826 VSS.n17967 VSS.n1182 0.00675
R25827 VSS.n1265 VSS.n1264 0.00675
R25828 VSS.n17963 VSS.n1186 0.00675
R25829 VSS.n914 VSS.n909 0.00675
R25830 VSS.n901 VSS.n469 0.00675
R25831 VSS.n991 VSS.n479 0.00675
R25832 VSS.n947 VSS.n946 0.00675
R25833 VSS.n16986 VSS.n16977 0.00675
R25834 VSS.n16980 VSS.n16978 0.00675
R25835 VSS.n17077 VSS.n16958 0.00675
R25836 VSS.n1095 VSS.n1090 0.00675
R25837 VSS.n1082 VSS.n1036 0.00675
R25838 VSS.n18017 VSS.n1046 0.00675
R25839 VSS.n1128 VSS.n1127 0.00675
R25840 VSS.n1038 VSS.n1035 0.00675
R25841 VSS.n18016 VSS.n18015 0.00675
R25842 VSS.n1130 VSS.n1049 0.00675
R25843 VSS.n17141 VSS.n17140 0.00675
R25844 VSS.n17159 VSS.n16909 0.00675
R25845 VSS.n17180 VSS.n16905 0.00675
R25846 VSS.n17182 VSS.n17181 0.00675
R25847 VSS.n17205 VSS.n17203 0.00675
R25848 VSS.n17251 VSS.n16873 0.00675
R25849 VSS.n17139 VSS.n16929 0.00675
R25850 VSS.n17158 VSS.n16908 0.00675
R25851 VSS.n17179 VSS.n17178 0.00675
R25852 VSS.n17206 VSS.n17193 0.00675
R25853 VSS.n17253 VSS.n17252 0.00675
R25854 VSS.n17248 VSS.n16861 0.00675
R25855 VSS.n16984 VSS.n16979 0.00675
R25856 VSS.n17043 VSS.n16981 0.00675
R25857 VSS.n16965 VSS.n16962 0.00675
R25858 VSS.n17076 VSS.n17075 0.00675
R25859 VSS.n17074 VSS.n17070 0.00675
R25860 VSS.n17400 VSS.n17391 0.00675
R25861 VSS.n17394 VSS.n17392 0.00675
R25862 VSS.n17669 VSS.n17372 0.00675
R25863 VSS.n17505 VSS.n17484 0.00675
R25864 VSS.n17476 VSS.n17475 0.00675
R25865 VSS.n17567 VSS.n17446 0.00675
R25866 VSS.n17454 VSS.n17453 0.00675
R25867 VSS.n17541 VSS.n17540 0.00675
R25868 VSS.n17568 VSS.n17444 0.00675
R25869 VSS.n17451 VSS.n17445 0.00675
R25870 VSS.n17733 VSS.n17732 0.00675
R25871 VSS.n17751 VSS.n17323 0.00675
R25872 VSS.n17772 VSS.n17319 0.00675
R25873 VSS.n17774 VSS.n17773 0.00675
R25874 VSS.n17797 VSS.n17795 0.00675
R25875 VSS.n17843 VSS.n17287 0.00675
R25876 VSS.n17731 VSS.n17343 0.00675
R25877 VSS.n17750 VSS.n17322 0.00675
R25878 VSS.n17771 VSS.n17770 0.00675
R25879 VSS.n17798 VSS.n17785 0.00675
R25880 VSS.n17845 VSS.n17844 0.00675
R25881 VSS.n17840 VSS.n17275 0.00675
R25882 VSS.n17398 VSS.n17393 0.00675
R25883 VSS.n17635 VSS.n17395 0.00675
R25884 VSS.n17379 VSS.n17376 0.00675
R25885 VSS.n17668 VSS.n17667 0.00675
R25886 VSS.n17666 VSS.n17662 0.00675
R25887 VSS.n18082 VSS.n276 0.00675
R25888 VSS.n268 VSS.n267 0.00675
R25889 VSS.n18144 VSS.n238 0.00675
R25890 VSS.n246 VSS.n245 0.00675
R25891 VSS.n18256 VSS.n18253 0.00675
R25892 VSS.n18567 VSS.n18566 0.00675
R25893 VSS.n18283 VSS.n18280 0.00675
R25894 VSS.n18255 VSS.n18254 0.00675
R25895 VSS.n18568 VSS.n18187 0.00675
R25896 VSS.n18556 VSS.n18199 0.00675
R25897 VSS.n18282 VSS.n18281 0.00675
R25898 VSS.n18552 VSS.n18203 0.00675
R25899 VSS.n18333 VSS.n18314 0.00675
R25900 VSS.n18513 VSS.n18512 0.00675
R25901 VSS.n18506 VSS.n18345 0.00675
R25902 VSS.n18378 VSS.n18377 0.00675
R25903 VSS.n18409 VSS.n18408 0.00675
R25904 VSS.n18473 VSS.n18472 0.00675
R25905 VSS.n18321 VSS.n18320 0.00675
R25906 VSS.n18514 VSS.n18341 0.00675
R25907 VSS.n18505 VSS.n18347 0.00675
R25908 VSS.n18410 VSS.n18393 0.00675
R25909 VSS.n18471 VSS.n18425 0.00675
R25910 VSS.n18467 VSS.n18431 0.00675
R25911 VSS.n18118 VSS.n18117 0.00675
R25912 VSS.n18145 VSS.n236 0.00675
R25913 VSS.n243 VSS.n237 0.00675
R25914 VSS.n9555 VSS.n9534 0.00675
R25915 VSS.n9526 VSS.n9525 0.00675
R25916 VSS.n9617 VSS.n9496 0.00675
R25917 VSS.n9504 VSS.n9503 0.00675
R25918 VSS.n9450 VSS.n9441 0.00675
R25919 VSS.n9444 VSS.n9442 0.00675
R25920 VSS.n9719 VSS.n9422 0.00675
R25921 VSS.n9448 VSS.n9443 0.00675
R25922 VSS.n9685 VSS.n9445 0.00675
R25923 VSS.n9429 VSS.n9426 0.00675
R25924 VSS.n9718 VSS.n9717 0.00675
R25925 VSS.n9716 VSS.n9712 0.00675
R25926 VSS.n9783 VSS.n9782 0.00675
R25927 VSS.n9801 VSS.n9373 0.00675
R25928 VSS.n9822 VSS.n9369 0.00675
R25929 VSS.n9824 VSS.n9823 0.00675
R25930 VSS.n9847 VSS.n9845 0.00675
R25931 VSS.n9895 VSS.n9894 0.00675
R25932 VSS.n9781 VSS.n9393 0.00675
R25933 VSS.n9800 VSS.n9372 0.00675
R25934 VSS.n9821 VSS.n9820 0.00675
R25935 VSS.n9848 VSS.n9835 0.00675
R25936 VSS.n9896 VSS.n9339 0.00675
R25937 VSS.n9891 VSS.n9326 0.00675
R25938 VSS.n9591 VSS.n9590 0.00675
R25939 VSS.n9618 VSS.n9494 0.00675
R25940 VSS.n9501 VSS.n9495 0.00675
R25941 VSS.n16491 VSS.n16472 0.00675
R25942 VSS.n16526 VSS.n16525 0.00675
R25943 VSS.n16546 VSS.n16545 0.00675
R25944 VSS.n16552 VSS.n16439 0.00675
R25945 VSS.n16392 VSS.n16383 0.00675
R25946 VSS.n16386 VSS.n16384 0.00675
R25947 VSS.n16662 VSS.n16364 0.00675
R25948 VSS.n16390 VSS.n16385 0.00675
R25949 VSS.n16628 VSS.n16387 0.00675
R25950 VSS.n16371 VSS.n16368 0.00675
R25951 VSS.n16661 VSS.n16660 0.00675
R25952 VSS.n16659 VSS.n16655 0.00675
R25953 VSS.n16726 VSS.n16725 0.00675
R25954 VSS.n16744 VSS.n16315 0.00675
R25955 VSS.n16765 VSS.n16311 0.00675
R25956 VSS.n16767 VSS.n16766 0.00675
R25957 VSS.n16790 VSS.n16788 0.00675
R25958 VSS.n16838 VSS.n16837 0.00675
R25959 VSS.n16724 VSS.n16335 0.00675
R25960 VSS.n16743 VSS.n16314 0.00675
R25961 VSS.n16764 VSS.n16763 0.00675
R25962 VSS.n16791 VSS.n16778 0.00675
R25963 VSS.n16839 VSS.n16281 0.00675
R25964 VSS.n16834 VSS.n16268 0.00675
R25965 VSS.n16520 VSS.n16464 0.00675
R25966 VSS.n16547 VSS.n16443 0.00675
R25967 VSS.n16556 VSS.n16440 0.00675
R25968 VSS.n1656 VSS.n1637 0.00675
R25969 VSS.n1691 VSS.n1690 0.00675
R25970 VSS.n1711 VSS.n1710 0.00675
R25971 VSS.n1717 VSS.n1604 0.00675
R25972 VSS.n1564 VSS.n1555 0.00675
R25973 VSS.n1558 VSS.n1556 0.00675
R25974 VSS.n16069 VSS.n1536 0.00675
R25975 VSS.n1562 VSS.n1557 0.00675
R25976 VSS.n16035 VSS.n1559 0.00675
R25977 VSS.n1543 VSS.n1540 0.00675
R25978 VSS.n16068 VSS.n16067 0.00675
R25979 VSS.n16066 VSS.n16062 0.00675
R25980 VSS.n16133 VSS.n16132 0.00675
R25981 VSS.n16151 VSS.n1487 0.00675
R25982 VSS.n16172 VSS.n1483 0.00675
R25983 VSS.n16174 VSS.n16173 0.00675
R25984 VSS.n16197 VSS.n16195 0.00675
R25985 VSS.n16245 VSS.n16244 0.00675
R25986 VSS.n16131 VSS.n1507 0.00675
R25987 VSS.n16150 VSS.n1486 0.00675
R25988 VSS.n16171 VSS.n16170 0.00675
R25989 VSS.n16198 VSS.n16185 0.00675
R25990 VSS.n16246 VSS.n1453 0.00675
R25991 VSS.n16241 VSS.n1440 0.00675
R25992 VSS.n1685 VSS.n1629 0.00675
R25993 VSS.n1712 VSS.n1608 0.00675
R25994 VSS.n1721 VSS.n1605 0.00675
R25995 VSS.n1847 VSS.n1826 0.00675
R25996 VSS.n1818 VSS.n1817 0.00675
R25997 VSS.n1909 VSS.n1788 0.00675
R25998 VSS.n1796 VSS.n1795 0.00675
R25999 VSS.n2021 VSS.n2018 0.00675
R26000 VSS.n2332 VSS.n2331 0.00675
R26001 VSS.n2048 VSS.n2045 0.00675
R26002 VSS.n2020 VSS.n2019 0.00675
R26003 VSS.n2333 VSS.n1952 0.00675
R26004 VSS.n2321 VSS.n1964 0.00675
R26005 VSS.n2047 VSS.n2046 0.00675
R26006 VSS.n2317 VSS.n1968 0.00675
R26007 VSS.n2097 VSS.n2079 0.00675
R26008 VSS.n2275 VSS.n2109 0.00675
R26009 VSS.n2140 VSS.n2134 0.00675
R26010 VSS.n2142 VSS.n2141 0.00675
R26011 VSS.n2253 VSS.n2155 0.00675
R26012 VSS.n2214 VSS.n2212 0.00675
R26013 VSS.n2085 VSS.n2081 0.00675
R26014 VSS.n2274 VSS.n2273 0.00675
R26015 VSS.n2139 VSS.n2138 0.00675
R26016 VSS.n2254 VSS.n2153 0.00675
R26017 VSS.n2215 VSS.n2208 0.00675
R26018 VSS.n2216 VSS.n2202 0.00675
R26019 VSS.n1883 VSS.n1882 0.00675
R26020 VSS.n1910 VSS.n1786 0.00675
R26021 VSS.n1793 VSS.n1787 0.00675
R26022 VSS.n3046 VSS.n3025 0.00675
R26023 VSS.n3017 VSS.n3016 0.00675
R26024 VSS.n3108 VSS.n2987 0.00675
R26025 VSS.n2995 VSS.n2994 0.00675
R26026 VSS.n2941 VSS.n2932 0.00675
R26027 VSS.n2935 VSS.n2933 0.00675
R26028 VSS.n3210 VSS.n2913 0.00675
R26029 VSS.n2939 VSS.n2934 0.00675
R26030 VSS.n3176 VSS.n2936 0.00675
R26031 VSS.n2920 VSS.n2917 0.00675
R26032 VSS.n3209 VSS.n3208 0.00675
R26033 VSS.n3207 VSS.n3203 0.00675
R26034 VSS.n3274 VSS.n3273 0.00675
R26035 VSS.n3292 VSS.n2864 0.00675
R26036 VSS.n3313 VSS.n2860 0.00675
R26037 VSS.n3315 VSS.n3314 0.00675
R26038 VSS.n3338 VSS.n3336 0.00675
R26039 VSS.n3386 VSS.n3385 0.00675
R26040 VSS.n3272 VSS.n2884 0.00675
R26041 VSS.n3291 VSS.n2863 0.00675
R26042 VSS.n3312 VSS.n3311 0.00675
R26043 VSS.n3339 VSS.n3326 0.00675
R26044 VSS.n3387 VSS.n2830 0.00675
R26045 VSS.n3382 VSS.n2817 0.00675
R26046 VSS.n3082 VSS.n3081 0.00675
R26047 VSS.n3109 VSS.n2985 0.00675
R26048 VSS.n2992 VSS.n2986 0.00675
R26049 VSS.n3638 VSS.n3617 0.00675
R26050 VSS.n3609 VSS.n3608 0.00675
R26051 VSS.n3700 VSS.n3579 0.00675
R26052 VSS.n3587 VSS.n3586 0.00675
R26053 VSS.n3533 VSS.n3524 0.00675
R26054 VSS.n3527 VSS.n3525 0.00675
R26055 VSS.n3802 VSS.n3505 0.00675
R26056 VSS.n3531 VSS.n3526 0.00675
R26057 VSS.n3768 VSS.n3528 0.00675
R26058 VSS.n3512 VSS.n3509 0.00675
R26059 VSS.n3801 VSS.n3800 0.00675
R26060 VSS.n3799 VSS.n3795 0.00675
R26061 VSS.n3866 VSS.n3865 0.00675
R26062 VSS.n3884 VSS.n3456 0.00675
R26063 VSS.n3905 VSS.n3452 0.00675
R26064 VSS.n3907 VSS.n3906 0.00675
R26065 VSS.n3930 VSS.n3928 0.00675
R26066 VSS.n3978 VSS.n3977 0.00675
R26067 VSS.n3864 VSS.n3476 0.00675
R26068 VSS.n3883 VSS.n3455 0.00675
R26069 VSS.n3904 VSS.n3903 0.00675
R26070 VSS.n3931 VSS.n3918 0.00675
R26071 VSS.n3979 VSS.n3422 0.00675
R26072 VSS.n3974 VSS.n3409 0.00675
R26073 VSS.n3674 VSS.n3673 0.00675
R26074 VSS.n3701 VSS.n3577 0.00675
R26075 VSS.n3584 VSS.n3578 0.00675
R26076 VSS.n4230 VSS.n4209 0.00675
R26077 VSS.n4201 VSS.n4200 0.00675
R26078 VSS.n4292 VSS.n4171 0.00675
R26079 VSS.n4179 VSS.n4178 0.00675
R26080 VSS.n4125 VSS.n4116 0.00675
R26081 VSS.n4119 VSS.n4117 0.00675
R26082 VSS.n4394 VSS.n4097 0.00675
R26083 VSS.n4123 VSS.n4118 0.00675
R26084 VSS.n4360 VSS.n4120 0.00675
R26085 VSS.n4104 VSS.n4101 0.00675
R26086 VSS.n4393 VSS.n4392 0.00675
R26087 VSS.n4391 VSS.n4387 0.00675
R26088 VSS.n4458 VSS.n4457 0.00675
R26089 VSS.n4476 VSS.n4048 0.00675
R26090 VSS.n4497 VSS.n4044 0.00675
R26091 VSS.n4499 VSS.n4498 0.00675
R26092 VSS.n4522 VSS.n4520 0.00675
R26093 VSS.n4570 VSS.n4569 0.00675
R26094 VSS.n4456 VSS.n4068 0.00675
R26095 VSS.n4475 VSS.n4047 0.00675
R26096 VSS.n4496 VSS.n4495 0.00675
R26097 VSS.n4523 VSS.n4510 0.00675
R26098 VSS.n4571 VSS.n4014 0.00675
R26099 VSS.n4566 VSS.n4001 0.00675
R26100 VSS.n4266 VSS.n4265 0.00675
R26101 VSS.n4293 VSS.n4169 0.00675
R26102 VSS.n4176 VSS.n4170 0.00675
R26103 VSS.n4822 VSS.n4801 0.00675
R26104 VSS.n4793 VSS.n4792 0.00675
R26105 VSS.n4884 VSS.n4763 0.00675
R26106 VSS.n4771 VSS.n4770 0.00675
R26107 VSS.n4717 VSS.n4708 0.00675
R26108 VSS.n4711 VSS.n4709 0.00675
R26109 VSS.n4986 VSS.n4689 0.00675
R26110 VSS.n4715 VSS.n4710 0.00675
R26111 VSS.n4952 VSS.n4712 0.00675
R26112 VSS.n4696 VSS.n4693 0.00675
R26113 VSS.n4985 VSS.n4984 0.00675
R26114 VSS.n4983 VSS.n4979 0.00675
R26115 VSS.n5050 VSS.n5049 0.00675
R26116 VSS.n5068 VSS.n4640 0.00675
R26117 VSS.n5089 VSS.n4636 0.00675
R26118 VSS.n5091 VSS.n5090 0.00675
R26119 VSS.n5114 VSS.n5112 0.00675
R26120 VSS.n5162 VSS.n5161 0.00675
R26121 VSS.n5048 VSS.n4660 0.00675
R26122 VSS.n5067 VSS.n4639 0.00675
R26123 VSS.n5088 VSS.n5087 0.00675
R26124 VSS.n5115 VSS.n5102 0.00675
R26125 VSS.n5163 VSS.n4606 0.00675
R26126 VSS.n5158 VSS.n4593 0.00675
R26127 VSS.n4858 VSS.n4857 0.00675
R26128 VSS.n4885 VSS.n4761 0.00675
R26129 VSS.n4768 VSS.n4762 0.00675
R26130 VSS.n2443 VSS.n2422 0.00675
R26131 VSS.n2414 VSS.n2413 0.00675
R26132 VSS.n2505 VSS.n2384 0.00675
R26133 VSS.n2392 VSS.n2391 0.00675
R26134 VSS.n2617 VSS.n2614 0.00675
R26135 VSS.n5297 VSS.n5296 0.00675
R26136 VSS.n2644 VSS.n2641 0.00675
R26137 VSS.n2616 VSS.n2615 0.00675
R26138 VSS.n5298 VSS.n2548 0.00675
R26139 VSS.n5286 VSS.n2560 0.00675
R26140 VSS.n2643 VSS.n2642 0.00675
R26141 VSS.n5282 VSS.n2564 0.00675
R26142 VSS.n2693 VSS.n2675 0.00675
R26143 VSS.n5240 VSS.n2705 0.00675
R26144 VSS.n2736 VSS.n2730 0.00675
R26145 VSS.n2738 VSS.n2737 0.00675
R26146 VSS.n5218 VSS.n2751 0.00675
R26147 VSS.n2810 VSS.n2808 0.00675
R26148 VSS.n2681 VSS.n2677 0.00675
R26149 VSS.n5239 VSS.n5238 0.00675
R26150 VSS.n2735 VSS.n2734 0.00675
R26151 VSS.n5219 VSS.n2749 0.00675
R26152 VSS.n2811 VSS.n2804 0.00675
R26153 VSS.n2812 VSS.n2798 0.00675
R26154 VSS.n2479 VSS.n2478 0.00675
R26155 VSS.n2506 VSS.n2382 0.00675
R26156 VSS.n2389 VSS.n2383 0.00675
R26157 VSS.n5404 VSS.n5383 0.00675
R26158 VSS.n5375 VSS.n5374 0.00675
R26159 VSS.n5466 VSS.n5345 0.00675
R26160 VSS.n5353 VSS.n5352 0.00675
R26161 VSS.n5578 VSS.n5575 0.00675
R26162 VSS.n5870 VSS.n5869 0.00675
R26163 VSS.n5605 VSS.n5602 0.00675
R26164 VSS.n5577 VSS.n5576 0.00675
R26165 VSS.n5871 VSS.n5509 0.00675
R26166 VSS.n5859 VSS.n5521 0.00675
R26167 VSS.n5604 VSS.n5603 0.00675
R26168 VSS.n5855 VSS.n5525 0.00675
R26169 VSS.n5654 VSS.n5636 0.00675
R26170 VSS.n5813 VSS.n5666 0.00675
R26171 VSS.n5697 VSS.n5691 0.00675
R26172 VSS.n5699 VSS.n5698 0.00675
R26173 VSS.n5791 VSS.n5712 0.00675
R26174 VSS.n5737 VSS.n5736 0.00675
R26175 VSS.n5642 VSS.n5638 0.00675
R26176 VSS.n5812 VSS.n5811 0.00675
R26177 VSS.n5696 VSS.n5695 0.00675
R26178 VSS.n5792 VSS.n5710 0.00675
R26179 VSS.n5738 VSS.n5730 0.00675
R26180 VSS.n5733 VSS.n2 0.00675
R26181 VSS.n5440 VSS.n5439 0.00675
R26182 VSS.n5467 VSS.n5343 0.00675
R26183 VSS.n5350 VSS.n5344 0.00675
R26184 VSS.n5977 VSS.n5956 0.00675
R26185 VSS.n5948 VSS.n5947 0.00675
R26186 VSS.n6039 VSS.n5918 0.00675
R26187 VSS.n5926 VSS.n5925 0.00675
R26188 VSS.n6151 VSS.n6148 0.00675
R26189 VSS.n6462 VSS.n6461 0.00675
R26190 VSS.n6178 VSS.n6175 0.00675
R26191 VSS.n6150 VSS.n6149 0.00675
R26192 VSS.n6463 VSS.n6082 0.00675
R26193 VSS.n6451 VSS.n6094 0.00675
R26194 VSS.n6177 VSS.n6176 0.00675
R26195 VSS.n6447 VSS.n6098 0.00675
R26196 VSS.n6227 VSS.n6209 0.00675
R26197 VSS.n6405 VSS.n6239 0.00675
R26198 VSS.n6270 VSS.n6264 0.00675
R26199 VSS.n6272 VSS.n6271 0.00675
R26200 VSS.n6383 VSS.n6285 0.00675
R26201 VSS.n6344 VSS.n6342 0.00675
R26202 VSS.n6215 VSS.n6211 0.00675
R26203 VSS.n6404 VSS.n6403 0.00675
R26204 VSS.n6269 VSS.n6268 0.00675
R26205 VSS.n6384 VSS.n6283 0.00675
R26206 VSS.n6345 VSS.n6338 0.00675
R26207 VSS.n6346 VSS.n6332 0.00675
R26208 VSS.n6013 VSS.n6012 0.00675
R26209 VSS.n6040 VSS.n5916 0.00675
R26210 VSS.n5923 VSS.n5917 0.00675
R26211 VSS.n7779 VSS.n7758 0.00675
R26212 VSS.n7750 VSS.n7749 0.00675
R26213 VSS.n7841 VSS.n7720 0.00675
R26214 VSS.n7728 VSS.n7727 0.00675
R26215 VSS.n7674 VSS.n7665 0.00675
R26216 VSS.n7668 VSS.n7666 0.00675
R26217 VSS.n7943 VSS.n7646 0.00675
R26218 VSS.n7672 VSS.n7667 0.00675
R26219 VSS.n7909 VSS.n7669 0.00675
R26220 VSS.n7653 VSS.n7650 0.00675
R26221 VSS.n7942 VSS.n7941 0.00675
R26222 VSS.n7940 VSS.n7936 0.00675
R26223 VSS.n8007 VSS.n8006 0.00675
R26224 VSS.n8025 VSS.n7597 0.00675
R26225 VSS.n8046 VSS.n7593 0.00675
R26226 VSS.n8048 VSS.n8047 0.00675
R26227 VSS.n8071 VSS.n8069 0.00675
R26228 VSS.n8119 VSS.n8118 0.00675
R26229 VSS.n8005 VSS.n7617 0.00675
R26230 VSS.n8024 VSS.n7596 0.00675
R26231 VSS.n8045 VSS.n8044 0.00675
R26232 VSS.n8072 VSS.n8059 0.00675
R26233 VSS.n8120 VSS.n7563 0.00675
R26234 VSS.n8115 VSS.n7550 0.00675
R26235 VSS.n7815 VSS.n7814 0.00675
R26236 VSS.n7842 VSS.n7718 0.00675
R26237 VSS.n7725 VSS.n7719 0.00675
R26238 VSS.n8371 VSS.n8350 0.00675
R26239 VSS.n8342 VSS.n8341 0.00675
R26240 VSS.n8433 VSS.n8312 0.00675
R26241 VSS.n8320 VSS.n8319 0.00675
R26242 VSS.n8266 VSS.n8257 0.00675
R26243 VSS.n8260 VSS.n8258 0.00675
R26244 VSS.n8535 VSS.n8238 0.00675
R26245 VSS.n8264 VSS.n8259 0.00675
R26246 VSS.n8501 VSS.n8261 0.00675
R26247 VSS.n8245 VSS.n8242 0.00675
R26248 VSS.n8534 VSS.n8533 0.00675
R26249 VSS.n8532 VSS.n8528 0.00675
R26250 VSS.n8599 VSS.n8598 0.00675
R26251 VSS.n8617 VSS.n8189 0.00675
R26252 VSS.n8638 VSS.n8185 0.00675
R26253 VSS.n8640 VSS.n8639 0.00675
R26254 VSS.n8663 VSS.n8661 0.00675
R26255 VSS.n8711 VSS.n8710 0.00675
R26256 VSS.n8597 VSS.n8209 0.00675
R26257 VSS.n8616 VSS.n8188 0.00675
R26258 VSS.n8637 VSS.n8636 0.00675
R26259 VSS.n8664 VSS.n8651 0.00675
R26260 VSS.n8712 VSS.n8155 0.00675
R26261 VSS.n8707 VSS.n8142 0.00675
R26262 VSS.n8407 VSS.n8406 0.00675
R26263 VSS.n8434 VSS.n8310 0.00675
R26264 VSS.n8317 VSS.n8311 0.00675
R26265 VSS.n8963 VSS.n8942 0.00675
R26266 VSS.n8934 VSS.n8933 0.00675
R26267 VSS.n9025 VSS.n8904 0.00675
R26268 VSS.n8912 VSS.n8911 0.00675
R26269 VSS.n8858 VSS.n8849 0.00675
R26270 VSS.n8852 VSS.n8850 0.00675
R26271 VSS.n9127 VSS.n8830 0.00675
R26272 VSS.n8856 VSS.n8851 0.00675
R26273 VSS.n9093 VSS.n8853 0.00675
R26274 VSS.n8837 VSS.n8834 0.00675
R26275 VSS.n9126 VSS.n9125 0.00675
R26276 VSS.n9124 VSS.n9120 0.00675
R26277 VSS.n9191 VSS.n9190 0.00675
R26278 VSS.n9209 VSS.n8781 0.00675
R26279 VSS.n9230 VSS.n8777 0.00675
R26280 VSS.n9232 VSS.n9231 0.00675
R26281 VSS.n9255 VSS.n9253 0.00675
R26282 VSS.n9303 VSS.n9302 0.00675
R26283 VSS.n9189 VSS.n8801 0.00675
R26284 VSS.n9208 VSS.n8780 0.00675
R26285 VSS.n9229 VSS.n9228 0.00675
R26286 VSS.n9256 VSS.n9243 0.00675
R26287 VSS.n9304 VSS.n8747 0.00675
R26288 VSS.n9299 VSS.n8734 0.00675
R26289 VSS.n8999 VSS.n8998 0.00675
R26290 VSS.n9026 VSS.n8902 0.00675
R26291 VSS.n8909 VSS.n8903 0.00675
R26292 VSS.n10147 VSS.n10126 0.00675
R26293 VSS.n10118 VSS.n10117 0.00675
R26294 VSS.n10209 VSS.n10088 0.00675
R26295 VSS.n10096 VSS.n10095 0.00675
R26296 VSS.n10042 VSS.n10033 0.00675
R26297 VSS.n10036 VSS.n10034 0.00675
R26298 VSS.n10311 VSS.n10014 0.00675
R26299 VSS.n10040 VSS.n10035 0.00675
R26300 VSS.n10277 VSS.n10037 0.00675
R26301 VSS.n10021 VSS.n10018 0.00675
R26302 VSS.n10310 VSS.n10309 0.00675
R26303 VSS.n10308 VSS.n10304 0.00675
R26304 VSS.n10375 VSS.n10374 0.00675
R26305 VSS.n10393 VSS.n9965 0.00675
R26306 VSS.n10414 VSS.n9961 0.00675
R26307 VSS.n10416 VSS.n10415 0.00675
R26308 VSS.n10439 VSS.n10437 0.00675
R26309 VSS.n10487 VSS.n10486 0.00675
R26310 VSS.n10373 VSS.n9985 0.00675
R26311 VSS.n10392 VSS.n9964 0.00675
R26312 VSS.n10413 VSS.n10412 0.00675
R26313 VSS.n10440 VSS.n10427 0.00675
R26314 VSS.n10488 VSS.n9931 0.00675
R26315 VSS.n10483 VSS.n9918 0.00675
R26316 VSS.n10183 VSS.n10182 0.00675
R26317 VSS.n10210 VSS.n10086 0.00675
R26318 VSS.n10093 VSS.n10087 0.00675
R26319 VSS.n10739 VSS.n10718 0.00675
R26320 VSS.n10710 VSS.n10709 0.00675
R26321 VSS.n10801 VSS.n10680 0.00675
R26322 VSS.n10688 VSS.n10687 0.00675
R26323 VSS.n10634 VSS.n10625 0.00675
R26324 VSS.n10628 VSS.n10626 0.00675
R26325 VSS.n10903 VSS.n10606 0.00675
R26326 VSS.n10632 VSS.n10627 0.00675
R26327 VSS.n10869 VSS.n10629 0.00675
R26328 VSS.n10613 VSS.n10610 0.00675
R26329 VSS.n10902 VSS.n10901 0.00675
R26330 VSS.n10900 VSS.n10896 0.00675
R26331 VSS.n10967 VSS.n10966 0.00675
R26332 VSS.n10985 VSS.n10557 0.00675
R26333 VSS.n11006 VSS.n10553 0.00675
R26334 VSS.n11008 VSS.n11007 0.00675
R26335 VSS.n11031 VSS.n11029 0.00675
R26336 VSS.n11079 VSS.n11078 0.00675
R26337 VSS.n10965 VSS.n10577 0.00675
R26338 VSS.n10984 VSS.n10556 0.00675
R26339 VSS.n11005 VSS.n11004 0.00675
R26340 VSS.n11032 VSS.n11019 0.00675
R26341 VSS.n11080 VSS.n10523 0.00675
R26342 VSS.n11075 VSS.n10510 0.00675
R26343 VSS.n10775 VSS.n10774 0.00675
R26344 VSS.n10802 VSS.n10678 0.00675
R26345 VSS.n10685 VSS.n10679 0.00675
R26346 VSS.n11331 VSS.n11310 0.00675
R26347 VSS.n11302 VSS.n11301 0.00675
R26348 VSS.n11393 VSS.n11272 0.00675
R26349 VSS.n11280 VSS.n11279 0.00675
R26350 VSS.n11226 VSS.n11217 0.00675
R26351 VSS.n11220 VSS.n11218 0.00675
R26352 VSS.n11495 VSS.n11198 0.00675
R26353 VSS.n11224 VSS.n11219 0.00675
R26354 VSS.n11461 VSS.n11221 0.00675
R26355 VSS.n11205 VSS.n11202 0.00675
R26356 VSS.n11494 VSS.n11493 0.00675
R26357 VSS.n11492 VSS.n11488 0.00675
R26358 VSS.n11559 VSS.n11558 0.00675
R26359 VSS.n11577 VSS.n11149 0.00675
R26360 VSS.n11598 VSS.n11145 0.00675
R26361 VSS.n11600 VSS.n11599 0.00675
R26362 VSS.n11623 VSS.n11621 0.00675
R26363 VSS.n11671 VSS.n11670 0.00675
R26364 VSS.n11557 VSS.n11169 0.00675
R26365 VSS.n11576 VSS.n11148 0.00675
R26366 VSS.n11597 VSS.n11596 0.00675
R26367 VSS.n11624 VSS.n11611 0.00675
R26368 VSS.n11672 VSS.n11115 0.00675
R26369 VSS.n11667 VSS.n11102 0.00675
R26370 VSS.n11367 VSS.n11366 0.00675
R26371 VSS.n11394 VSS.n11270 0.00675
R26372 VSS.n11277 VSS.n11271 0.00675
R26373 VSS.n11923 VSS.n11902 0.00675
R26374 VSS.n11894 VSS.n11893 0.00675
R26375 VSS.n11985 VSS.n11864 0.00675
R26376 VSS.n11872 VSS.n11871 0.00675
R26377 VSS.n11818 VSS.n11809 0.00675
R26378 VSS.n11812 VSS.n11810 0.00675
R26379 VSS.n12087 VSS.n11790 0.00675
R26380 VSS.n11816 VSS.n11811 0.00675
R26381 VSS.n12053 VSS.n11813 0.00675
R26382 VSS.n11797 VSS.n11794 0.00675
R26383 VSS.n12086 VSS.n12085 0.00675
R26384 VSS.n12084 VSS.n12080 0.00675
R26385 VSS.n12151 VSS.n12150 0.00675
R26386 VSS.n12169 VSS.n11741 0.00675
R26387 VSS.n12190 VSS.n11737 0.00675
R26388 VSS.n12192 VSS.n12191 0.00675
R26389 VSS.n12215 VSS.n12213 0.00675
R26390 VSS.n12263 VSS.n12262 0.00675
R26391 VSS.n12149 VSS.n11761 0.00675
R26392 VSS.n12168 VSS.n11740 0.00675
R26393 VSS.n12189 VSS.n12188 0.00675
R26394 VSS.n12216 VSS.n12203 0.00675
R26395 VSS.n12264 VSS.n11707 0.00675
R26396 VSS.n12259 VSS.n11694 0.00675
R26397 VSS.n11959 VSS.n11958 0.00675
R26398 VSS.n11986 VSS.n11862 0.00675
R26399 VSS.n11869 VSS.n11863 0.00675
R26400 VSS.n12515 VSS.n12494 0.00675
R26401 VSS.n12486 VSS.n12485 0.00675
R26402 VSS.n12577 VSS.n12456 0.00675
R26403 VSS.n12464 VSS.n12463 0.00675
R26404 VSS.n12410 VSS.n12401 0.00675
R26405 VSS.n12404 VSS.n12402 0.00675
R26406 VSS.n12679 VSS.n12382 0.00675
R26407 VSS.n12408 VSS.n12403 0.00675
R26408 VSS.n12645 VSS.n12405 0.00675
R26409 VSS.n12389 VSS.n12386 0.00675
R26410 VSS.n12678 VSS.n12677 0.00675
R26411 VSS.n12676 VSS.n12672 0.00675
R26412 VSS.n12743 VSS.n12742 0.00675
R26413 VSS.n12761 VSS.n12333 0.00675
R26414 VSS.n12782 VSS.n12329 0.00675
R26415 VSS.n12784 VSS.n12783 0.00675
R26416 VSS.n12807 VSS.n12805 0.00675
R26417 VSS.n12855 VSS.n12854 0.00675
R26418 VSS.n12741 VSS.n12353 0.00675
R26419 VSS.n12760 VSS.n12332 0.00675
R26420 VSS.n12781 VSS.n12780 0.00675
R26421 VSS.n12808 VSS.n12795 0.00675
R26422 VSS.n12856 VSS.n12299 0.00675
R26423 VSS.n12851 VSS.n12286 0.00675
R26424 VSS.n12551 VSS.n12550 0.00675
R26425 VSS.n12578 VSS.n12454 0.00675
R26426 VSS.n12461 VSS.n12455 0.00675
R26427 VSS.n13107 VSS.n13086 0.00675
R26428 VSS.n13078 VSS.n13077 0.00675
R26429 VSS.n13169 VSS.n13048 0.00675
R26430 VSS.n13056 VSS.n13055 0.00675
R26431 VSS.n13002 VSS.n12993 0.00675
R26432 VSS.n12996 VSS.n12994 0.00675
R26433 VSS.n13271 VSS.n12974 0.00675
R26434 VSS.n13000 VSS.n12995 0.00675
R26435 VSS.n13237 VSS.n12997 0.00675
R26436 VSS.n12981 VSS.n12978 0.00675
R26437 VSS.n13270 VSS.n13269 0.00675
R26438 VSS.n13268 VSS.n13264 0.00675
R26439 VSS.n13335 VSS.n13334 0.00675
R26440 VSS.n13353 VSS.n12925 0.00675
R26441 VSS.n13374 VSS.n12921 0.00675
R26442 VSS.n13376 VSS.n13375 0.00675
R26443 VSS.n13399 VSS.n13397 0.00675
R26444 VSS.n13447 VSS.n13446 0.00675
R26445 VSS.n13333 VSS.n12945 0.00675
R26446 VSS.n13352 VSS.n12924 0.00675
R26447 VSS.n13373 VSS.n13372 0.00675
R26448 VSS.n13400 VSS.n13387 0.00675
R26449 VSS.n13448 VSS.n12891 0.00675
R26450 VSS.n13443 VSS.n12878 0.00675
R26451 VSS.n13143 VSS.n13142 0.00675
R26452 VSS.n13170 VSS.n13046 0.00675
R26453 VSS.n13053 VSS.n13047 0.00675
R26454 VSS.n13699 VSS.n13678 0.00675
R26455 VSS.n13670 VSS.n13669 0.00675
R26456 VSS.n13761 VSS.n13640 0.00675
R26457 VSS.n13648 VSS.n13647 0.00675
R26458 VSS.n13594 VSS.n13585 0.00675
R26459 VSS.n13588 VSS.n13586 0.00675
R26460 VSS.n13863 VSS.n13566 0.00675
R26461 VSS.n13592 VSS.n13587 0.00675
R26462 VSS.n13829 VSS.n13589 0.00675
R26463 VSS.n13573 VSS.n13570 0.00675
R26464 VSS.n13862 VSS.n13861 0.00675
R26465 VSS.n13860 VSS.n13856 0.00675
R26466 VSS.n13927 VSS.n13926 0.00675
R26467 VSS.n13945 VSS.n13517 0.00675
R26468 VSS.n13966 VSS.n13513 0.00675
R26469 VSS.n13968 VSS.n13967 0.00675
R26470 VSS.n13991 VSS.n13989 0.00675
R26471 VSS.n14039 VSS.n14038 0.00675
R26472 VSS.n13925 VSS.n13537 0.00675
R26473 VSS.n13944 VSS.n13516 0.00675
R26474 VSS.n13965 VSS.n13964 0.00675
R26475 VSS.n13992 VSS.n13979 0.00675
R26476 VSS.n14040 VSS.n13483 0.00675
R26477 VSS.n14035 VSS.n13470 0.00675
R26478 VSS.n13735 VSS.n13734 0.00675
R26479 VSS.n13762 VSS.n13638 0.00675
R26480 VSS.n13645 VSS.n13639 0.00675
R26481 VSS.n14291 VSS.n14270 0.00675
R26482 VSS.n14262 VSS.n14261 0.00675
R26483 VSS.n14353 VSS.n14232 0.00675
R26484 VSS.n14240 VSS.n14239 0.00675
R26485 VSS.n14186 VSS.n14177 0.00675
R26486 VSS.n14180 VSS.n14178 0.00675
R26487 VSS.n14455 VSS.n14158 0.00675
R26488 VSS.n14184 VSS.n14179 0.00675
R26489 VSS.n14421 VSS.n14181 0.00675
R26490 VSS.n14165 VSS.n14162 0.00675
R26491 VSS.n14454 VSS.n14453 0.00675
R26492 VSS.n14452 VSS.n14448 0.00675
R26493 VSS.n14519 VSS.n14518 0.00675
R26494 VSS.n14537 VSS.n14109 0.00675
R26495 VSS.n14558 VSS.n14105 0.00675
R26496 VSS.n14560 VSS.n14559 0.00675
R26497 VSS.n14583 VSS.n14581 0.00675
R26498 VSS.n14631 VSS.n14630 0.00675
R26499 VSS.n14517 VSS.n14129 0.00675
R26500 VSS.n14536 VSS.n14108 0.00675
R26501 VSS.n14557 VSS.n14556 0.00675
R26502 VSS.n14584 VSS.n14571 0.00675
R26503 VSS.n14632 VSS.n14075 0.00675
R26504 VSS.n14627 VSS.n14062 0.00675
R26505 VSS.n14327 VSS.n14326 0.00675
R26506 VSS.n14354 VSS.n14230 0.00675
R26507 VSS.n14237 VSS.n14231 0.00675
R26508 VSS.n14883 VSS.n14862 0.00675
R26509 VSS.n14854 VSS.n14853 0.00675
R26510 VSS.n14945 VSS.n14824 0.00675
R26511 VSS.n14832 VSS.n14831 0.00675
R26512 VSS.n14778 VSS.n14769 0.00675
R26513 VSS.n14772 VSS.n14770 0.00675
R26514 VSS.n15047 VSS.n14750 0.00675
R26515 VSS.n14776 VSS.n14771 0.00675
R26516 VSS.n15013 VSS.n14773 0.00675
R26517 VSS.n14757 VSS.n14754 0.00675
R26518 VSS.n15046 VSS.n15045 0.00675
R26519 VSS.n15044 VSS.n15040 0.00675
R26520 VSS.n15111 VSS.n15110 0.00675
R26521 VSS.n15129 VSS.n14701 0.00675
R26522 VSS.n15150 VSS.n14697 0.00675
R26523 VSS.n15152 VSS.n15151 0.00675
R26524 VSS.n15175 VSS.n15173 0.00675
R26525 VSS.n15223 VSS.n15222 0.00675
R26526 VSS.n15109 VSS.n14721 0.00675
R26527 VSS.n15128 VSS.n14700 0.00675
R26528 VSS.n15149 VSS.n15148 0.00675
R26529 VSS.n15176 VSS.n15163 0.00675
R26530 VSS.n15224 VSS.n14667 0.00675
R26531 VSS.n15219 VSS.n14654 0.00675
R26532 VSS.n14919 VSS.n14918 0.00675
R26533 VSS.n14946 VSS.n14822 0.00675
R26534 VSS.n14829 VSS.n14823 0.00675
R26535 VSS.n15475 VSS.n15454 0.00675
R26536 VSS.n15446 VSS.n15445 0.00675
R26537 VSS.n15537 VSS.n15416 0.00675
R26538 VSS.n15424 VSS.n15423 0.00675
R26539 VSS.n15370 VSS.n15361 0.00675
R26540 VSS.n15364 VSS.n15362 0.00675
R26541 VSS.n15639 VSS.n15342 0.00675
R26542 VSS.n15368 VSS.n15363 0.00675
R26543 VSS.n15605 VSS.n15365 0.00675
R26544 VSS.n15349 VSS.n15346 0.00675
R26545 VSS.n15638 VSS.n15637 0.00675
R26546 VSS.n15636 VSS.n15632 0.00675
R26547 VSS.n15703 VSS.n15702 0.00675
R26548 VSS.n15721 VSS.n15293 0.00675
R26549 VSS.n15742 VSS.n15289 0.00675
R26550 VSS.n15744 VSS.n15743 0.00675
R26551 VSS.n15767 VSS.n15765 0.00675
R26552 VSS.n15815 VSS.n15814 0.00675
R26553 VSS.n15701 VSS.n15313 0.00675
R26554 VSS.n15720 VSS.n15292 0.00675
R26555 VSS.n15741 VSS.n15740 0.00675
R26556 VSS.n15768 VSS.n15755 0.00675
R26557 VSS.n15816 VSS.n15259 0.00675
R26558 VSS.n15811 VSS.n15246 0.00675
R26559 VSS.n15511 VSS.n15510 0.00675
R26560 VSS.n15538 VSS.n15414 0.00675
R26561 VSS.n15421 VSS.n15415 0.00675
R26562 VSS.n6583 VSS.n6562 0.00675
R26563 VSS.n6554 VSS.n6553 0.00675
R26564 VSS.n6645 VSS.n6524 0.00675
R26565 VSS.n6532 VSS.n6531 0.00675
R26566 VSS.n6757 VSS.n6754 0.00675
R26567 VSS.n15950 VSS.n15949 0.00675
R26568 VSS.n6784 VSS.n6781 0.00675
R26569 VSS.n6756 VSS.n6755 0.00675
R26570 VSS.n15951 VSS.n6688 0.00675
R26571 VSS.n15939 VSS.n6700 0.00675
R26572 VSS.n6783 VSS.n6782 0.00675
R26573 VSS.n15935 VSS.n6704 0.00675
R26574 VSS.n6833 VSS.n6815 0.00675
R26575 VSS.n15893 VSS.n6845 0.00675
R26576 VSS.n6876 VSS.n6870 0.00675
R26577 VSS.n6878 VSS.n6877 0.00675
R26578 VSS.n15871 VSS.n6891 0.00675
R26579 VSS.n6950 VSS.n6948 0.00675
R26580 VSS.n6821 VSS.n6817 0.00675
R26581 VSS.n15892 VSS.n15891 0.00675
R26582 VSS.n6875 VSS.n6874 0.00675
R26583 VSS.n15872 VSS.n6889 0.00675
R26584 VSS.n6951 VSS.n6944 0.00675
R26585 VSS.n6952 VSS.n6938 0.00675
R26586 VSS.n6619 VSS.n6618 0.00675
R26587 VSS.n6646 VSS.n6522 0.00675
R26588 VSS.n6529 VSS.n6523 0.00675
R26589 VSS.n7180 VSS.n7161 0.00675
R26590 VSS.n7215 VSS.n7214 0.00675
R26591 VSS.n7235 VSS.n7234 0.00675
R26592 VSS.n7241 VSS.n7128 0.00675
R26593 VSS.n7081 VSS.n7072 0.00675
R26594 VSS.n7075 VSS.n7073 0.00675
R26595 VSS.n7351 VSS.n7053 0.00675
R26596 VSS.n7079 VSS.n7074 0.00675
R26597 VSS.n7317 VSS.n7076 0.00675
R26598 VSS.n7060 VSS.n7057 0.00675
R26599 VSS.n7350 VSS.n7349 0.00675
R26600 VSS.n7348 VSS.n7344 0.00675
R26601 VSS.n7415 VSS.n7414 0.00675
R26602 VSS.n7433 VSS.n7004 0.00675
R26603 VSS.n7454 VSS.n7000 0.00675
R26604 VSS.n7456 VSS.n7455 0.00675
R26605 VSS.n7479 VSS.n7477 0.00675
R26606 VSS.n7527 VSS.n7526 0.00675
R26607 VSS.n7413 VSS.n7024 0.00675
R26608 VSS.n7432 VSS.n7003 0.00675
R26609 VSS.n7453 VSS.n7452 0.00675
R26610 VSS.n7480 VSS.n7467 0.00675
R26611 VSS.n7528 VSS.n6970 0.00675
R26612 VSS.n7523 VSS.n6957 0.00675
R26613 VSS.n7209 VSS.n7153 0.00675
R26614 VSS.n7236 VSS.n7132 0.00675
R26615 VSS.n7245 VSS.n7129 0.00675
R26616 VSS.n355 VSS.n354 0.00675
R26617 VSS.n370 VSS.n303 0.00675
R26618 VSS.n426 VSS.n313 0.00675
R26619 VSS.n392 VSS.n391 0.00675
R26620 VSS.n179 VSS.n170 0.00675
R26621 VSS.n173 VSS.n171 0.00675
R26622 VSS.n18663 VSS.n151 0.00675
R26623 VSS.n177 VSS.n172 0.00675
R26624 VSS.n18629 VSS.n174 0.00675
R26625 VSS.n158 VSS.n155 0.00675
R26626 VSS.n18662 VSS.n18661 0.00675
R26627 VSS.n18660 VSS.n18656 0.00675
R26628 VSS.n18727 VSS.n18726 0.00675
R26629 VSS.n18745 VSS.n102 0.00675
R26630 VSS.n18766 VSS.n98 0.00675
R26631 VSS.n18768 VSS.n18767 0.00675
R26632 VSS.n18791 VSS.n18789 0.00675
R26633 VSS.n18839 VSS.n18838 0.00675
R26634 VSS.n18725 VSS.n122 0.00675
R26635 VSS.n18744 VSS.n101 0.00675
R26636 VSS.n18765 VSS.n18764 0.00675
R26637 VSS.n18792 VSS.n18779 0.00675
R26638 VSS.n18840 VSS.n68 0.00675
R26639 VSS.n18835 VSS.n55 0.00675
R26640 VSS.n305 VSS.n302 0.00675
R26641 VSS.n425 VSS.n424 0.00675
R26642 VSS.n389 VSS.n316 0.00675
R26643 VSS.n580 VSS.n577 0.00675
R26644 VSS.n864 VSS.n863 0.00675
R26645 VSS.n607 VSS.n604 0.00675
R26646 VSS.n579 VSS.n578 0.00675
R26647 VSS.n865 VSS.n508 0.00675
R26648 VSS.n853 VSS.n520 0.00675
R26649 VSS.n606 VSS.n605 0.00675
R26650 VSS.n849 VSS.n524 0.00675
R26651 VSS.n656 VSS.n638 0.00675
R26652 VSS.n807 VSS.n668 0.00675
R26653 VSS.n699 VSS.n693 0.00675
R26654 VSS.n701 VSS.n700 0.00675
R26655 VSS.n785 VSS.n714 0.00675
R26656 VSS.n738 VSS.n737 0.00675
R26657 VSS.n644 VSS.n640 0.00675
R26658 VSS.n806 VSS.n805 0.00675
R26659 VSS.n698 VSS.n697 0.00675
R26660 VSS.n786 VSS.n712 0.00675
R26661 VSS.n739 VSS.n735 0.00675
R26662 VSS.n732 VSS.n51 0.00675
R26663 VSS.n471 VSS.n468 0.00675
R26664 VSS.n990 VSS.n989 0.00675
R26665 VSS.n949 VSS.n482 0.00675
R26666 VSS.n1315 VSS.n1297 0.00675
R26667 VSS.n17921 VSS.n1327 0.00675
R26668 VSS.n1358 VSS.n1352 0.00675
R26669 VSS.n1360 VSS.n1359 0.00675
R26670 VSS.n17899 VSS.n1373 0.00675
R26671 VSS.n1432 VSS.n1430 0.00675
R26672 VSS.n1303 VSS.n1299 0.00675
R26673 VSS.n17920 VSS.n17919 0.00675
R26674 VSS.n1357 VSS.n1356 0.00675
R26675 VSS.n17900 VSS.n1371 0.00675
R26676 VSS.n1433 VSS.n1426 0.00675
R26677 VSS.n1434 VSS.n1420 0.00675
R26678 VSS.n17110 VSS.n17109 0.00636816
R26679 VSS.n17702 VSS.n17701 0.00636816
R26680 VSS.n18324 VSS.n18308 0.00636816
R26681 VSS.n9752 VSS.n9751 0.00636816
R26682 VSS.n16695 VSS.n16694 0.00636816
R26683 VSS.n16102 VSS.n16101 0.00636816
R26684 VSS.n2088 VSS.n2073 0.00636816
R26685 VSS.n3243 VSS.n3242 0.00636816
R26686 VSS.n3835 VSS.n3834 0.00636816
R26687 VSS.n4427 VSS.n4426 0.00636816
R26688 VSS.n5019 VSS.n5018 0.00636816
R26689 VSS.n2684 VSS.n2669 0.00636816
R26690 VSS.n5645 VSS.n5630 0.00636816
R26691 VSS.n6218 VSS.n6203 0.00636816
R26692 VSS.n7976 VSS.n7975 0.00636816
R26693 VSS.n8568 VSS.n8567 0.00636816
R26694 VSS.n9160 VSS.n9159 0.00636816
R26695 VSS.n10344 VSS.n10343 0.00636816
R26696 VSS.n10936 VSS.n10935 0.00636816
R26697 VSS.n11528 VSS.n11527 0.00636816
R26698 VSS.n12120 VSS.n12119 0.00636816
R26699 VSS.n12712 VSS.n12711 0.00636816
R26700 VSS.n13304 VSS.n13303 0.00636816
R26701 VSS.n13896 VSS.n13895 0.00636816
R26702 VSS.n14488 VSS.n14487 0.00636816
R26703 VSS.n15080 VSS.n15079 0.00636816
R26704 VSS.n15672 VSS.n15671 0.00636816
R26705 VSS.n6824 VSS.n6809 0.00636816
R26706 VSS.n7384 VSS.n7383 0.00636816
R26707 VSS.n18696 VSS.n18695 0.00636816
R26708 VSS.n647 VSS.n632 0.00636816
R26709 VSS.n1306 VSS.n1291 0.00636816
R26710 VSS.n17268 VSS.n16862 0.00636785
R26711 VSS.n17860 VSS.n17276 0.00636785
R26712 VSS.n18464 VSS.n18432 0.00636785
R26713 VSS.n9911 VSS.n9327 0.00636785
R26714 VSS.n16854 VSS.n16269 0.00636785
R26715 VSS.n16261 VSS.n1441 0.00636785
R26716 VSS.n2207 VSS.n2201 0.00636785
R26717 VSS.n3402 VSS.n2818 0.00636785
R26718 VSS.n3994 VSS.n3410 0.00636785
R26719 VSS.n4586 VSS.n4002 0.00636785
R26720 VSS.n5178 VSS.n4594 0.00636785
R26721 VSS.n2803 VSS.n2797 0.00636785
R26722 VSS.n18884 VSS.n3 0.00636785
R26723 VSS.n6337 VSS.n6331 0.00636785
R26724 VSS.n8135 VSS.n7551 0.00636785
R26725 VSS.n8727 VSS.n8143 0.00636785
R26726 VSS.n9319 VSS.n8735 0.00636785
R26727 VSS.n10503 VSS.n9919 0.00636785
R26728 VSS.n11095 VSS.n10511 0.00636785
R26729 VSS.n11687 VSS.n11103 0.00636785
R26730 VSS.n12279 VSS.n11695 0.00636785
R26731 VSS.n12871 VSS.n12287 0.00636785
R26732 VSS.n13463 VSS.n12879 0.00636785
R26733 VSS.n14055 VSS.n13471 0.00636785
R26734 VSS.n14647 VSS.n14063 0.00636785
R26735 VSS.n15239 VSS.n14655 0.00636785
R26736 VSS.n15831 VSS.n15247 0.00636785
R26737 VSS.n6943 VSS.n6937 0.00636785
R26738 VSS.n7543 VSS.n6958 0.00636785
R26739 VSS.n18855 VSS.n56 0.00636785
R26740 VSS.n50 VSS.n44 0.00636785
R26741 VSS.n1425 VSS.n1419 0.00636785
R26742 VSS.n17146 VSS.n17145 0.00620714
R26743 VSS.n17145 VSS.n16907 0.00620714
R26744 VSS.n17227 VSS.n16875 0.00620714
R26745 VSS.n17245 VSS.n16875 0.00620714
R26746 VSS.n17738 VSS.n17737 0.00620714
R26747 VSS.n17737 VSS.n17321 0.00620714
R26748 VSS.n17819 VSS.n17289 0.00620714
R26749 VSS.n17837 VSS.n17289 0.00620714
R26750 VSS.n18522 VSS.n18521 0.00620714
R26751 VSS.n18521 VSS.n18520 0.00620714
R26752 VSS.n18485 VSS.n18415 0.00620714
R26753 VSS.n18428 VSS.n18415 0.00620714
R26754 VSS.n9788 VSS.n9787 0.00620714
R26755 VSS.n9787 VSS.n9371 0.00620714
R26756 VSS.n9869 VSS.n9340 0.00620714
R26757 VSS.n9887 VSS.n9340 0.00620714
R26758 VSS.n16731 VSS.n16730 0.00620714
R26759 VSS.n16730 VSS.n16313 0.00620714
R26760 VSS.n16812 VSS.n16282 0.00620714
R26761 VSS.n16830 VSS.n16282 0.00620714
R26762 VSS.n16138 VSS.n16137 0.00620714
R26763 VSS.n16137 VSS.n1485 0.00620714
R26764 VSS.n16219 VSS.n1454 0.00620714
R26765 VSS.n16237 VSS.n1454 0.00620714
R26766 VSS.n2112 VSS.n2101 0.00620714
R26767 VSS.n2117 VSS.n2112 0.00620714
R26768 VSS.n2239 VSS.n2238 0.00620714
R26769 VSS.n2238 VSS.n2237 0.00620714
R26770 VSS.n3279 VSS.n3278 0.00620714
R26771 VSS.n3278 VSS.n2862 0.00620714
R26772 VSS.n3360 VSS.n2831 0.00620714
R26773 VSS.n3378 VSS.n2831 0.00620714
R26774 VSS.n3871 VSS.n3870 0.00620714
R26775 VSS.n3870 VSS.n3454 0.00620714
R26776 VSS.n3952 VSS.n3423 0.00620714
R26777 VSS.n3970 VSS.n3423 0.00620714
R26778 VSS.n4463 VSS.n4462 0.00620714
R26779 VSS.n4462 VSS.n4046 0.00620714
R26780 VSS.n4544 VSS.n4015 0.00620714
R26781 VSS.n4562 VSS.n4015 0.00620714
R26782 VSS.n5055 VSS.n5054 0.00620714
R26783 VSS.n5054 VSS.n4638 0.00620714
R26784 VSS.n5136 VSS.n4607 0.00620714
R26785 VSS.n5154 VSS.n4607 0.00620714
R26786 VSS.n2708 VSS.n2697 0.00620714
R26787 VSS.n2713 VSS.n2708 0.00620714
R26788 VSS.n5204 VSS.n5203 0.00620714
R26789 VSS.n5203 VSS.n5202 0.00620714
R26790 VSS.n5669 VSS.n5658 0.00620714
R26791 VSS.n5674 VSS.n5669 0.00620714
R26792 VSS.n5777 VSS.n5776 0.00620714
R26793 VSS.n5776 VSS.n5775 0.00620714
R26794 VSS.n6242 VSS.n6231 0.00620714
R26795 VSS.n6247 VSS.n6242 0.00620714
R26796 VSS.n6369 VSS.n6368 0.00620714
R26797 VSS.n6368 VSS.n6367 0.00620714
R26798 VSS.n8012 VSS.n8011 0.00620714
R26799 VSS.n8011 VSS.n7595 0.00620714
R26800 VSS.n8093 VSS.n7564 0.00620714
R26801 VSS.n8111 VSS.n7564 0.00620714
R26802 VSS.n8604 VSS.n8603 0.00620714
R26803 VSS.n8603 VSS.n8187 0.00620714
R26804 VSS.n8685 VSS.n8156 0.00620714
R26805 VSS.n8703 VSS.n8156 0.00620714
R26806 VSS.n9196 VSS.n9195 0.00620714
R26807 VSS.n9195 VSS.n8779 0.00620714
R26808 VSS.n9277 VSS.n8748 0.00620714
R26809 VSS.n9295 VSS.n8748 0.00620714
R26810 VSS.n10380 VSS.n10379 0.00620714
R26811 VSS.n10379 VSS.n9963 0.00620714
R26812 VSS.n10461 VSS.n9932 0.00620714
R26813 VSS.n10479 VSS.n9932 0.00620714
R26814 VSS.n10972 VSS.n10971 0.00620714
R26815 VSS.n10971 VSS.n10555 0.00620714
R26816 VSS.n11053 VSS.n10524 0.00620714
R26817 VSS.n11071 VSS.n10524 0.00620714
R26818 VSS.n11564 VSS.n11563 0.00620714
R26819 VSS.n11563 VSS.n11147 0.00620714
R26820 VSS.n11645 VSS.n11116 0.00620714
R26821 VSS.n11663 VSS.n11116 0.00620714
R26822 VSS.n12156 VSS.n12155 0.00620714
R26823 VSS.n12155 VSS.n11739 0.00620714
R26824 VSS.n12237 VSS.n11708 0.00620714
R26825 VSS.n12255 VSS.n11708 0.00620714
R26826 VSS.n12748 VSS.n12747 0.00620714
R26827 VSS.n12747 VSS.n12331 0.00620714
R26828 VSS.n12829 VSS.n12300 0.00620714
R26829 VSS.n12847 VSS.n12300 0.00620714
R26830 VSS.n13340 VSS.n13339 0.00620714
R26831 VSS.n13339 VSS.n12923 0.00620714
R26832 VSS.n13421 VSS.n12892 0.00620714
R26833 VSS.n13439 VSS.n12892 0.00620714
R26834 VSS.n13932 VSS.n13931 0.00620714
R26835 VSS.n13931 VSS.n13515 0.00620714
R26836 VSS.n14013 VSS.n13484 0.00620714
R26837 VSS.n14031 VSS.n13484 0.00620714
R26838 VSS.n14524 VSS.n14523 0.00620714
R26839 VSS.n14523 VSS.n14107 0.00620714
R26840 VSS.n14605 VSS.n14076 0.00620714
R26841 VSS.n14623 VSS.n14076 0.00620714
R26842 VSS.n15116 VSS.n15115 0.00620714
R26843 VSS.n15115 VSS.n14699 0.00620714
R26844 VSS.n15197 VSS.n14668 0.00620714
R26845 VSS.n15215 VSS.n14668 0.00620714
R26846 VSS.n15708 VSS.n15707 0.00620714
R26847 VSS.n15707 VSS.n15291 0.00620714
R26848 VSS.n15789 VSS.n15260 0.00620714
R26849 VSS.n15807 VSS.n15260 0.00620714
R26850 VSS.n6848 VSS.n6837 0.00620714
R26851 VSS.n6853 VSS.n6848 0.00620714
R26852 VSS.n15857 VSS.n15856 0.00620714
R26853 VSS.n15856 VSS.n15855 0.00620714
R26854 VSS.n7420 VSS.n7419 0.00620714
R26855 VSS.n7419 VSS.n7002 0.00620714
R26856 VSS.n7501 VSS.n6971 0.00620714
R26857 VSS.n7519 VSS.n6971 0.00620714
R26858 VSS.n18732 VSS.n18731 0.00620714
R26859 VSS.n18731 VSS.n100 0.00620714
R26860 VSS.n18813 VSS.n69 0.00620714
R26861 VSS.n18831 VSS.n69 0.00620714
R26862 VSS.n671 VSS.n660 0.00620714
R26863 VSS.n676 VSS.n671 0.00620714
R26864 VSS.n771 VSS.n770 0.00620714
R26865 VSS.n770 VSS.n769 0.00620714
R26866 VSS.n1330 VSS.n1319 0.00620714
R26867 VSS.n1335 VSS.n1330 0.00620714
R26868 VSS.n17885 VSS.n17884 0.00620714
R26869 VSS.n17884 VSS.n17883 0.00620714
R26870 VSS.n17135 VSS.n16927 0.00587143
R26871 VSS.n17176 VSS.n17175 0.00587143
R26872 VSS.n17192 VSS.n16887 0.00587143
R26873 VSS.n17246 VSS.n16860 0.00587143
R26874 VSS.n17727 VSS.n17341 0.00587143
R26875 VSS.n17768 VSS.n17767 0.00587143
R26876 VSS.n17784 VSS.n17301 0.00587143
R26877 VSS.n17838 VSS.n17274 0.00587143
R26878 VSS.n18329 VSS.n18318 0.00587143
R26879 VSS.n18351 VSS.n18350 0.00587143
R26880 VSS.n18414 VSS.n18413 0.00587143
R26881 VSS.n18469 VSS.n18468 0.00587143
R26882 VSS.n9777 VSS.n9391 0.00587143
R26883 VSS.n9818 VSS.n9817 0.00587143
R26884 VSS.n9834 VSS.n9351 0.00587143
R26885 VSS.n9889 VSS.n9325 0.00587143
R26886 VSS.n16720 VSS.n16333 0.00587143
R26887 VSS.n16761 VSS.n16760 0.00587143
R26888 VSS.n16777 VSS.n16293 0.00587143
R26889 VSS.n16832 VSS.n16267 0.00587143
R26890 VSS.n16127 VSS.n1505 0.00587143
R26891 VSS.n16168 VSS.n16167 0.00587143
R26892 VSS.n16184 VSS.n1465 0.00587143
R26893 VSS.n16239 VSS.n1439 0.00587143
R26894 VSS.n2093 VSS.n2083 0.00587143
R26895 VSS.n2136 VSS.n2135 0.00587143
R26896 VSS.n2167 VSS.n2152 0.00587143
R26897 VSS.n2219 VSS.n2218 0.00587143
R26898 VSS.n3268 VSS.n2882 0.00587143
R26899 VSS.n3309 VSS.n3308 0.00587143
R26900 VSS.n3325 VSS.n2842 0.00587143
R26901 VSS.n3380 VSS.n2816 0.00587143
R26902 VSS.n3860 VSS.n3474 0.00587143
R26903 VSS.n3901 VSS.n3900 0.00587143
R26904 VSS.n3917 VSS.n3434 0.00587143
R26905 VSS.n3972 VSS.n3408 0.00587143
R26906 VSS.n4452 VSS.n4066 0.00587143
R26907 VSS.n4493 VSS.n4492 0.00587143
R26908 VSS.n4509 VSS.n4026 0.00587143
R26909 VSS.n4564 VSS.n4000 0.00587143
R26910 VSS.n5044 VSS.n4658 0.00587143
R26911 VSS.n5085 VSS.n5084 0.00587143
R26912 VSS.n5101 VSS.n4618 0.00587143
R26913 VSS.n5156 VSS.n4592 0.00587143
R26914 VSS.n2689 VSS.n2679 0.00587143
R26915 VSS.n2732 VSS.n2731 0.00587143
R26916 VSS.n2763 VSS.n2748 0.00587143
R26917 VSS.n2815 VSS.n2814 0.00587143
R26918 VSS.n5650 VSS.n5640 0.00587143
R26919 VSS.n5693 VSS.n5692 0.00587143
R26920 VSS.n5724 VSS.n5709 0.00587143
R26921 VSS.n5731 VSS.n1 0.00587143
R26922 VSS.n6223 VSS.n6213 0.00587143
R26923 VSS.n6266 VSS.n6265 0.00587143
R26924 VSS.n6297 VSS.n6282 0.00587143
R26925 VSS.n6349 VSS.n6348 0.00587143
R26926 VSS.n8001 VSS.n7615 0.00587143
R26927 VSS.n8042 VSS.n8041 0.00587143
R26928 VSS.n8058 VSS.n7575 0.00587143
R26929 VSS.n8113 VSS.n7549 0.00587143
R26930 VSS.n8593 VSS.n8207 0.00587143
R26931 VSS.n8634 VSS.n8633 0.00587143
R26932 VSS.n8650 VSS.n8167 0.00587143
R26933 VSS.n8705 VSS.n8141 0.00587143
R26934 VSS.n9185 VSS.n8799 0.00587143
R26935 VSS.n9226 VSS.n9225 0.00587143
R26936 VSS.n9242 VSS.n8759 0.00587143
R26937 VSS.n9297 VSS.n8733 0.00587143
R26938 VSS.n10369 VSS.n9983 0.00587143
R26939 VSS.n10410 VSS.n10409 0.00587143
R26940 VSS.n10426 VSS.n9943 0.00587143
R26941 VSS.n10481 VSS.n9917 0.00587143
R26942 VSS.n10961 VSS.n10575 0.00587143
R26943 VSS.n11002 VSS.n11001 0.00587143
R26944 VSS.n11018 VSS.n10535 0.00587143
R26945 VSS.n11073 VSS.n10509 0.00587143
R26946 VSS.n11553 VSS.n11167 0.00587143
R26947 VSS.n11594 VSS.n11593 0.00587143
R26948 VSS.n11610 VSS.n11127 0.00587143
R26949 VSS.n11665 VSS.n11101 0.00587143
R26950 VSS.n12145 VSS.n11759 0.00587143
R26951 VSS.n12186 VSS.n12185 0.00587143
R26952 VSS.n12202 VSS.n11719 0.00587143
R26953 VSS.n12257 VSS.n11693 0.00587143
R26954 VSS.n12737 VSS.n12351 0.00587143
R26955 VSS.n12778 VSS.n12777 0.00587143
R26956 VSS.n12794 VSS.n12311 0.00587143
R26957 VSS.n12849 VSS.n12285 0.00587143
R26958 VSS.n13329 VSS.n12943 0.00587143
R26959 VSS.n13370 VSS.n13369 0.00587143
R26960 VSS.n13386 VSS.n12903 0.00587143
R26961 VSS.n13441 VSS.n12877 0.00587143
R26962 VSS.n13921 VSS.n13535 0.00587143
R26963 VSS.n13962 VSS.n13961 0.00587143
R26964 VSS.n13978 VSS.n13495 0.00587143
R26965 VSS.n14033 VSS.n13469 0.00587143
R26966 VSS.n14513 VSS.n14127 0.00587143
R26967 VSS.n14554 VSS.n14553 0.00587143
R26968 VSS.n14570 VSS.n14087 0.00587143
R26969 VSS.n14625 VSS.n14061 0.00587143
R26970 VSS.n15105 VSS.n14719 0.00587143
R26971 VSS.n15146 VSS.n15145 0.00587143
R26972 VSS.n15162 VSS.n14679 0.00587143
R26973 VSS.n15217 VSS.n14653 0.00587143
R26974 VSS.n15697 VSS.n15311 0.00587143
R26975 VSS.n15738 VSS.n15737 0.00587143
R26976 VSS.n15754 VSS.n15271 0.00587143
R26977 VSS.n15809 VSS.n15245 0.00587143
R26978 VSS.n6829 VSS.n6819 0.00587143
R26979 VSS.n6872 VSS.n6871 0.00587143
R26980 VSS.n6903 VSS.n6888 0.00587143
R26981 VSS.n6955 VSS.n6954 0.00587143
R26982 VSS.n7409 VSS.n7022 0.00587143
R26983 VSS.n7450 VSS.n7449 0.00587143
R26984 VSS.n7466 VSS.n6982 0.00587143
R26985 VSS.n7521 VSS.n6956 0.00587143
R26986 VSS.n18721 VSS.n120 0.00587143
R26987 VSS.n18762 VSS.n18761 0.00587143
R26988 VSS.n18778 VSS.n80 0.00587143
R26989 VSS.n18833 VSS.n54 0.00587143
R26990 VSS.n652 VSS.n642 0.00587143
R26991 VSS.n695 VSS.n694 0.00587143
R26992 VSS.n726 VSS.n711 0.00587143
R26993 VSS.n733 VSS.n52 0.00587143
R26994 VSS.n1311 VSS.n1301 0.00587143
R26995 VSS.n1354 VSS.n1353 0.00587143
R26996 VSS.n1385 VSS.n1370 0.00587143
R26997 VSS.n1437 VSS.n1436 0.00587143
R26998 VSS.n1228 VSS.n1223 0.00585714
R26999 VSS.n1215 VSS.n1171 0.00585714
R27000 VSS.n17968 VSS.n1180 0.00585714
R27001 VSS.n1267 VSS.n1260 0.00585714
R27002 VSS.n1277 VSS.n1202 0.00585714
R27003 VSS.n17983 VSS.n1164 0.00585714
R27004 VSS.n1173 VSS.n1170 0.00585714
R27005 VSS.n17967 VSS.n17966 0.00585714
R27006 VSS.n923 VSS.n922 0.00585714
R27007 VSS.n1001 VSS.n1000 0.00585714
R27008 VSS.n17011 VSS.n16991 0.00585714
R27009 VSS.n17046 VSS.n17045 0.00585714
R27010 VSS.n17066 VSS.n17065 0.00585714
R27011 VSS.n17078 VSS.n16957 0.00585714
R27012 VSS.n16948 VSS.n16941 0.00585714
R27013 VSS.n1104 VSS.n1103 0.00585714
R27014 VSS.n18027 VSS.n18026 0.00585714
R27015 VSS.n1102 VSS.n1032 0.00585714
R27016 VSS.n18028 VSS.n1035 0.00585714
R27017 VSS.n18016 VSS.n1048 0.00585714
R27018 VSS.n18011 VSS.n1053 0.00585714
R27019 VSS.n17160 VSS.n16919 0.00585714
R27020 VSS.n17202 VSS.n17201 0.00585714
R27021 VSS.n17223 VSS.n16884 0.00585714
R27022 VSS.n17233 VSS.n17232 0.00585714
R27023 VSS.n16889 VSS.n16886 0.00585714
R27024 VSS.n16995 VSS.n16983 0.00585714
R27025 VSS.n17040 VSS.n16981 0.00585714
R27026 VSS.n17067 VSS.n16962 0.00585714
R27027 VSS.n17603 VSS.n17405 0.00585714
R27028 VSS.n17638 VSS.n17637 0.00585714
R27029 VSS.n17658 VSS.n17657 0.00585714
R27030 VSS.n17670 VSS.n17371 0.00585714
R27031 VSS.n17362 VSS.n17355 0.00585714
R27032 VSS.n17534 VSS.n17533 0.00585714
R27033 VSS.n17542 VSS.n17468 0.00585714
R27034 VSS.n17535 VSS.n17472 0.00585714
R27035 VSS.n17541 VSS.n17469 0.00585714
R27036 VSS.n17547 VSS.n17444 0.00585714
R27037 VSS.n17572 VSS.n17440 0.00585714
R27038 VSS.n17752 VSS.n17333 0.00585714
R27039 VSS.n17794 VSS.n17793 0.00585714
R27040 VSS.n17815 VSS.n17298 0.00585714
R27041 VSS.n17825 VSS.n17824 0.00585714
R27042 VSS.n17303 VSS.n17300 0.00585714
R27043 VSS.n17409 VSS.n17397 0.00585714
R27044 VSS.n17632 VSS.n17395 0.00585714
R27045 VSS.n17659 VSS.n17376 0.00585714
R27046 VSS.n18111 VSS.n18110 0.00585714
R27047 VSS.n18119 VSS.n260 0.00585714
R27048 VSS.n18245 VSS.n18240 0.00585714
R27049 VSS.n18232 VSS.n18188 0.00585714
R27050 VSS.n18557 VSS.n18197 0.00585714
R27051 VSS.n18284 VSS.n18277 0.00585714
R27052 VSS.n18294 VSS.n18219 0.00585714
R27053 VSS.n18572 VSS.n18181 0.00585714
R27054 VSS.n18190 VSS.n18187 0.00585714
R27055 VSS.n18556 VSS.n18555 0.00585714
R27056 VSS.n18516 VSS.n18340 0.00585714
R27057 VSS.n18407 VSS.n18406 0.00585714
R27058 VSS.n18443 VSS.n18389 0.00585714
R27059 VSS.n18447 VSS.n18446 0.00585714
R27060 VSS.n18444 VSS.n18391 0.00585714
R27061 VSS.n18112 VSS.n264 0.00585714
R27062 VSS.n18118 VSS.n261 0.00585714
R27063 VSS.n18124 VSS.n236 0.00585714
R27064 VSS.n18149 VSS.n232 0.00585714
R27065 VSS.n9584 VSS.n9583 0.00585714
R27066 VSS.n9592 VSS.n9518 0.00585714
R27067 VSS.n9653 VSS.n9455 0.00585714
R27068 VSS.n9688 VSS.n9687 0.00585714
R27069 VSS.n9708 VSS.n9707 0.00585714
R27070 VSS.n9720 VSS.n9421 0.00585714
R27071 VSS.n9412 VSS.n9405 0.00585714
R27072 VSS.n9459 VSS.n9447 0.00585714
R27073 VSS.n9682 VSS.n9445 0.00585714
R27074 VSS.n9709 VSS.n9426 0.00585714
R27075 VSS.n9802 VSS.n9383 0.00585714
R27076 VSS.n9844 VSS.n9843 0.00585714
R27077 VSS.n9865 VSS.n9348 0.00585714
R27078 VSS.n9875 VSS.n9874 0.00585714
R27079 VSS.n9353 VSS.n9350 0.00585714
R27080 VSS.n9585 VSS.n9522 0.00585714
R27081 VSS.n9591 VSS.n9519 0.00585714
R27082 VSS.n9597 VSS.n9494 0.00585714
R27083 VSS.n9622 VSS.n9490 0.00585714
R27084 VSS.n16515 VSS.n16460 0.00585714
R27085 VSS.n16463 VSS.n16461 0.00585714
R27086 VSS.n16596 VSS.n16397 0.00585714
R27087 VSS.n16631 VSS.n16630 0.00585714
R27088 VSS.n16651 VSS.n16650 0.00585714
R27089 VSS.n16663 VSS.n16363 0.00585714
R27090 VSS.n16354 VSS.n16347 0.00585714
R27091 VSS.n16401 VSS.n16389 0.00585714
R27092 VSS.n16625 VSS.n16387 0.00585714
R27093 VSS.n16652 VSS.n16368 0.00585714
R27094 VSS.n16745 VSS.n16325 0.00585714
R27095 VSS.n16787 VSS.n16786 0.00585714
R27096 VSS.n16808 VSS.n16290 0.00585714
R27097 VSS.n16818 VSS.n16817 0.00585714
R27098 VSS.n16295 VSS.n16292 0.00585714
R27099 VSS.n16516 VSS.n16462 0.00585714
R27100 VSS.n16523 VSS.n16464 0.00585714
R27101 VSS.n16446 VSS.n16443 0.00585714
R27102 VSS.n16441 VSS.n16426 0.00585714
R27103 VSS.n1680 VSS.n1625 0.00585714
R27104 VSS.n1628 VSS.n1626 0.00585714
R27105 VSS.n16003 VSS.n1569 0.00585714
R27106 VSS.n16038 VSS.n16037 0.00585714
R27107 VSS.n16058 VSS.n16057 0.00585714
R27108 VSS.n16070 VSS.n1535 0.00585714
R27109 VSS.n1526 VSS.n1519 0.00585714
R27110 VSS.n1573 VSS.n1561 0.00585714
R27111 VSS.n16032 VSS.n1559 0.00585714
R27112 VSS.n16059 VSS.n1540 0.00585714
R27113 VSS.n16152 VSS.n1497 0.00585714
R27114 VSS.n16194 VSS.n16193 0.00585714
R27115 VSS.n16215 VSS.n1462 0.00585714
R27116 VSS.n16225 VSS.n16224 0.00585714
R27117 VSS.n1467 VSS.n1464 0.00585714
R27118 VSS.n1681 VSS.n1627 0.00585714
R27119 VSS.n1688 VSS.n1629 0.00585714
R27120 VSS.n1611 VSS.n1608 0.00585714
R27121 VSS.n1606 VSS.n1591 0.00585714
R27122 VSS.n1876 VSS.n1875 0.00585714
R27123 VSS.n1884 VSS.n1810 0.00585714
R27124 VSS.n2010 VSS.n2005 0.00585714
R27125 VSS.n1997 VSS.n1953 0.00585714
R27126 VSS.n2322 VSS.n1962 0.00585714
R27127 VSS.n2049 VSS.n2042 0.00585714
R27128 VSS.n2059 VSS.n1984 0.00585714
R27129 VSS.n2337 VSS.n1946 0.00585714
R27130 VSS.n1955 VSS.n1952 0.00585714
R27131 VSS.n2321 VSS.n2320 0.00585714
R27132 VSS.n2276 VSS.n2108 0.00585714
R27133 VSS.n2184 VSS.n2183 0.00585714
R27134 VSS.n2247 VSS.n2159 0.00585714
R27135 VSS.n2243 VSS.n2162 0.00585714
R27136 VSS.n2246 VSS.n2245 0.00585714
R27137 VSS.n1877 VSS.n1814 0.00585714
R27138 VSS.n1883 VSS.n1811 0.00585714
R27139 VSS.n1889 VSS.n1786 0.00585714
R27140 VSS.n1914 VSS.n1782 0.00585714
R27141 VSS.n3075 VSS.n3074 0.00585714
R27142 VSS.n3083 VSS.n3009 0.00585714
R27143 VSS.n3144 VSS.n2946 0.00585714
R27144 VSS.n3179 VSS.n3178 0.00585714
R27145 VSS.n3199 VSS.n3198 0.00585714
R27146 VSS.n3211 VSS.n2912 0.00585714
R27147 VSS.n2903 VSS.n2896 0.00585714
R27148 VSS.n2950 VSS.n2938 0.00585714
R27149 VSS.n3173 VSS.n2936 0.00585714
R27150 VSS.n3200 VSS.n2917 0.00585714
R27151 VSS.n3293 VSS.n2874 0.00585714
R27152 VSS.n3335 VSS.n3334 0.00585714
R27153 VSS.n3356 VSS.n2839 0.00585714
R27154 VSS.n3366 VSS.n3365 0.00585714
R27155 VSS.n2844 VSS.n2841 0.00585714
R27156 VSS.n3076 VSS.n3013 0.00585714
R27157 VSS.n3082 VSS.n3010 0.00585714
R27158 VSS.n3088 VSS.n2985 0.00585714
R27159 VSS.n3113 VSS.n2981 0.00585714
R27160 VSS.n3667 VSS.n3666 0.00585714
R27161 VSS.n3675 VSS.n3601 0.00585714
R27162 VSS.n3736 VSS.n3538 0.00585714
R27163 VSS.n3771 VSS.n3770 0.00585714
R27164 VSS.n3791 VSS.n3790 0.00585714
R27165 VSS.n3803 VSS.n3504 0.00585714
R27166 VSS.n3495 VSS.n3488 0.00585714
R27167 VSS.n3542 VSS.n3530 0.00585714
R27168 VSS.n3765 VSS.n3528 0.00585714
R27169 VSS.n3792 VSS.n3509 0.00585714
R27170 VSS.n3885 VSS.n3466 0.00585714
R27171 VSS.n3927 VSS.n3926 0.00585714
R27172 VSS.n3948 VSS.n3431 0.00585714
R27173 VSS.n3958 VSS.n3957 0.00585714
R27174 VSS.n3436 VSS.n3433 0.00585714
R27175 VSS.n3668 VSS.n3605 0.00585714
R27176 VSS.n3674 VSS.n3602 0.00585714
R27177 VSS.n3680 VSS.n3577 0.00585714
R27178 VSS.n3705 VSS.n3573 0.00585714
R27179 VSS.n4259 VSS.n4258 0.00585714
R27180 VSS.n4267 VSS.n4193 0.00585714
R27181 VSS.n4328 VSS.n4130 0.00585714
R27182 VSS.n4363 VSS.n4362 0.00585714
R27183 VSS.n4383 VSS.n4382 0.00585714
R27184 VSS.n4395 VSS.n4096 0.00585714
R27185 VSS.n4087 VSS.n4080 0.00585714
R27186 VSS.n4134 VSS.n4122 0.00585714
R27187 VSS.n4357 VSS.n4120 0.00585714
R27188 VSS.n4384 VSS.n4101 0.00585714
R27189 VSS.n4477 VSS.n4058 0.00585714
R27190 VSS.n4519 VSS.n4518 0.00585714
R27191 VSS.n4540 VSS.n4023 0.00585714
R27192 VSS.n4550 VSS.n4549 0.00585714
R27193 VSS.n4028 VSS.n4025 0.00585714
R27194 VSS.n4260 VSS.n4197 0.00585714
R27195 VSS.n4266 VSS.n4194 0.00585714
R27196 VSS.n4272 VSS.n4169 0.00585714
R27197 VSS.n4297 VSS.n4165 0.00585714
R27198 VSS.n4851 VSS.n4850 0.00585714
R27199 VSS.n4859 VSS.n4785 0.00585714
R27200 VSS.n4920 VSS.n4722 0.00585714
R27201 VSS.n4955 VSS.n4954 0.00585714
R27202 VSS.n4975 VSS.n4974 0.00585714
R27203 VSS.n4987 VSS.n4688 0.00585714
R27204 VSS.n4679 VSS.n4672 0.00585714
R27205 VSS.n4726 VSS.n4714 0.00585714
R27206 VSS.n4949 VSS.n4712 0.00585714
R27207 VSS.n4976 VSS.n4693 0.00585714
R27208 VSS.n5069 VSS.n4650 0.00585714
R27209 VSS.n5111 VSS.n5110 0.00585714
R27210 VSS.n5132 VSS.n4615 0.00585714
R27211 VSS.n5142 VSS.n5141 0.00585714
R27212 VSS.n4620 VSS.n4617 0.00585714
R27213 VSS.n4852 VSS.n4789 0.00585714
R27214 VSS.n4858 VSS.n4786 0.00585714
R27215 VSS.n4864 VSS.n4761 0.00585714
R27216 VSS.n4889 VSS.n4757 0.00585714
R27217 VSS.n2472 VSS.n2471 0.00585714
R27218 VSS.n2480 VSS.n2406 0.00585714
R27219 VSS.n2606 VSS.n2601 0.00585714
R27220 VSS.n2593 VSS.n2549 0.00585714
R27221 VSS.n5287 VSS.n2558 0.00585714
R27222 VSS.n2645 VSS.n2638 0.00585714
R27223 VSS.n2655 VSS.n2580 0.00585714
R27224 VSS.n5302 VSS.n2542 0.00585714
R27225 VSS.n2551 VSS.n2548 0.00585714
R27226 VSS.n5286 VSS.n5285 0.00585714
R27227 VSS.n5241 VSS.n2704 0.00585714
R27228 VSS.n2780 VSS.n2779 0.00585714
R27229 VSS.n5212 VSS.n2755 0.00585714
R27230 VSS.n5208 VSS.n2758 0.00585714
R27231 VSS.n5211 VSS.n5210 0.00585714
R27232 VSS.n2473 VSS.n2410 0.00585714
R27233 VSS.n2479 VSS.n2407 0.00585714
R27234 VSS.n2485 VSS.n2382 0.00585714
R27235 VSS.n2510 VSS.n2378 0.00585714
R27236 VSS.n5433 VSS.n5432 0.00585714
R27237 VSS.n5441 VSS.n5367 0.00585714
R27238 VSS.n5567 VSS.n5562 0.00585714
R27239 VSS.n5554 VSS.n5510 0.00585714
R27240 VSS.n5860 VSS.n5519 0.00585714
R27241 VSS.n5606 VSS.n5599 0.00585714
R27242 VSS.n5616 VSS.n5541 0.00585714
R27243 VSS.n5875 VSS.n5503 0.00585714
R27244 VSS.n5512 VSS.n5509 0.00585714
R27245 VSS.n5859 VSS.n5858 0.00585714
R27246 VSS.n5814 VSS.n5665 0.00585714
R27247 VSS.n5754 VSS.n5753 0.00585714
R27248 VSS.n5785 VSS.n5716 0.00585714
R27249 VSS.n5781 VSS.n5719 0.00585714
R27250 VSS.n5784 VSS.n5783 0.00585714
R27251 VSS.n5434 VSS.n5371 0.00585714
R27252 VSS.n5440 VSS.n5368 0.00585714
R27253 VSS.n5446 VSS.n5343 0.00585714
R27254 VSS.n5471 VSS.n5339 0.00585714
R27255 VSS.n6006 VSS.n6005 0.00585714
R27256 VSS.n6014 VSS.n5940 0.00585714
R27257 VSS.n6140 VSS.n6135 0.00585714
R27258 VSS.n6127 VSS.n6083 0.00585714
R27259 VSS.n6452 VSS.n6092 0.00585714
R27260 VSS.n6179 VSS.n6172 0.00585714
R27261 VSS.n6189 VSS.n6114 0.00585714
R27262 VSS.n6467 VSS.n6076 0.00585714
R27263 VSS.n6085 VSS.n6082 0.00585714
R27264 VSS.n6451 VSS.n6450 0.00585714
R27265 VSS.n6406 VSS.n6238 0.00585714
R27266 VSS.n6314 VSS.n6313 0.00585714
R27267 VSS.n6377 VSS.n6289 0.00585714
R27268 VSS.n6373 VSS.n6292 0.00585714
R27269 VSS.n6376 VSS.n6375 0.00585714
R27270 VSS.n6007 VSS.n5944 0.00585714
R27271 VSS.n6013 VSS.n5941 0.00585714
R27272 VSS.n6019 VSS.n5916 0.00585714
R27273 VSS.n6044 VSS.n5912 0.00585714
R27274 VSS.n7808 VSS.n7807 0.00585714
R27275 VSS.n7816 VSS.n7742 0.00585714
R27276 VSS.n7877 VSS.n7679 0.00585714
R27277 VSS.n7912 VSS.n7911 0.00585714
R27278 VSS.n7932 VSS.n7931 0.00585714
R27279 VSS.n7944 VSS.n7645 0.00585714
R27280 VSS.n7636 VSS.n7629 0.00585714
R27281 VSS.n7683 VSS.n7671 0.00585714
R27282 VSS.n7906 VSS.n7669 0.00585714
R27283 VSS.n7933 VSS.n7650 0.00585714
R27284 VSS.n8026 VSS.n7607 0.00585714
R27285 VSS.n8068 VSS.n8067 0.00585714
R27286 VSS.n8089 VSS.n7572 0.00585714
R27287 VSS.n8099 VSS.n8098 0.00585714
R27288 VSS.n7577 VSS.n7574 0.00585714
R27289 VSS.n7809 VSS.n7746 0.00585714
R27290 VSS.n7815 VSS.n7743 0.00585714
R27291 VSS.n7821 VSS.n7718 0.00585714
R27292 VSS.n7846 VSS.n7714 0.00585714
R27293 VSS.n8400 VSS.n8399 0.00585714
R27294 VSS.n8408 VSS.n8334 0.00585714
R27295 VSS.n8469 VSS.n8271 0.00585714
R27296 VSS.n8504 VSS.n8503 0.00585714
R27297 VSS.n8524 VSS.n8523 0.00585714
R27298 VSS.n8536 VSS.n8237 0.00585714
R27299 VSS.n8228 VSS.n8221 0.00585714
R27300 VSS.n8275 VSS.n8263 0.00585714
R27301 VSS.n8498 VSS.n8261 0.00585714
R27302 VSS.n8525 VSS.n8242 0.00585714
R27303 VSS.n8618 VSS.n8199 0.00585714
R27304 VSS.n8660 VSS.n8659 0.00585714
R27305 VSS.n8681 VSS.n8164 0.00585714
R27306 VSS.n8691 VSS.n8690 0.00585714
R27307 VSS.n8169 VSS.n8166 0.00585714
R27308 VSS.n8401 VSS.n8338 0.00585714
R27309 VSS.n8407 VSS.n8335 0.00585714
R27310 VSS.n8413 VSS.n8310 0.00585714
R27311 VSS.n8438 VSS.n8306 0.00585714
R27312 VSS.n8992 VSS.n8991 0.00585714
R27313 VSS.n9000 VSS.n8926 0.00585714
R27314 VSS.n9061 VSS.n8863 0.00585714
R27315 VSS.n9096 VSS.n9095 0.00585714
R27316 VSS.n9116 VSS.n9115 0.00585714
R27317 VSS.n9128 VSS.n8829 0.00585714
R27318 VSS.n8820 VSS.n8813 0.00585714
R27319 VSS.n8867 VSS.n8855 0.00585714
R27320 VSS.n9090 VSS.n8853 0.00585714
R27321 VSS.n9117 VSS.n8834 0.00585714
R27322 VSS.n9210 VSS.n8791 0.00585714
R27323 VSS.n9252 VSS.n9251 0.00585714
R27324 VSS.n9273 VSS.n8756 0.00585714
R27325 VSS.n9283 VSS.n9282 0.00585714
R27326 VSS.n8761 VSS.n8758 0.00585714
R27327 VSS.n8993 VSS.n8930 0.00585714
R27328 VSS.n8999 VSS.n8927 0.00585714
R27329 VSS.n9005 VSS.n8902 0.00585714
R27330 VSS.n9030 VSS.n8898 0.00585714
R27331 VSS.n10176 VSS.n10175 0.00585714
R27332 VSS.n10184 VSS.n10110 0.00585714
R27333 VSS.n10245 VSS.n10047 0.00585714
R27334 VSS.n10280 VSS.n10279 0.00585714
R27335 VSS.n10300 VSS.n10299 0.00585714
R27336 VSS.n10312 VSS.n10013 0.00585714
R27337 VSS.n10004 VSS.n9997 0.00585714
R27338 VSS.n10051 VSS.n10039 0.00585714
R27339 VSS.n10274 VSS.n10037 0.00585714
R27340 VSS.n10301 VSS.n10018 0.00585714
R27341 VSS.n10394 VSS.n9975 0.00585714
R27342 VSS.n10436 VSS.n10435 0.00585714
R27343 VSS.n10457 VSS.n9940 0.00585714
R27344 VSS.n10467 VSS.n10466 0.00585714
R27345 VSS.n9945 VSS.n9942 0.00585714
R27346 VSS.n10177 VSS.n10114 0.00585714
R27347 VSS.n10183 VSS.n10111 0.00585714
R27348 VSS.n10189 VSS.n10086 0.00585714
R27349 VSS.n10214 VSS.n10082 0.00585714
R27350 VSS.n10768 VSS.n10767 0.00585714
R27351 VSS.n10776 VSS.n10702 0.00585714
R27352 VSS.n10837 VSS.n10639 0.00585714
R27353 VSS.n10872 VSS.n10871 0.00585714
R27354 VSS.n10892 VSS.n10891 0.00585714
R27355 VSS.n10904 VSS.n10605 0.00585714
R27356 VSS.n10596 VSS.n10589 0.00585714
R27357 VSS.n10643 VSS.n10631 0.00585714
R27358 VSS.n10866 VSS.n10629 0.00585714
R27359 VSS.n10893 VSS.n10610 0.00585714
R27360 VSS.n10986 VSS.n10567 0.00585714
R27361 VSS.n11028 VSS.n11027 0.00585714
R27362 VSS.n11049 VSS.n10532 0.00585714
R27363 VSS.n11059 VSS.n11058 0.00585714
R27364 VSS.n10537 VSS.n10534 0.00585714
R27365 VSS.n10769 VSS.n10706 0.00585714
R27366 VSS.n10775 VSS.n10703 0.00585714
R27367 VSS.n10781 VSS.n10678 0.00585714
R27368 VSS.n10806 VSS.n10674 0.00585714
R27369 VSS.n11360 VSS.n11359 0.00585714
R27370 VSS.n11368 VSS.n11294 0.00585714
R27371 VSS.n11429 VSS.n11231 0.00585714
R27372 VSS.n11464 VSS.n11463 0.00585714
R27373 VSS.n11484 VSS.n11483 0.00585714
R27374 VSS.n11496 VSS.n11197 0.00585714
R27375 VSS.n11188 VSS.n11181 0.00585714
R27376 VSS.n11235 VSS.n11223 0.00585714
R27377 VSS.n11458 VSS.n11221 0.00585714
R27378 VSS.n11485 VSS.n11202 0.00585714
R27379 VSS.n11578 VSS.n11159 0.00585714
R27380 VSS.n11620 VSS.n11619 0.00585714
R27381 VSS.n11641 VSS.n11124 0.00585714
R27382 VSS.n11651 VSS.n11650 0.00585714
R27383 VSS.n11129 VSS.n11126 0.00585714
R27384 VSS.n11361 VSS.n11298 0.00585714
R27385 VSS.n11367 VSS.n11295 0.00585714
R27386 VSS.n11373 VSS.n11270 0.00585714
R27387 VSS.n11398 VSS.n11266 0.00585714
R27388 VSS.n11952 VSS.n11951 0.00585714
R27389 VSS.n11960 VSS.n11886 0.00585714
R27390 VSS.n12021 VSS.n11823 0.00585714
R27391 VSS.n12056 VSS.n12055 0.00585714
R27392 VSS.n12076 VSS.n12075 0.00585714
R27393 VSS.n12088 VSS.n11789 0.00585714
R27394 VSS.n11780 VSS.n11773 0.00585714
R27395 VSS.n11827 VSS.n11815 0.00585714
R27396 VSS.n12050 VSS.n11813 0.00585714
R27397 VSS.n12077 VSS.n11794 0.00585714
R27398 VSS.n12170 VSS.n11751 0.00585714
R27399 VSS.n12212 VSS.n12211 0.00585714
R27400 VSS.n12233 VSS.n11716 0.00585714
R27401 VSS.n12243 VSS.n12242 0.00585714
R27402 VSS.n11721 VSS.n11718 0.00585714
R27403 VSS.n11953 VSS.n11890 0.00585714
R27404 VSS.n11959 VSS.n11887 0.00585714
R27405 VSS.n11965 VSS.n11862 0.00585714
R27406 VSS.n11990 VSS.n11858 0.00585714
R27407 VSS.n12544 VSS.n12543 0.00585714
R27408 VSS.n12552 VSS.n12478 0.00585714
R27409 VSS.n12613 VSS.n12415 0.00585714
R27410 VSS.n12648 VSS.n12647 0.00585714
R27411 VSS.n12668 VSS.n12667 0.00585714
R27412 VSS.n12680 VSS.n12381 0.00585714
R27413 VSS.n12372 VSS.n12365 0.00585714
R27414 VSS.n12419 VSS.n12407 0.00585714
R27415 VSS.n12642 VSS.n12405 0.00585714
R27416 VSS.n12669 VSS.n12386 0.00585714
R27417 VSS.n12762 VSS.n12343 0.00585714
R27418 VSS.n12804 VSS.n12803 0.00585714
R27419 VSS.n12825 VSS.n12308 0.00585714
R27420 VSS.n12835 VSS.n12834 0.00585714
R27421 VSS.n12313 VSS.n12310 0.00585714
R27422 VSS.n12545 VSS.n12482 0.00585714
R27423 VSS.n12551 VSS.n12479 0.00585714
R27424 VSS.n12557 VSS.n12454 0.00585714
R27425 VSS.n12582 VSS.n12450 0.00585714
R27426 VSS.n13136 VSS.n13135 0.00585714
R27427 VSS.n13144 VSS.n13070 0.00585714
R27428 VSS.n13205 VSS.n13007 0.00585714
R27429 VSS.n13240 VSS.n13239 0.00585714
R27430 VSS.n13260 VSS.n13259 0.00585714
R27431 VSS.n13272 VSS.n12973 0.00585714
R27432 VSS.n12964 VSS.n12957 0.00585714
R27433 VSS.n13011 VSS.n12999 0.00585714
R27434 VSS.n13234 VSS.n12997 0.00585714
R27435 VSS.n13261 VSS.n12978 0.00585714
R27436 VSS.n13354 VSS.n12935 0.00585714
R27437 VSS.n13396 VSS.n13395 0.00585714
R27438 VSS.n13417 VSS.n12900 0.00585714
R27439 VSS.n13427 VSS.n13426 0.00585714
R27440 VSS.n12905 VSS.n12902 0.00585714
R27441 VSS.n13137 VSS.n13074 0.00585714
R27442 VSS.n13143 VSS.n13071 0.00585714
R27443 VSS.n13149 VSS.n13046 0.00585714
R27444 VSS.n13174 VSS.n13042 0.00585714
R27445 VSS.n13728 VSS.n13727 0.00585714
R27446 VSS.n13736 VSS.n13662 0.00585714
R27447 VSS.n13797 VSS.n13599 0.00585714
R27448 VSS.n13832 VSS.n13831 0.00585714
R27449 VSS.n13852 VSS.n13851 0.00585714
R27450 VSS.n13864 VSS.n13565 0.00585714
R27451 VSS.n13556 VSS.n13549 0.00585714
R27452 VSS.n13603 VSS.n13591 0.00585714
R27453 VSS.n13826 VSS.n13589 0.00585714
R27454 VSS.n13853 VSS.n13570 0.00585714
R27455 VSS.n13946 VSS.n13527 0.00585714
R27456 VSS.n13988 VSS.n13987 0.00585714
R27457 VSS.n14009 VSS.n13492 0.00585714
R27458 VSS.n14019 VSS.n14018 0.00585714
R27459 VSS.n13497 VSS.n13494 0.00585714
R27460 VSS.n13729 VSS.n13666 0.00585714
R27461 VSS.n13735 VSS.n13663 0.00585714
R27462 VSS.n13741 VSS.n13638 0.00585714
R27463 VSS.n13766 VSS.n13634 0.00585714
R27464 VSS.n14320 VSS.n14319 0.00585714
R27465 VSS.n14328 VSS.n14254 0.00585714
R27466 VSS.n14389 VSS.n14191 0.00585714
R27467 VSS.n14424 VSS.n14423 0.00585714
R27468 VSS.n14444 VSS.n14443 0.00585714
R27469 VSS.n14456 VSS.n14157 0.00585714
R27470 VSS.n14148 VSS.n14141 0.00585714
R27471 VSS.n14195 VSS.n14183 0.00585714
R27472 VSS.n14418 VSS.n14181 0.00585714
R27473 VSS.n14445 VSS.n14162 0.00585714
R27474 VSS.n14538 VSS.n14119 0.00585714
R27475 VSS.n14580 VSS.n14579 0.00585714
R27476 VSS.n14601 VSS.n14084 0.00585714
R27477 VSS.n14611 VSS.n14610 0.00585714
R27478 VSS.n14089 VSS.n14086 0.00585714
R27479 VSS.n14321 VSS.n14258 0.00585714
R27480 VSS.n14327 VSS.n14255 0.00585714
R27481 VSS.n14333 VSS.n14230 0.00585714
R27482 VSS.n14358 VSS.n14226 0.00585714
R27483 VSS.n14912 VSS.n14911 0.00585714
R27484 VSS.n14920 VSS.n14846 0.00585714
R27485 VSS.n14981 VSS.n14783 0.00585714
R27486 VSS.n15016 VSS.n15015 0.00585714
R27487 VSS.n15036 VSS.n15035 0.00585714
R27488 VSS.n15048 VSS.n14749 0.00585714
R27489 VSS.n14740 VSS.n14733 0.00585714
R27490 VSS.n14787 VSS.n14775 0.00585714
R27491 VSS.n15010 VSS.n14773 0.00585714
R27492 VSS.n15037 VSS.n14754 0.00585714
R27493 VSS.n15130 VSS.n14711 0.00585714
R27494 VSS.n15172 VSS.n15171 0.00585714
R27495 VSS.n15193 VSS.n14676 0.00585714
R27496 VSS.n15203 VSS.n15202 0.00585714
R27497 VSS.n14681 VSS.n14678 0.00585714
R27498 VSS.n14913 VSS.n14850 0.00585714
R27499 VSS.n14919 VSS.n14847 0.00585714
R27500 VSS.n14925 VSS.n14822 0.00585714
R27501 VSS.n14950 VSS.n14818 0.00585714
R27502 VSS.n15504 VSS.n15503 0.00585714
R27503 VSS.n15512 VSS.n15438 0.00585714
R27504 VSS.n15573 VSS.n15375 0.00585714
R27505 VSS.n15608 VSS.n15607 0.00585714
R27506 VSS.n15628 VSS.n15627 0.00585714
R27507 VSS.n15640 VSS.n15341 0.00585714
R27508 VSS.n15332 VSS.n15325 0.00585714
R27509 VSS.n15379 VSS.n15367 0.00585714
R27510 VSS.n15602 VSS.n15365 0.00585714
R27511 VSS.n15629 VSS.n15346 0.00585714
R27512 VSS.n15722 VSS.n15303 0.00585714
R27513 VSS.n15764 VSS.n15763 0.00585714
R27514 VSS.n15785 VSS.n15268 0.00585714
R27515 VSS.n15795 VSS.n15794 0.00585714
R27516 VSS.n15273 VSS.n15270 0.00585714
R27517 VSS.n15505 VSS.n15442 0.00585714
R27518 VSS.n15511 VSS.n15439 0.00585714
R27519 VSS.n15517 VSS.n15414 0.00585714
R27520 VSS.n15542 VSS.n15410 0.00585714
R27521 VSS.n6612 VSS.n6611 0.00585714
R27522 VSS.n6620 VSS.n6546 0.00585714
R27523 VSS.n6746 VSS.n6741 0.00585714
R27524 VSS.n6733 VSS.n6689 0.00585714
R27525 VSS.n15940 VSS.n6698 0.00585714
R27526 VSS.n6785 VSS.n6778 0.00585714
R27527 VSS.n6795 VSS.n6720 0.00585714
R27528 VSS.n15955 VSS.n6682 0.00585714
R27529 VSS.n6691 VSS.n6688 0.00585714
R27530 VSS.n15939 VSS.n15938 0.00585714
R27531 VSS.n15894 VSS.n6844 0.00585714
R27532 VSS.n6920 VSS.n6919 0.00585714
R27533 VSS.n15865 VSS.n6895 0.00585714
R27534 VSS.n15861 VSS.n6898 0.00585714
R27535 VSS.n15864 VSS.n15863 0.00585714
R27536 VSS.n6613 VSS.n6550 0.00585714
R27537 VSS.n6619 VSS.n6547 0.00585714
R27538 VSS.n6625 VSS.n6522 0.00585714
R27539 VSS.n6650 VSS.n6518 0.00585714
R27540 VSS.n7204 VSS.n7149 0.00585714
R27541 VSS.n7152 VSS.n7150 0.00585714
R27542 VSS.n7285 VSS.n7086 0.00585714
R27543 VSS.n7320 VSS.n7319 0.00585714
R27544 VSS.n7340 VSS.n7339 0.00585714
R27545 VSS.n7352 VSS.n7052 0.00585714
R27546 VSS.n7043 VSS.n7036 0.00585714
R27547 VSS.n7090 VSS.n7078 0.00585714
R27548 VSS.n7314 VSS.n7076 0.00585714
R27549 VSS.n7341 VSS.n7057 0.00585714
R27550 VSS.n7434 VSS.n7014 0.00585714
R27551 VSS.n7476 VSS.n7475 0.00585714
R27552 VSS.n7497 VSS.n6979 0.00585714
R27553 VSS.n7507 VSS.n7506 0.00585714
R27554 VSS.n6984 VSS.n6981 0.00585714
R27555 VSS.n7205 VSS.n7151 0.00585714
R27556 VSS.n7212 VSS.n7153 0.00585714
R27557 VSS.n7135 VSS.n7132 0.00585714
R27558 VSS.n7130 VSS.n7115 0.00585714
R27559 VSS.n369 VSS.n367 0.00585714
R27560 VSS.n436 VSS.n435 0.00585714
R27561 VSS.n18597 VSS.n184 0.00585714
R27562 VSS.n18632 VSS.n18631 0.00585714
R27563 VSS.n18652 VSS.n18651 0.00585714
R27564 VSS.n18664 VSS.n150 0.00585714
R27565 VSS.n141 VSS.n134 0.00585714
R27566 VSS.n188 VSS.n176 0.00585714
R27567 VSS.n18626 VSS.n174 0.00585714
R27568 VSS.n18653 VSS.n155 0.00585714
R27569 VSS.n18746 VSS.n112 0.00585714
R27570 VSS.n18788 VSS.n18787 0.00585714
R27571 VSS.n18809 VSS.n77 0.00585714
R27572 VSS.n18819 VSS.n18818 0.00585714
R27573 VSS.n82 VSS.n79 0.00585714
R27574 VSS.n368 VSS.n299 0.00585714
R27575 VSS.n437 VSS.n302 0.00585714
R27576 VSS.n425 VSS.n315 0.00585714
R27577 VSS.n420 VSS.n320 0.00585714
R27578 VSS.n569 VSS.n566 0.00585714
R27579 VSS.n553 VSS.n509 0.00585714
R27580 VSS.n854 VSS.n518 0.00585714
R27581 VSS.n608 VSS.n601 0.00585714
R27582 VSS.n618 VSS.n540 0.00585714
R27583 VSS.n869 VSS.n502 0.00585714
R27584 VSS.n511 VSS.n508 0.00585714
R27585 VSS.n853 VSS.n852 0.00585714
R27586 VSS.n808 VSS.n667 0.00585714
R27587 VSS.n752 VSS.n751 0.00585714
R27588 VSS.n779 VSS.n718 0.00585714
R27589 VSS.n775 VSS.n721 0.00585714
R27590 VSS.n778 VSS.n777 0.00585714
R27591 VSS.n921 VSS.n465 0.00585714
R27592 VSS.n1002 VSS.n468 0.00585714
R27593 VSS.n990 VSS.n481 0.00585714
R27594 VSS.n985 VSS.n486 0.00585714
R27595 VSS.n17922 VSS.n1326 0.00585714
R27596 VSS.n1402 VSS.n1401 0.00585714
R27597 VSS.n17893 VSS.n1377 0.00585714
R27598 VSS.n17889 VSS.n1380 0.00585714
R27599 VSS.n17892 VSS.n17891 0.00585714
R27600 VSS.n977 VSS.n494 0.00565497
R27601 VSS.n18003 VSS.n1061 0.00565497
R27602 VSS.n17597 VSS.n17424 0.00565497
R27603 VSS.n18174 VSS.n216 0.00565497
R27604 VSS.n9647 VSS.n9474 0.00565497
R27605 VSS.n16590 VSS.n16416 0.00565497
R27606 VSS.n15997 VSS.n1581 0.00565497
R27607 VSS.n1939 VSS.n1766 0.00565497
R27608 VSS.n3138 VSS.n2965 0.00565497
R27609 VSS.n3730 VSS.n3557 0.00565497
R27610 VSS.n4322 VSS.n4149 0.00565497
R27611 VSS.n4914 VSS.n4741 0.00565497
R27612 VSS.n2535 VSS.n2362 0.00565497
R27613 VSS.n5496 VSS.n5323 0.00565497
R27614 VSS.n6069 VSS.n5896 0.00565497
R27615 VSS.n7871 VSS.n7698 0.00565497
R27616 VSS.n8463 VSS.n8290 0.00565497
R27617 VSS.n9055 VSS.n8882 0.00565497
R27618 VSS.n10239 VSS.n10066 0.00565497
R27619 VSS.n10831 VSS.n10658 0.00565497
R27620 VSS.n11423 VSS.n11250 0.00565497
R27621 VSS.n12015 VSS.n11842 0.00565497
R27622 VSS.n12607 VSS.n12434 0.00565497
R27623 VSS.n13199 VSS.n13026 0.00565497
R27624 VSS.n13791 VSS.n13618 0.00565497
R27625 VSS.n14383 VSS.n14210 0.00565497
R27626 VSS.n14975 VSS.n14802 0.00565497
R27627 VSS.n15567 VSS.n15394 0.00565497
R27628 VSS.n6675 VSS.n6502 0.00565497
R27629 VSS.n7279 VSS.n7105 0.00565497
R27630 VSS.n18591 VSS.n196 0.00565497
R27631 VSS.n17954 VSS.n1195 0.00511752
R27632 VSS.n17131 VSS.n16935 0.00511752
R27633 VSS.n17723 VSS.n17349 0.00511752
R27634 VSS.n18543 VSS.n18212 0.00511752
R27635 VSS.n9773 VSS.n9399 0.00511752
R27636 VSS.n16716 VSS.n16341 0.00511752
R27637 VSS.n16123 VSS.n1513 0.00511752
R27638 VSS.n2308 VSS.n1977 0.00511752
R27639 VSS.n3264 VSS.n2890 0.00511752
R27640 VSS.n3856 VSS.n3482 0.00511752
R27641 VSS.n4448 VSS.n4074 0.00511752
R27642 VSS.n5040 VSS.n4666 0.00511752
R27643 VSS.n5273 VSS.n2573 0.00511752
R27644 VSS.n5846 VSS.n5534 0.00511752
R27645 VSS.n6438 VSS.n6107 0.00511752
R27646 VSS.n7997 VSS.n7623 0.00511752
R27647 VSS.n8589 VSS.n8215 0.00511752
R27648 VSS.n9181 VSS.n8807 0.00511752
R27649 VSS.n10365 VSS.n9991 0.00511752
R27650 VSS.n10957 VSS.n10583 0.00511752
R27651 VSS.n11549 VSS.n11175 0.00511752
R27652 VSS.n12141 VSS.n11767 0.00511752
R27653 VSS.n12733 VSS.n12359 0.00511752
R27654 VSS.n13325 VSS.n12951 0.00511752
R27655 VSS.n13917 VSS.n13543 0.00511752
R27656 VSS.n14509 VSS.n14135 0.00511752
R27657 VSS.n15101 VSS.n14727 0.00511752
R27658 VSS.n15693 VSS.n15319 0.00511752
R27659 VSS.n15926 VSS.n6713 0.00511752
R27660 VSS.n7405 VSS.n7030 0.00511752
R27661 VSS.n18717 VSS.n128 0.00511752
R27662 VSS.n840 VSS.n533 0.00511752
R27663 VSS.n17990 VSS.n1161 0.00496429
R27664 VSS.n17986 VSS.n1164 0.00496429
R27665 VSS.n17962 VSS.n1187 0.00496429
R27666 VSS.n17959 VSS.n1187 0.00496429
R27667 VSS.n17956 VSS.n1193 0.00496429
R27668 VSS.n951 VSS.n944 0.00496429
R27669 VSS.n962 VSS.n887 0.00496429
R27670 VSS.n1132 VSS.n1125 0.00496429
R27671 VSS.n1143 VSS.n1068 0.00496429
R27672 VSS.n18039 VSS.n1026 0.00496429
R27673 VSS.n18035 VSS.n1029 0.00496429
R27674 VSS.n18032 VSS.n1029 0.00496429
R27675 VSS.n18008 VSS.n1053 0.00496429
R27676 VSS.n18005 VSS.n1059 0.00496429
R27677 VSS.n17243 VSS.n16871 0.00496429
R27678 VSS.n17189 VSS.n17188 0.00496429
R27679 VSS.n17244 VSS.n16877 0.00496429
R27680 VSS.n17019 VSS.n16997 0.00496429
R27681 VSS.n17022 VSS.n16995 0.00496429
R27682 VSS.n16960 VSS.n16945 0.00496429
R27683 VSS.n17090 VSS.n16945 0.00496429
R27684 VSS.n17093 VSS.n16933 0.00496429
R27685 VSS.n17566 VSS.n17565 0.00496429
R27686 VSS.n17434 VSS.n17431 0.00496429
R27687 VSS.n17513 VSS.n17491 0.00496429
R27688 VSS.n17516 VSS.n17489 0.00496429
R27689 VSS.n17489 VSS.n17471 0.00496429
R27690 VSS.n17575 VSS.n17440 0.00496429
R27691 VSS.n17578 VSS.n17422 0.00496429
R27692 VSS.n17835 VSS.n17285 0.00496429
R27693 VSS.n17781 VSS.n17780 0.00496429
R27694 VSS.n17836 VSS.n17291 0.00496429
R27695 VSS.n17611 VSS.n17411 0.00496429
R27696 VSS.n17614 VSS.n17409 0.00496429
R27697 VSS.n17374 VSS.n17359 0.00496429
R27698 VSS.n17682 VSS.n17359 0.00496429
R27699 VSS.n17685 VSS.n17347 0.00496429
R27700 VSS.n18143 VSS.n18142 0.00496429
R27701 VSS.n226 VSS.n223 0.00496429
R27702 VSS.n18579 VSS.n18178 0.00496429
R27703 VSS.n18575 VSS.n18181 0.00496429
R27704 VSS.n18551 VSS.n18204 0.00496429
R27705 VSS.n18548 VSS.n18204 0.00496429
R27706 VSS.n18545 VSS.n18210 0.00496429
R27707 VSS.n18478 VSS.n18422 0.00496429
R27708 VSS.n18502 VSS.n18501 0.00496429
R27709 VSS.n18477 VSS.n18424 0.00496429
R27710 VSS.n18090 VSS.n283 0.00496429
R27711 VSS.n18093 VSS.n281 0.00496429
R27712 VSS.n281 VSS.n263 0.00496429
R27713 VSS.n18152 VSS.n232 0.00496429
R27714 VSS.n18155 VSS.n214 0.00496429
R27715 VSS.n9616 VSS.n9615 0.00496429
R27716 VSS.n9484 VSS.n9481 0.00496429
R27717 VSS.n9661 VSS.n9461 0.00496429
R27718 VSS.n9664 VSS.n9459 0.00496429
R27719 VSS.n9424 VSS.n9409 0.00496429
R27720 VSS.n9732 VSS.n9409 0.00496429
R27721 VSS.n9735 VSS.n9397 0.00496429
R27722 VSS.n9885 VSS.n9336 0.00496429
R27723 VSS.n9831 VSS.n9830 0.00496429
R27724 VSS.n9886 VSS.n9338 0.00496429
R27725 VSS.n9563 VSS.n9541 0.00496429
R27726 VSS.n9566 VSS.n9539 0.00496429
R27727 VSS.n9539 VSS.n9521 0.00496429
R27728 VSS.n9625 VSS.n9490 0.00496429
R27729 VSS.n9628 VSS.n9472 0.00496429
R27730 VSS.n16558 VSS.n16438 0.00496429
R27731 VSS.n16429 VSS.n16422 0.00496429
R27732 VSS.n16604 VSS.n16403 0.00496429
R27733 VSS.n16607 VSS.n16401 0.00496429
R27734 VSS.n16366 VSS.n16351 0.00496429
R27735 VSS.n16675 VSS.n16351 0.00496429
R27736 VSS.n16678 VSS.n16339 0.00496429
R27737 VSS.n16828 VSS.n16278 0.00496429
R27738 VSS.n16774 VSS.n16773 0.00496429
R27739 VSS.n16829 VSS.n16280 0.00496429
R27740 VSS.n16499 VSS.n16478 0.00496429
R27741 VSS.n16502 VSS.n16476 0.00496429
R27742 VSS.n16476 VSS.n16466 0.00496429
R27743 VSS.n16571 VSS.n16426 0.00496429
R27744 VSS.n16574 VSS.n16414 0.00496429
R27745 VSS.n1723 VSS.n1603 0.00496429
R27746 VSS.n1594 VSS.n1587 0.00496429
R27747 VSS.n16011 VSS.n1575 0.00496429
R27748 VSS.n16014 VSS.n1573 0.00496429
R27749 VSS.n1538 VSS.n1523 0.00496429
R27750 VSS.n16082 VSS.n1523 0.00496429
R27751 VSS.n16085 VSS.n1511 0.00496429
R27752 VSS.n16235 VSS.n1450 0.00496429
R27753 VSS.n16181 VSS.n16180 0.00496429
R27754 VSS.n16236 VSS.n1452 0.00496429
R27755 VSS.n1664 VSS.n1643 0.00496429
R27756 VSS.n1667 VSS.n1641 0.00496429
R27757 VSS.n1641 VSS.n1631 0.00496429
R27758 VSS.n1736 VSS.n1591 0.00496429
R27759 VSS.n1739 VSS.n1579 0.00496429
R27760 VSS.n1908 VSS.n1907 0.00496429
R27761 VSS.n1776 VSS.n1773 0.00496429
R27762 VSS.n2344 VSS.n1943 0.00496429
R27763 VSS.n2340 VSS.n1946 0.00496429
R27764 VSS.n2316 VSS.n1969 0.00496429
R27765 VSS.n2313 VSS.n1969 0.00496429
R27766 VSS.n2310 VSS.n1975 0.00496429
R27767 VSS.n2235 VSS.n2234 0.00496429
R27768 VSS.n2149 VSS.n2148 0.00496429
R27769 VSS.n2236 VSS.n2170 0.00496429
R27770 VSS.n1855 VSS.n1833 0.00496429
R27771 VSS.n1858 VSS.n1831 0.00496429
R27772 VSS.n1831 VSS.n1813 0.00496429
R27773 VSS.n1917 VSS.n1782 0.00496429
R27774 VSS.n1920 VSS.n1764 0.00496429
R27775 VSS.n3107 VSS.n3106 0.00496429
R27776 VSS.n2975 VSS.n2972 0.00496429
R27777 VSS.n3152 VSS.n2952 0.00496429
R27778 VSS.n3155 VSS.n2950 0.00496429
R27779 VSS.n2915 VSS.n2900 0.00496429
R27780 VSS.n3223 VSS.n2900 0.00496429
R27781 VSS.n3226 VSS.n2888 0.00496429
R27782 VSS.n3376 VSS.n2827 0.00496429
R27783 VSS.n3322 VSS.n3321 0.00496429
R27784 VSS.n3377 VSS.n2829 0.00496429
R27785 VSS.n3054 VSS.n3032 0.00496429
R27786 VSS.n3057 VSS.n3030 0.00496429
R27787 VSS.n3030 VSS.n3012 0.00496429
R27788 VSS.n3116 VSS.n2981 0.00496429
R27789 VSS.n3119 VSS.n2963 0.00496429
R27790 VSS.n3699 VSS.n3698 0.00496429
R27791 VSS.n3567 VSS.n3564 0.00496429
R27792 VSS.n3744 VSS.n3544 0.00496429
R27793 VSS.n3747 VSS.n3542 0.00496429
R27794 VSS.n3507 VSS.n3492 0.00496429
R27795 VSS.n3815 VSS.n3492 0.00496429
R27796 VSS.n3818 VSS.n3480 0.00496429
R27797 VSS.n3968 VSS.n3419 0.00496429
R27798 VSS.n3914 VSS.n3913 0.00496429
R27799 VSS.n3969 VSS.n3421 0.00496429
R27800 VSS.n3646 VSS.n3624 0.00496429
R27801 VSS.n3649 VSS.n3622 0.00496429
R27802 VSS.n3622 VSS.n3604 0.00496429
R27803 VSS.n3708 VSS.n3573 0.00496429
R27804 VSS.n3711 VSS.n3555 0.00496429
R27805 VSS.n4291 VSS.n4290 0.00496429
R27806 VSS.n4159 VSS.n4156 0.00496429
R27807 VSS.n4336 VSS.n4136 0.00496429
R27808 VSS.n4339 VSS.n4134 0.00496429
R27809 VSS.n4099 VSS.n4084 0.00496429
R27810 VSS.n4407 VSS.n4084 0.00496429
R27811 VSS.n4410 VSS.n4072 0.00496429
R27812 VSS.n4560 VSS.n4011 0.00496429
R27813 VSS.n4506 VSS.n4505 0.00496429
R27814 VSS.n4561 VSS.n4013 0.00496429
R27815 VSS.n4238 VSS.n4216 0.00496429
R27816 VSS.n4241 VSS.n4214 0.00496429
R27817 VSS.n4214 VSS.n4196 0.00496429
R27818 VSS.n4300 VSS.n4165 0.00496429
R27819 VSS.n4303 VSS.n4147 0.00496429
R27820 VSS.n4883 VSS.n4882 0.00496429
R27821 VSS.n4751 VSS.n4748 0.00496429
R27822 VSS.n4928 VSS.n4728 0.00496429
R27823 VSS.n4931 VSS.n4726 0.00496429
R27824 VSS.n4691 VSS.n4676 0.00496429
R27825 VSS.n4999 VSS.n4676 0.00496429
R27826 VSS.n5002 VSS.n4664 0.00496429
R27827 VSS.n5152 VSS.n4603 0.00496429
R27828 VSS.n5098 VSS.n5097 0.00496429
R27829 VSS.n5153 VSS.n4605 0.00496429
R27830 VSS.n4830 VSS.n4808 0.00496429
R27831 VSS.n4833 VSS.n4806 0.00496429
R27832 VSS.n4806 VSS.n4788 0.00496429
R27833 VSS.n4892 VSS.n4757 0.00496429
R27834 VSS.n4895 VSS.n4739 0.00496429
R27835 VSS.n2504 VSS.n2503 0.00496429
R27836 VSS.n2372 VSS.n2369 0.00496429
R27837 VSS.n5309 VSS.n2539 0.00496429
R27838 VSS.n5305 VSS.n2542 0.00496429
R27839 VSS.n5281 VSS.n2565 0.00496429
R27840 VSS.n5278 VSS.n2565 0.00496429
R27841 VSS.n5275 VSS.n2571 0.00496429
R27842 VSS.n5200 VSS.n5199 0.00496429
R27843 VSS.n2745 VSS.n2744 0.00496429
R27844 VSS.n5201 VSS.n2766 0.00496429
R27845 VSS.n2451 VSS.n2429 0.00496429
R27846 VSS.n2454 VSS.n2427 0.00496429
R27847 VSS.n2427 VSS.n2409 0.00496429
R27848 VSS.n2513 VSS.n2378 0.00496429
R27849 VSS.n2516 VSS.n2360 0.00496429
R27850 VSS.n5465 VSS.n5464 0.00496429
R27851 VSS.n5333 VSS.n5330 0.00496429
R27852 VSS.n5882 VSS.n5500 0.00496429
R27853 VSS.n5878 VSS.n5503 0.00496429
R27854 VSS.n5854 VSS.n5526 0.00496429
R27855 VSS.n5851 VSS.n5526 0.00496429
R27856 VSS.n5848 VSS.n5532 0.00496429
R27857 VSS.n5773 VSS.n5772 0.00496429
R27858 VSS.n5706 VSS.n5705 0.00496429
R27859 VSS.n5774 VSS.n5727 0.00496429
R27860 VSS.n5412 VSS.n5390 0.00496429
R27861 VSS.n5415 VSS.n5388 0.00496429
R27862 VSS.n5388 VSS.n5370 0.00496429
R27863 VSS.n5474 VSS.n5339 0.00496429
R27864 VSS.n5477 VSS.n5321 0.00496429
R27865 VSS.n6038 VSS.n6037 0.00496429
R27866 VSS.n5906 VSS.n5903 0.00496429
R27867 VSS.n6474 VSS.n6073 0.00496429
R27868 VSS.n6470 VSS.n6076 0.00496429
R27869 VSS.n6446 VSS.n6099 0.00496429
R27870 VSS.n6443 VSS.n6099 0.00496429
R27871 VSS.n6440 VSS.n6105 0.00496429
R27872 VSS.n6365 VSS.n6364 0.00496429
R27873 VSS.n6279 VSS.n6278 0.00496429
R27874 VSS.n6366 VSS.n6300 0.00496429
R27875 VSS.n5985 VSS.n5963 0.00496429
R27876 VSS.n5988 VSS.n5961 0.00496429
R27877 VSS.n5961 VSS.n5943 0.00496429
R27878 VSS.n6047 VSS.n5912 0.00496429
R27879 VSS.n6050 VSS.n5894 0.00496429
R27880 VSS.n7840 VSS.n7839 0.00496429
R27881 VSS.n7708 VSS.n7705 0.00496429
R27882 VSS.n7885 VSS.n7685 0.00496429
R27883 VSS.n7888 VSS.n7683 0.00496429
R27884 VSS.n7648 VSS.n7633 0.00496429
R27885 VSS.n7956 VSS.n7633 0.00496429
R27886 VSS.n7959 VSS.n7621 0.00496429
R27887 VSS.n8109 VSS.n7560 0.00496429
R27888 VSS.n8055 VSS.n8054 0.00496429
R27889 VSS.n8110 VSS.n7562 0.00496429
R27890 VSS.n7787 VSS.n7765 0.00496429
R27891 VSS.n7790 VSS.n7763 0.00496429
R27892 VSS.n7763 VSS.n7745 0.00496429
R27893 VSS.n7849 VSS.n7714 0.00496429
R27894 VSS.n7852 VSS.n7696 0.00496429
R27895 VSS.n8432 VSS.n8431 0.00496429
R27896 VSS.n8300 VSS.n8297 0.00496429
R27897 VSS.n8477 VSS.n8277 0.00496429
R27898 VSS.n8480 VSS.n8275 0.00496429
R27899 VSS.n8240 VSS.n8225 0.00496429
R27900 VSS.n8548 VSS.n8225 0.00496429
R27901 VSS.n8551 VSS.n8213 0.00496429
R27902 VSS.n8701 VSS.n8152 0.00496429
R27903 VSS.n8647 VSS.n8646 0.00496429
R27904 VSS.n8702 VSS.n8154 0.00496429
R27905 VSS.n8379 VSS.n8357 0.00496429
R27906 VSS.n8382 VSS.n8355 0.00496429
R27907 VSS.n8355 VSS.n8337 0.00496429
R27908 VSS.n8441 VSS.n8306 0.00496429
R27909 VSS.n8444 VSS.n8288 0.00496429
R27910 VSS.n9024 VSS.n9023 0.00496429
R27911 VSS.n8892 VSS.n8889 0.00496429
R27912 VSS.n9069 VSS.n8869 0.00496429
R27913 VSS.n9072 VSS.n8867 0.00496429
R27914 VSS.n8832 VSS.n8817 0.00496429
R27915 VSS.n9140 VSS.n8817 0.00496429
R27916 VSS.n9143 VSS.n8805 0.00496429
R27917 VSS.n9293 VSS.n8744 0.00496429
R27918 VSS.n9239 VSS.n9238 0.00496429
R27919 VSS.n9294 VSS.n8746 0.00496429
R27920 VSS.n8971 VSS.n8949 0.00496429
R27921 VSS.n8974 VSS.n8947 0.00496429
R27922 VSS.n8947 VSS.n8929 0.00496429
R27923 VSS.n9033 VSS.n8898 0.00496429
R27924 VSS.n9036 VSS.n8880 0.00496429
R27925 VSS.n10208 VSS.n10207 0.00496429
R27926 VSS.n10076 VSS.n10073 0.00496429
R27927 VSS.n10253 VSS.n10053 0.00496429
R27928 VSS.n10256 VSS.n10051 0.00496429
R27929 VSS.n10016 VSS.n10001 0.00496429
R27930 VSS.n10324 VSS.n10001 0.00496429
R27931 VSS.n10327 VSS.n9989 0.00496429
R27932 VSS.n10477 VSS.n9928 0.00496429
R27933 VSS.n10423 VSS.n10422 0.00496429
R27934 VSS.n10478 VSS.n9930 0.00496429
R27935 VSS.n10155 VSS.n10133 0.00496429
R27936 VSS.n10158 VSS.n10131 0.00496429
R27937 VSS.n10131 VSS.n10113 0.00496429
R27938 VSS.n10217 VSS.n10082 0.00496429
R27939 VSS.n10220 VSS.n10064 0.00496429
R27940 VSS.n10800 VSS.n10799 0.00496429
R27941 VSS.n10668 VSS.n10665 0.00496429
R27942 VSS.n10845 VSS.n10645 0.00496429
R27943 VSS.n10848 VSS.n10643 0.00496429
R27944 VSS.n10608 VSS.n10593 0.00496429
R27945 VSS.n10916 VSS.n10593 0.00496429
R27946 VSS.n10919 VSS.n10581 0.00496429
R27947 VSS.n11069 VSS.n10520 0.00496429
R27948 VSS.n11015 VSS.n11014 0.00496429
R27949 VSS.n11070 VSS.n10522 0.00496429
R27950 VSS.n10747 VSS.n10725 0.00496429
R27951 VSS.n10750 VSS.n10723 0.00496429
R27952 VSS.n10723 VSS.n10705 0.00496429
R27953 VSS.n10809 VSS.n10674 0.00496429
R27954 VSS.n10812 VSS.n10656 0.00496429
R27955 VSS.n11392 VSS.n11391 0.00496429
R27956 VSS.n11260 VSS.n11257 0.00496429
R27957 VSS.n11437 VSS.n11237 0.00496429
R27958 VSS.n11440 VSS.n11235 0.00496429
R27959 VSS.n11200 VSS.n11185 0.00496429
R27960 VSS.n11508 VSS.n11185 0.00496429
R27961 VSS.n11511 VSS.n11173 0.00496429
R27962 VSS.n11661 VSS.n11112 0.00496429
R27963 VSS.n11607 VSS.n11606 0.00496429
R27964 VSS.n11662 VSS.n11114 0.00496429
R27965 VSS.n11339 VSS.n11317 0.00496429
R27966 VSS.n11342 VSS.n11315 0.00496429
R27967 VSS.n11315 VSS.n11297 0.00496429
R27968 VSS.n11401 VSS.n11266 0.00496429
R27969 VSS.n11404 VSS.n11248 0.00496429
R27970 VSS.n11984 VSS.n11983 0.00496429
R27971 VSS.n11852 VSS.n11849 0.00496429
R27972 VSS.n12029 VSS.n11829 0.00496429
R27973 VSS.n12032 VSS.n11827 0.00496429
R27974 VSS.n11792 VSS.n11777 0.00496429
R27975 VSS.n12100 VSS.n11777 0.00496429
R27976 VSS.n12103 VSS.n11765 0.00496429
R27977 VSS.n12253 VSS.n11704 0.00496429
R27978 VSS.n12199 VSS.n12198 0.00496429
R27979 VSS.n12254 VSS.n11706 0.00496429
R27980 VSS.n11931 VSS.n11909 0.00496429
R27981 VSS.n11934 VSS.n11907 0.00496429
R27982 VSS.n11907 VSS.n11889 0.00496429
R27983 VSS.n11993 VSS.n11858 0.00496429
R27984 VSS.n11996 VSS.n11840 0.00496429
R27985 VSS.n12576 VSS.n12575 0.00496429
R27986 VSS.n12444 VSS.n12441 0.00496429
R27987 VSS.n12621 VSS.n12421 0.00496429
R27988 VSS.n12624 VSS.n12419 0.00496429
R27989 VSS.n12384 VSS.n12369 0.00496429
R27990 VSS.n12692 VSS.n12369 0.00496429
R27991 VSS.n12695 VSS.n12357 0.00496429
R27992 VSS.n12845 VSS.n12296 0.00496429
R27993 VSS.n12791 VSS.n12790 0.00496429
R27994 VSS.n12846 VSS.n12298 0.00496429
R27995 VSS.n12523 VSS.n12501 0.00496429
R27996 VSS.n12526 VSS.n12499 0.00496429
R27997 VSS.n12499 VSS.n12481 0.00496429
R27998 VSS.n12585 VSS.n12450 0.00496429
R27999 VSS.n12588 VSS.n12432 0.00496429
R28000 VSS.n13168 VSS.n13167 0.00496429
R28001 VSS.n13036 VSS.n13033 0.00496429
R28002 VSS.n13213 VSS.n13013 0.00496429
R28003 VSS.n13216 VSS.n13011 0.00496429
R28004 VSS.n12976 VSS.n12961 0.00496429
R28005 VSS.n13284 VSS.n12961 0.00496429
R28006 VSS.n13287 VSS.n12949 0.00496429
R28007 VSS.n13437 VSS.n12888 0.00496429
R28008 VSS.n13383 VSS.n13382 0.00496429
R28009 VSS.n13438 VSS.n12890 0.00496429
R28010 VSS.n13115 VSS.n13093 0.00496429
R28011 VSS.n13118 VSS.n13091 0.00496429
R28012 VSS.n13091 VSS.n13073 0.00496429
R28013 VSS.n13177 VSS.n13042 0.00496429
R28014 VSS.n13180 VSS.n13024 0.00496429
R28015 VSS.n13760 VSS.n13759 0.00496429
R28016 VSS.n13628 VSS.n13625 0.00496429
R28017 VSS.n13805 VSS.n13605 0.00496429
R28018 VSS.n13808 VSS.n13603 0.00496429
R28019 VSS.n13568 VSS.n13553 0.00496429
R28020 VSS.n13876 VSS.n13553 0.00496429
R28021 VSS.n13879 VSS.n13541 0.00496429
R28022 VSS.n14029 VSS.n13480 0.00496429
R28023 VSS.n13975 VSS.n13974 0.00496429
R28024 VSS.n14030 VSS.n13482 0.00496429
R28025 VSS.n13707 VSS.n13685 0.00496429
R28026 VSS.n13710 VSS.n13683 0.00496429
R28027 VSS.n13683 VSS.n13665 0.00496429
R28028 VSS.n13769 VSS.n13634 0.00496429
R28029 VSS.n13772 VSS.n13616 0.00496429
R28030 VSS.n14352 VSS.n14351 0.00496429
R28031 VSS.n14220 VSS.n14217 0.00496429
R28032 VSS.n14397 VSS.n14197 0.00496429
R28033 VSS.n14400 VSS.n14195 0.00496429
R28034 VSS.n14160 VSS.n14145 0.00496429
R28035 VSS.n14468 VSS.n14145 0.00496429
R28036 VSS.n14471 VSS.n14133 0.00496429
R28037 VSS.n14621 VSS.n14072 0.00496429
R28038 VSS.n14567 VSS.n14566 0.00496429
R28039 VSS.n14622 VSS.n14074 0.00496429
R28040 VSS.n14299 VSS.n14277 0.00496429
R28041 VSS.n14302 VSS.n14275 0.00496429
R28042 VSS.n14275 VSS.n14257 0.00496429
R28043 VSS.n14361 VSS.n14226 0.00496429
R28044 VSS.n14364 VSS.n14208 0.00496429
R28045 VSS.n14944 VSS.n14943 0.00496429
R28046 VSS.n14812 VSS.n14809 0.00496429
R28047 VSS.n14989 VSS.n14789 0.00496429
R28048 VSS.n14992 VSS.n14787 0.00496429
R28049 VSS.n14752 VSS.n14737 0.00496429
R28050 VSS.n15060 VSS.n14737 0.00496429
R28051 VSS.n15063 VSS.n14725 0.00496429
R28052 VSS.n15213 VSS.n14664 0.00496429
R28053 VSS.n15159 VSS.n15158 0.00496429
R28054 VSS.n15214 VSS.n14666 0.00496429
R28055 VSS.n14891 VSS.n14869 0.00496429
R28056 VSS.n14894 VSS.n14867 0.00496429
R28057 VSS.n14867 VSS.n14849 0.00496429
R28058 VSS.n14953 VSS.n14818 0.00496429
R28059 VSS.n14956 VSS.n14800 0.00496429
R28060 VSS.n15536 VSS.n15535 0.00496429
R28061 VSS.n15404 VSS.n15401 0.00496429
R28062 VSS.n15581 VSS.n15381 0.00496429
R28063 VSS.n15584 VSS.n15379 0.00496429
R28064 VSS.n15344 VSS.n15329 0.00496429
R28065 VSS.n15652 VSS.n15329 0.00496429
R28066 VSS.n15655 VSS.n15317 0.00496429
R28067 VSS.n15805 VSS.n15256 0.00496429
R28068 VSS.n15751 VSS.n15750 0.00496429
R28069 VSS.n15806 VSS.n15258 0.00496429
R28070 VSS.n15483 VSS.n15461 0.00496429
R28071 VSS.n15486 VSS.n15459 0.00496429
R28072 VSS.n15459 VSS.n15441 0.00496429
R28073 VSS.n15545 VSS.n15410 0.00496429
R28074 VSS.n15548 VSS.n15392 0.00496429
R28075 VSS.n6644 VSS.n6643 0.00496429
R28076 VSS.n6512 VSS.n6509 0.00496429
R28077 VSS.n15962 VSS.n6679 0.00496429
R28078 VSS.n15958 VSS.n6682 0.00496429
R28079 VSS.n15934 VSS.n6705 0.00496429
R28080 VSS.n15931 VSS.n6705 0.00496429
R28081 VSS.n15928 VSS.n6711 0.00496429
R28082 VSS.n15853 VSS.n15852 0.00496429
R28083 VSS.n6885 VSS.n6884 0.00496429
R28084 VSS.n15854 VSS.n6906 0.00496429
R28085 VSS.n6591 VSS.n6569 0.00496429
R28086 VSS.n6594 VSS.n6567 0.00496429
R28087 VSS.n6567 VSS.n6549 0.00496429
R28088 VSS.n6653 VSS.n6518 0.00496429
R28089 VSS.n6656 VSS.n6500 0.00496429
R28090 VSS.n7247 VSS.n7127 0.00496429
R28091 VSS.n7118 VSS.n7111 0.00496429
R28092 VSS.n7293 VSS.n7092 0.00496429
R28093 VSS.n7296 VSS.n7090 0.00496429
R28094 VSS.n7055 VSS.n7040 0.00496429
R28095 VSS.n7364 VSS.n7040 0.00496429
R28096 VSS.n7367 VSS.n7028 0.00496429
R28097 VSS.n7517 VSS.n6967 0.00496429
R28098 VSS.n7463 VSS.n7462 0.00496429
R28099 VSS.n7518 VSS.n6969 0.00496429
R28100 VSS.n7188 VSS.n7167 0.00496429
R28101 VSS.n7191 VSS.n7165 0.00496429
R28102 VSS.n7165 VSS.n7155 0.00496429
R28103 VSS.n7260 VSS.n7115 0.00496429
R28104 VSS.n7263 VSS.n7103 0.00496429
R28105 VSS.n387 VSS.n333 0.00496429
R28106 VSS.n407 VSS.n406 0.00496429
R28107 VSS.n18605 VSS.n190 0.00496429
R28108 VSS.n18608 VSS.n188 0.00496429
R28109 VSS.n153 VSS.n138 0.00496429
R28110 VSS.n18676 VSS.n138 0.00496429
R28111 VSS.n18679 VSS.n126 0.00496429
R28112 VSS.n18829 VSS.n65 0.00496429
R28113 VSS.n18775 VSS.n18774 0.00496429
R28114 VSS.n18830 VSS.n67 0.00496429
R28115 VSS.n448 VSS.n293 0.00496429
R28116 VSS.n444 VSS.n296 0.00496429
R28117 VSS.n441 VSS.n296 0.00496429
R28118 VSS.n417 VSS.n320 0.00496429
R28119 VSS.n414 VSS.n194 0.00496429
R28120 VSS.n875 VSS.n496 0.00496429
R28121 VSS.n872 VSS.n502 0.00496429
R28122 VSS.n848 VSS.n525 0.00496429
R28123 VSS.n845 VSS.n525 0.00496429
R28124 VSS.n842 VSS.n531 0.00496429
R28125 VSS.n767 VSS.n766 0.00496429
R28126 VSS.n708 VSS.n707 0.00496429
R28127 VSS.n768 VSS.n729 0.00496429
R28128 VSS.n1013 VSS.n459 0.00496429
R28129 VSS.n1009 VSS.n462 0.00496429
R28130 VSS.n1006 VSS.n462 0.00496429
R28131 VSS.n982 VSS.n486 0.00496429
R28132 VSS.n979 VSS.n492 0.00496429
R28133 VSS.n17881 VSS.n17880 0.00496429
R28134 VSS.n1367 VSS.n1366 0.00496429
R28135 VSS.n17882 VSS.n1388 0.00496429
R28136 VSS.n18029 VSS.n1033 0.00486429
R28137 VSS.n18022 VSS.n1041 0.00486429
R28138 VSS.n18021 VSS.n1042 0.00486429
R28139 VSS.n18014 VSS.n1050 0.00486429
R28140 VSS.n17042 VSS.n17041 0.00486429
R28141 VSS.n17059 VSS.n16966 0.00486429
R28142 VSS.n17061 VSS.n17060 0.00486429
R28143 VSS.n17068 VSS.n16961 0.00486429
R28144 VSS.n17539 VSS.n17538 0.00486429
R28145 VSS.n17546 VSS.n17466 0.00486429
R28146 VSS.n17550 VSS.n17549 0.00486429
R28147 VSS.n17569 VSS.n17443 0.00486429
R28148 VSS.n17634 VSS.n17633 0.00486429
R28149 VSS.n17651 VSS.n17380 0.00486429
R28150 VSS.n17653 VSS.n17652 0.00486429
R28151 VSS.n17660 VSS.n17375 0.00486429
R28152 VSS.n18116 VSS.n18115 0.00486429
R28153 VSS.n18123 VSS.n258 0.00486429
R28154 VSS.n18127 VSS.n18126 0.00486429
R28155 VSS.n18146 VSS.n235 0.00486429
R28156 VSS.n18569 VSS.n18185 0.00486429
R28157 VSS.n18562 VSS.n18193 0.00486429
R28158 VSS.n18561 VSS.n18194 0.00486429
R28159 VSS.n18554 VSS.n18201 0.00486429
R28160 VSS.n9684 VSS.n9683 0.00486429
R28161 VSS.n9701 VSS.n9430 0.00486429
R28162 VSS.n9703 VSS.n9702 0.00486429
R28163 VSS.n9710 VSS.n9425 0.00486429
R28164 VSS.n16522 VSS.n16521 0.00486429
R28165 VSS.n16539 VSS.n16447 0.00486429
R28166 VSS.n16541 VSS.n16540 0.00486429
R28167 VSS.n16548 VSS.n16442 0.00486429
R28168 VSS.n16627 VSS.n16626 0.00486429
R28169 VSS.n16644 VSS.n16372 0.00486429
R28170 VSS.n16646 VSS.n16645 0.00486429
R28171 VSS.n16653 VSS.n16367 0.00486429
R28172 VSS.n1687 VSS.n1686 0.00486429
R28173 VSS.n1704 VSS.n1612 0.00486429
R28174 VSS.n1706 VSS.n1705 0.00486429
R28175 VSS.n1713 VSS.n1607 0.00486429
R28176 VSS.n16034 VSS.n16033 0.00486429
R28177 VSS.n16051 VSS.n1544 0.00486429
R28178 VSS.n16053 VSS.n16052 0.00486429
R28179 VSS.n16060 VSS.n1539 0.00486429
R28180 VSS.n1881 VSS.n1880 0.00486429
R28181 VSS.n1888 VSS.n1808 0.00486429
R28182 VSS.n1892 VSS.n1891 0.00486429
R28183 VSS.n1911 VSS.n1785 0.00486429
R28184 VSS.n2334 VSS.n1950 0.00486429
R28185 VSS.n2327 VSS.n1958 0.00486429
R28186 VSS.n2326 VSS.n1959 0.00486429
R28187 VSS.n2319 VSS.n1966 0.00486429
R28188 VSS.n3080 VSS.n3079 0.00486429
R28189 VSS.n3087 VSS.n3007 0.00486429
R28190 VSS.n3091 VSS.n3090 0.00486429
R28191 VSS.n3110 VSS.n2984 0.00486429
R28192 VSS.n3175 VSS.n3174 0.00486429
R28193 VSS.n3192 VSS.n2921 0.00486429
R28194 VSS.n3194 VSS.n3193 0.00486429
R28195 VSS.n3201 VSS.n2916 0.00486429
R28196 VSS.n3672 VSS.n3671 0.00486429
R28197 VSS.n3679 VSS.n3599 0.00486429
R28198 VSS.n3683 VSS.n3682 0.00486429
R28199 VSS.n3702 VSS.n3576 0.00486429
R28200 VSS.n3767 VSS.n3766 0.00486429
R28201 VSS.n3784 VSS.n3513 0.00486429
R28202 VSS.n3786 VSS.n3785 0.00486429
R28203 VSS.n3793 VSS.n3508 0.00486429
R28204 VSS.n4264 VSS.n4263 0.00486429
R28205 VSS.n4271 VSS.n4191 0.00486429
R28206 VSS.n4275 VSS.n4274 0.00486429
R28207 VSS.n4294 VSS.n4168 0.00486429
R28208 VSS.n4359 VSS.n4358 0.00486429
R28209 VSS.n4376 VSS.n4105 0.00486429
R28210 VSS.n4378 VSS.n4377 0.00486429
R28211 VSS.n4385 VSS.n4100 0.00486429
R28212 VSS.n4856 VSS.n4855 0.00486429
R28213 VSS.n4863 VSS.n4783 0.00486429
R28214 VSS.n4867 VSS.n4866 0.00486429
R28215 VSS.n4886 VSS.n4760 0.00486429
R28216 VSS.n4951 VSS.n4950 0.00486429
R28217 VSS.n4968 VSS.n4697 0.00486429
R28218 VSS.n4970 VSS.n4969 0.00486429
R28219 VSS.n4977 VSS.n4692 0.00486429
R28220 VSS.n2477 VSS.n2476 0.00486429
R28221 VSS.n2484 VSS.n2404 0.00486429
R28222 VSS.n2488 VSS.n2487 0.00486429
R28223 VSS.n2507 VSS.n2381 0.00486429
R28224 VSS.n5299 VSS.n2546 0.00486429
R28225 VSS.n5292 VSS.n2554 0.00486429
R28226 VSS.n5291 VSS.n2555 0.00486429
R28227 VSS.n5284 VSS.n2562 0.00486429
R28228 VSS.n5438 VSS.n5437 0.00486429
R28229 VSS.n5445 VSS.n5365 0.00486429
R28230 VSS.n5449 VSS.n5448 0.00486429
R28231 VSS.n5468 VSS.n5342 0.00486429
R28232 VSS.n5872 VSS.n5507 0.00486429
R28233 VSS.n5865 VSS.n5515 0.00486429
R28234 VSS.n5864 VSS.n5516 0.00486429
R28235 VSS.n5857 VSS.n5523 0.00486429
R28236 VSS.n6011 VSS.n6010 0.00486429
R28237 VSS.n6018 VSS.n5938 0.00486429
R28238 VSS.n6022 VSS.n6021 0.00486429
R28239 VSS.n6041 VSS.n5915 0.00486429
R28240 VSS.n6464 VSS.n6080 0.00486429
R28241 VSS.n6457 VSS.n6088 0.00486429
R28242 VSS.n6456 VSS.n6089 0.00486429
R28243 VSS.n6449 VSS.n6096 0.00486429
R28244 VSS.n7813 VSS.n7812 0.00486429
R28245 VSS.n7820 VSS.n7740 0.00486429
R28246 VSS.n7824 VSS.n7823 0.00486429
R28247 VSS.n7843 VSS.n7717 0.00486429
R28248 VSS.n7908 VSS.n7907 0.00486429
R28249 VSS.n7925 VSS.n7654 0.00486429
R28250 VSS.n7927 VSS.n7926 0.00486429
R28251 VSS.n7934 VSS.n7649 0.00486429
R28252 VSS.n8405 VSS.n8404 0.00486429
R28253 VSS.n8412 VSS.n8332 0.00486429
R28254 VSS.n8416 VSS.n8415 0.00486429
R28255 VSS.n8435 VSS.n8309 0.00486429
R28256 VSS.n8500 VSS.n8499 0.00486429
R28257 VSS.n8517 VSS.n8246 0.00486429
R28258 VSS.n8519 VSS.n8518 0.00486429
R28259 VSS.n8526 VSS.n8241 0.00486429
R28260 VSS.n8997 VSS.n8996 0.00486429
R28261 VSS.n9004 VSS.n8924 0.00486429
R28262 VSS.n9008 VSS.n9007 0.00486429
R28263 VSS.n9027 VSS.n8901 0.00486429
R28264 VSS.n9092 VSS.n9091 0.00486429
R28265 VSS.n9109 VSS.n8838 0.00486429
R28266 VSS.n9111 VSS.n9110 0.00486429
R28267 VSS.n9118 VSS.n8833 0.00486429
R28268 VSS.n10181 VSS.n10180 0.00486429
R28269 VSS.n10188 VSS.n10108 0.00486429
R28270 VSS.n10192 VSS.n10191 0.00486429
R28271 VSS.n10211 VSS.n10085 0.00486429
R28272 VSS.n10276 VSS.n10275 0.00486429
R28273 VSS.n10293 VSS.n10022 0.00486429
R28274 VSS.n10295 VSS.n10294 0.00486429
R28275 VSS.n10302 VSS.n10017 0.00486429
R28276 VSS.n10773 VSS.n10772 0.00486429
R28277 VSS.n10780 VSS.n10700 0.00486429
R28278 VSS.n10784 VSS.n10783 0.00486429
R28279 VSS.n10803 VSS.n10677 0.00486429
R28280 VSS.n10868 VSS.n10867 0.00486429
R28281 VSS.n10885 VSS.n10614 0.00486429
R28282 VSS.n10887 VSS.n10886 0.00486429
R28283 VSS.n10894 VSS.n10609 0.00486429
R28284 VSS.n11365 VSS.n11364 0.00486429
R28285 VSS.n11372 VSS.n11292 0.00486429
R28286 VSS.n11376 VSS.n11375 0.00486429
R28287 VSS.n11395 VSS.n11269 0.00486429
R28288 VSS.n11460 VSS.n11459 0.00486429
R28289 VSS.n11477 VSS.n11206 0.00486429
R28290 VSS.n11479 VSS.n11478 0.00486429
R28291 VSS.n11486 VSS.n11201 0.00486429
R28292 VSS.n11957 VSS.n11956 0.00486429
R28293 VSS.n11964 VSS.n11884 0.00486429
R28294 VSS.n11968 VSS.n11967 0.00486429
R28295 VSS.n11987 VSS.n11861 0.00486429
R28296 VSS.n12052 VSS.n12051 0.00486429
R28297 VSS.n12069 VSS.n11798 0.00486429
R28298 VSS.n12071 VSS.n12070 0.00486429
R28299 VSS.n12078 VSS.n11793 0.00486429
R28300 VSS.n12549 VSS.n12548 0.00486429
R28301 VSS.n12556 VSS.n12476 0.00486429
R28302 VSS.n12560 VSS.n12559 0.00486429
R28303 VSS.n12579 VSS.n12453 0.00486429
R28304 VSS.n12644 VSS.n12643 0.00486429
R28305 VSS.n12661 VSS.n12390 0.00486429
R28306 VSS.n12663 VSS.n12662 0.00486429
R28307 VSS.n12670 VSS.n12385 0.00486429
R28308 VSS.n13141 VSS.n13140 0.00486429
R28309 VSS.n13148 VSS.n13068 0.00486429
R28310 VSS.n13152 VSS.n13151 0.00486429
R28311 VSS.n13171 VSS.n13045 0.00486429
R28312 VSS.n13236 VSS.n13235 0.00486429
R28313 VSS.n13253 VSS.n12982 0.00486429
R28314 VSS.n13255 VSS.n13254 0.00486429
R28315 VSS.n13262 VSS.n12977 0.00486429
R28316 VSS.n13733 VSS.n13732 0.00486429
R28317 VSS.n13740 VSS.n13660 0.00486429
R28318 VSS.n13744 VSS.n13743 0.00486429
R28319 VSS.n13763 VSS.n13637 0.00486429
R28320 VSS.n13828 VSS.n13827 0.00486429
R28321 VSS.n13845 VSS.n13574 0.00486429
R28322 VSS.n13847 VSS.n13846 0.00486429
R28323 VSS.n13854 VSS.n13569 0.00486429
R28324 VSS.n14325 VSS.n14324 0.00486429
R28325 VSS.n14332 VSS.n14252 0.00486429
R28326 VSS.n14336 VSS.n14335 0.00486429
R28327 VSS.n14355 VSS.n14229 0.00486429
R28328 VSS.n14420 VSS.n14419 0.00486429
R28329 VSS.n14437 VSS.n14166 0.00486429
R28330 VSS.n14439 VSS.n14438 0.00486429
R28331 VSS.n14446 VSS.n14161 0.00486429
R28332 VSS.n14917 VSS.n14916 0.00486429
R28333 VSS.n14924 VSS.n14844 0.00486429
R28334 VSS.n14928 VSS.n14927 0.00486429
R28335 VSS.n14947 VSS.n14821 0.00486429
R28336 VSS.n15012 VSS.n15011 0.00486429
R28337 VSS.n15029 VSS.n14758 0.00486429
R28338 VSS.n15031 VSS.n15030 0.00486429
R28339 VSS.n15038 VSS.n14753 0.00486429
R28340 VSS.n15509 VSS.n15508 0.00486429
R28341 VSS.n15516 VSS.n15436 0.00486429
R28342 VSS.n15520 VSS.n15519 0.00486429
R28343 VSS.n15539 VSS.n15413 0.00486429
R28344 VSS.n15604 VSS.n15603 0.00486429
R28345 VSS.n15621 VSS.n15350 0.00486429
R28346 VSS.n15623 VSS.n15622 0.00486429
R28347 VSS.n15630 VSS.n15345 0.00486429
R28348 VSS.n6617 VSS.n6616 0.00486429
R28349 VSS.n6624 VSS.n6544 0.00486429
R28350 VSS.n6628 VSS.n6627 0.00486429
R28351 VSS.n6647 VSS.n6521 0.00486429
R28352 VSS.n15952 VSS.n6686 0.00486429
R28353 VSS.n15945 VSS.n6694 0.00486429
R28354 VSS.n15944 VSS.n6695 0.00486429
R28355 VSS.n15937 VSS.n6702 0.00486429
R28356 VSS.n7211 VSS.n7210 0.00486429
R28357 VSS.n7228 VSS.n7136 0.00486429
R28358 VSS.n7230 VSS.n7229 0.00486429
R28359 VSS.n7237 VSS.n7131 0.00486429
R28360 VSS.n7316 VSS.n7315 0.00486429
R28361 VSS.n7333 VSS.n7061 0.00486429
R28362 VSS.n7335 VSS.n7334 0.00486429
R28363 VSS.n7342 VSS.n7056 0.00486429
R28364 VSS.n438 VSS.n300 0.00486429
R28365 VSS.n431 VSS.n308 0.00486429
R28366 VSS.n430 VSS.n309 0.00486429
R28367 VSS.n423 VSS.n317 0.00486429
R28368 VSS.n18628 VSS.n18627 0.00486429
R28369 VSS.n18645 VSS.n159 0.00486429
R28370 VSS.n18647 VSS.n18646 0.00486429
R28371 VSS.n18654 VSS.n154 0.00486429
R28372 VSS.n1003 VSS.n466 0.00486429
R28373 VSS.n996 VSS.n474 0.00486429
R28374 VSS.n995 VSS.n475 0.00486429
R28375 VSS.n988 VSS.n483 0.00486429
R28376 VSS.n866 VSS.n506 0.00486429
R28377 VSS.n859 VSS.n514 0.00486429
R28378 VSS.n858 VSS.n515 0.00486429
R28379 VSS.n851 VSS.n522 0.00486429
R28380 VSS.n17980 VSS.n1168 0.00486429
R28381 VSS.n17973 VSS.n1176 0.00486429
R28382 VSS.n17972 VSS.n1177 0.00486429
R28383 VSS.n17965 VSS.n1184 0.00486429
R28384 VSS.n9589 VSS.n9588 0.00483333
R28385 VSS.n9596 VSS.n9516 0.00483333
R28386 VSS.n9600 VSS.n9599 0.00483333
R28387 VSS.n9619 VSS.n9493 0.00483333
R28388 VSS.n17272 VSS 0.00452857
R28389 VSS.n17864 VSS 0.00452857
R28390 VSS.n18429 VSS 0.00452857
R28391 VSS.n9915 VSS 0.00452857
R28392 VSS.n16858 VSS 0.00452857
R28393 VSS.n16265 VSS 0.00452857
R28394 VSS.n2220 VSS 0.00452857
R28395 VSS.n3406 VSS 0.00452857
R28396 VSS.n3998 VSS 0.00452857
R28397 VSS.n4590 VSS 0.00452857
R28398 VSS.n5182 VSS 0.00452857
R28399 VSS.n5185 VSS 0.00452857
R28400 VSS.n18888 VSS 0.00452857
R28401 VSS.n6350 VSS 0.00452857
R28402 VSS.n8139 VSS 0.00452857
R28403 VSS.n8731 VSS 0.00452857
R28404 VSS.n9323 VSS 0.00452857
R28405 VSS.n10507 VSS 0.00452857
R28406 VSS.n11099 VSS 0.00452857
R28407 VSS.n11691 VSS 0.00452857
R28408 VSS.n12283 VSS 0.00452857
R28409 VSS.n12875 VSS 0.00452857
R28410 VSS.n13467 VSS 0.00452857
R28411 VSS.n14059 VSS 0.00452857
R28412 VSS.n14651 VSS 0.00452857
R28413 VSS.n15243 VSS 0.00452857
R28414 VSS.n15835 VSS 0.00452857
R28415 VSS.n15838 VSS 0.00452857
R28416 VSS.n7547 VSS 0.00452857
R28417 VSS.n18859 VSS 0.00452857
R28418 VSS.n18861 VSS 0.00452857
R28419 VSS.n17866 VSS 0.00452857
R28420 VSS.n924 VSS.n464 0.00407143
R28421 VSS.n1105 VSS.n1031 0.00407143
R28422 VSS.n17108 VSS.n16930 0.00407143
R28423 VSS.n17149 VSS.n16924 0.00407143
R28424 VSS.n17155 VSS.n17154 0.00407143
R28425 VSS.n17269 VSS.n16863 0.00407143
R28426 VSS.n17148 VSS.n17147 0.00407143
R28427 VSS.n17156 VSS.n16920 0.00407143
R28428 VSS.n17210 VSS.n17209 0.00407143
R28429 VSS.n17486 VSS.n17473 0.00407143
R28430 VSS.n17700 VSS.n17344 0.00407143
R28431 VSS.n17741 VSS.n17338 0.00407143
R28432 VSS.n17747 VSS.n17746 0.00407143
R28433 VSS.n17861 VSS.n17277 0.00407143
R28434 VSS.n17740 VSS.n17739 0.00407143
R28435 VSS.n17748 VSS.n17334 0.00407143
R28436 VSS.n17802 VSS.n17801 0.00407143
R28437 VSS.n278 VSS.n265 0.00407143
R28438 VSS.n18325 VSS.n18323 0.00407143
R28439 VSS.n18525 VSS.n18316 0.00407143
R28440 VSS.n18518 VSS.n18517 0.00407143
R28441 VSS.n18465 VSS.n18434 0.00407143
R28442 VSS.n18524 VSS.n18523 0.00407143
R28443 VSS.n18519 VSS.n18338 0.00407143
R28444 VSS.n18400 VSS.n18399 0.00407143
R28445 VSS.n9536 VSS.n9523 0.00407143
R28446 VSS.n9750 VSS.n9394 0.00407143
R28447 VSS.n9791 VSS.n9388 0.00407143
R28448 VSS.n9797 VSS.n9796 0.00407143
R28449 VSS.n9912 VSS.n9328 0.00407143
R28450 VSS.n9790 VSS.n9789 0.00407143
R28451 VSS.n9798 VSS.n9384 0.00407143
R28452 VSS.n9852 VSS.n9851 0.00407143
R28453 VSS.n16514 VSS.n16467 0.00407143
R28454 VSS.n16693 VSS.n16336 0.00407143
R28455 VSS.n16734 VSS.n16330 0.00407143
R28456 VSS.n16740 VSS.n16739 0.00407143
R28457 VSS.n16855 VSS.n16270 0.00407143
R28458 VSS.n16733 VSS.n16732 0.00407143
R28459 VSS.n16741 VSS.n16326 0.00407143
R28460 VSS.n16795 VSS.n16794 0.00407143
R28461 VSS.n1679 VSS.n1632 0.00407143
R28462 VSS.n16100 VSS.n1508 0.00407143
R28463 VSS.n16141 VSS.n1502 0.00407143
R28464 VSS.n16147 VSS.n16146 0.00407143
R28465 VSS.n16262 VSS.n1442 0.00407143
R28466 VSS.n16140 VSS.n16139 0.00407143
R28467 VSS.n16148 VSS.n1498 0.00407143
R28468 VSS.n16202 VSS.n16201 0.00407143
R28469 VSS.n1828 VSS.n1815 0.00407143
R28470 VSS.n2089 VSS.n2087 0.00407143
R28471 VSS.n2287 VSS.n2080 0.00407143
R28472 VSS.n2115 VSS.n2114 0.00407143
R28473 VSS.n2224 VSS.n2223 0.00407143
R28474 VSS.n2289 VSS.n2288 0.00407143
R28475 VSS.n2116 VSS.n2113 0.00407143
R28476 VSS.n2258 VSS.n2257 0.00407143
R28477 VSS.n3027 VSS.n3014 0.00407143
R28478 VSS.n3241 VSS.n2885 0.00407143
R28479 VSS.n3282 VSS.n2879 0.00407143
R28480 VSS.n3288 VSS.n3287 0.00407143
R28481 VSS.n3403 VSS.n2819 0.00407143
R28482 VSS.n3281 VSS.n3280 0.00407143
R28483 VSS.n3289 VSS.n2875 0.00407143
R28484 VSS.n3343 VSS.n3342 0.00407143
R28485 VSS.n3619 VSS.n3606 0.00407143
R28486 VSS.n3833 VSS.n3477 0.00407143
R28487 VSS.n3874 VSS.n3471 0.00407143
R28488 VSS.n3880 VSS.n3879 0.00407143
R28489 VSS.n3995 VSS.n3411 0.00407143
R28490 VSS.n3873 VSS.n3872 0.00407143
R28491 VSS.n3881 VSS.n3467 0.00407143
R28492 VSS.n3935 VSS.n3934 0.00407143
R28493 VSS.n4211 VSS.n4198 0.00407143
R28494 VSS.n4425 VSS.n4069 0.00407143
R28495 VSS.n4466 VSS.n4063 0.00407143
R28496 VSS.n4472 VSS.n4471 0.00407143
R28497 VSS.n4587 VSS.n4003 0.00407143
R28498 VSS.n4465 VSS.n4464 0.00407143
R28499 VSS.n4473 VSS.n4059 0.00407143
R28500 VSS.n4527 VSS.n4526 0.00407143
R28501 VSS.n4803 VSS.n4790 0.00407143
R28502 VSS.n5017 VSS.n4661 0.00407143
R28503 VSS.n5058 VSS.n4655 0.00407143
R28504 VSS.n5064 VSS.n5063 0.00407143
R28505 VSS.n5179 VSS.n4595 0.00407143
R28506 VSS.n5057 VSS.n5056 0.00407143
R28507 VSS.n5065 VSS.n4651 0.00407143
R28508 VSS.n5119 VSS.n5118 0.00407143
R28509 VSS.n2424 VSS.n2411 0.00407143
R28510 VSS.n2685 VSS.n2683 0.00407143
R28511 VSS.n5252 VSS.n2676 0.00407143
R28512 VSS.n2711 VSS.n2710 0.00407143
R28513 VSS.n5189 VSS.n5188 0.00407143
R28514 VSS.n5254 VSS.n5253 0.00407143
R28515 VSS.n2712 VSS.n2709 0.00407143
R28516 VSS.n5223 VSS.n5222 0.00407143
R28517 VSS.n5385 VSS.n5372 0.00407143
R28518 VSS.n5646 VSS.n5644 0.00407143
R28519 VSS.n5825 VSS.n5637 0.00407143
R28520 VSS.n5672 VSS.n5671 0.00407143
R28521 VSS.n18885 VSS.n4 0.00407143
R28522 VSS.n5827 VSS.n5826 0.00407143
R28523 VSS.n5673 VSS.n5670 0.00407143
R28524 VSS.n5796 VSS.n5795 0.00407143
R28525 VSS.n5958 VSS.n5945 0.00407143
R28526 VSS.n6219 VSS.n6217 0.00407143
R28527 VSS.n6417 VSS.n6210 0.00407143
R28528 VSS.n6245 VSS.n6244 0.00407143
R28529 VSS.n6354 VSS.n6353 0.00407143
R28530 VSS.n6419 VSS.n6418 0.00407143
R28531 VSS.n6246 VSS.n6243 0.00407143
R28532 VSS.n6388 VSS.n6387 0.00407143
R28533 VSS.n7760 VSS.n7747 0.00407143
R28534 VSS.n7974 VSS.n7618 0.00407143
R28535 VSS.n8015 VSS.n7612 0.00407143
R28536 VSS.n8021 VSS.n8020 0.00407143
R28537 VSS.n8136 VSS.n7552 0.00407143
R28538 VSS.n8014 VSS.n8013 0.00407143
R28539 VSS.n8022 VSS.n7608 0.00407143
R28540 VSS.n8076 VSS.n8075 0.00407143
R28541 VSS.n8352 VSS.n8339 0.00407143
R28542 VSS.n8566 VSS.n8210 0.00407143
R28543 VSS.n8607 VSS.n8204 0.00407143
R28544 VSS.n8613 VSS.n8612 0.00407143
R28545 VSS.n8728 VSS.n8144 0.00407143
R28546 VSS.n8606 VSS.n8605 0.00407143
R28547 VSS.n8614 VSS.n8200 0.00407143
R28548 VSS.n8668 VSS.n8667 0.00407143
R28549 VSS.n8944 VSS.n8931 0.00407143
R28550 VSS.n9158 VSS.n8802 0.00407143
R28551 VSS.n9199 VSS.n8796 0.00407143
R28552 VSS.n9205 VSS.n9204 0.00407143
R28553 VSS.n9320 VSS.n8736 0.00407143
R28554 VSS.n9198 VSS.n9197 0.00407143
R28555 VSS.n9206 VSS.n8792 0.00407143
R28556 VSS.n9260 VSS.n9259 0.00407143
R28557 VSS.n10128 VSS.n10115 0.00407143
R28558 VSS.n10342 VSS.n9986 0.00407143
R28559 VSS.n10383 VSS.n9980 0.00407143
R28560 VSS.n10389 VSS.n10388 0.00407143
R28561 VSS.n10504 VSS.n9920 0.00407143
R28562 VSS.n10382 VSS.n10381 0.00407143
R28563 VSS.n10390 VSS.n9976 0.00407143
R28564 VSS.n10444 VSS.n10443 0.00407143
R28565 VSS.n10720 VSS.n10707 0.00407143
R28566 VSS.n10934 VSS.n10578 0.00407143
R28567 VSS.n10975 VSS.n10572 0.00407143
R28568 VSS.n10981 VSS.n10980 0.00407143
R28569 VSS.n11096 VSS.n10512 0.00407143
R28570 VSS.n10974 VSS.n10973 0.00407143
R28571 VSS.n10982 VSS.n10568 0.00407143
R28572 VSS.n11036 VSS.n11035 0.00407143
R28573 VSS.n11312 VSS.n11299 0.00407143
R28574 VSS.n11526 VSS.n11170 0.00407143
R28575 VSS.n11567 VSS.n11164 0.00407143
R28576 VSS.n11573 VSS.n11572 0.00407143
R28577 VSS.n11688 VSS.n11104 0.00407143
R28578 VSS.n11566 VSS.n11565 0.00407143
R28579 VSS.n11574 VSS.n11160 0.00407143
R28580 VSS.n11628 VSS.n11627 0.00407143
R28581 VSS.n11904 VSS.n11891 0.00407143
R28582 VSS.n12118 VSS.n11762 0.00407143
R28583 VSS.n12159 VSS.n11756 0.00407143
R28584 VSS.n12165 VSS.n12164 0.00407143
R28585 VSS.n12280 VSS.n11696 0.00407143
R28586 VSS.n12158 VSS.n12157 0.00407143
R28587 VSS.n12166 VSS.n11752 0.00407143
R28588 VSS.n12220 VSS.n12219 0.00407143
R28589 VSS.n12496 VSS.n12483 0.00407143
R28590 VSS.n12710 VSS.n12354 0.00407143
R28591 VSS.n12751 VSS.n12348 0.00407143
R28592 VSS.n12757 VSS.n12756 0.00407143
R28593 VSS.n12872 VSS.n12288 0.00407143
R28594 VSS.n12750 VSS.n12749 0.00407143
R28595 VSS.n12758 VSS.n12344 0.00407143
R28596 VSS.n12812 VSS.n12811 0.00407143
R28597 VSS.n13088 VSS.n13075 0.00407143
R28598 VSS.n13302 VSS.n12946 0.00407143
R28599 VSS.n13343 VSS.n12940 0.00407143
R28600 VSS.n13349 VSS.n13348 0.00407143
R28601 VSS.n13464 VSS.n12880 0.00407143
R28602 VSS.n13342 VSS.n13341 0.00407143
R28603 VSS.n13350 VSS.n12936 0.00407143
R28604 VSS.n13404 VSS.n13403 0.00407143
R28605 VSS.n13680 VSS.n13667 0.00407143
R28606 VSS.n13894 VSS.n13538 0.00407143
R28607 VSS.n13935 VSS.n13532 0.00407143
R28608 VSS.n13941 VSS.n13940 0.00407143
R28609 VSS.n14056 VSS.n13472 0.00407143
R28610 VSS.n13934 VSS.n13933 0.00407143
R28611 VSS.n13942 VSS.n13528 0.00407143
R28612 VSS.n13996 VSS.n13995 0.00407143
R28613 VSS.n14272 VSS.n14259 0.00407143
R28614 VSS.n14486 VSS.n14130 0.00407143
R28615 VSS.n14527 VSS.n14124 0.00407143
R28616 VSS.n14533 VSS.n14532 0.00407143
R28617 VSS.n14648 VSS.n14064 0.00407143
R28618 VSS.n14526 VSS.n14525 0.00407143
R28619 VSS.n14534 VSS.n14120 0.00407143
R28620 VSS.n14588 VSS.n14587 0.00407143
R28621 VSS.n14864 VSS.n14851 0.00407143
R28622 VSS.n15078 VSS.n14722 0.00407143
R28623 VSS.n15119 VSS.n14716 0.00407143
R28624 VSS.n15125 VSS.n15124 0.00407143
R28625 VSS.n15240 VSS.n14656 0.00407143
R28626 VSS.n15118 VSS.n15117 0.00407143
R28627 VSS.n15126 VSS.n14712 0.00407143
R28628 VSS.n15180 VSS.n15179 0.00407143
R28629 VSS.n15456 VSS.n15443 0.00407143
R28630 VSS.n15670 VSS.n15314 0.00407143
R28631 VSS.n15711 VSS.n15308 0.00407143
R28632 VSS.n15717 VSS.n15716 0.00407143
R28633 VSS.n15832 VSS.n15248 0.00407143
R28634 VSS.n15710 VSS.n15709 0.00407143
R28635 VSS.n15718 VSS.n15304 0.00407143
R28636 VSS.n15772 VSS.n15771 0.00407143
R28637 VSS.n6564 VSS.n6551 0.00407143
R28638 VSS.n6825 VSS.n6823 0.00407143
R28639 VSS.n15905 VSS.n6816 0.00407143
R28640 VSS.n6851 VSS.n6850 0.00407143
R28641 VSS.n15842 VSS.n15841 0.00407143
R28642 VSS.n15907 VSS.n15906 0.00407143
R28643 VSS.n6852 VSS.n6849 0.00407143
R28644 VSS.n15876 VSS.n15875 0.00407143
R28645 VSS.n7203 VSS.n7156 0.00407143
R28646 VSS.n7382 VSS.n7025 0.00407143
R28647 VSS.n7423 VSS.n7019 0.00407143
R28648 VSS.n7429 VSS.n7428 0.00407143
R28649 VSS.n7544 VSS.n6959 0.00407143
R28650 VSS.n7422 VSS.n7421 0.00407143
R28651 VSS.n7430 VSS.n7015 0.00407143
R28652 VSS.n7484 VSS.n7483 0.00407143
R28653 VSS.n366 VSS.n298 0.00407143
R28654 VSS.n18694 VSS.n123 0.00407143
R28655 VSS.n18735 VSS.n117 0.00407143
R28656 VSS.n18741 VSS.n18740 0.00407143
R28657 VSS.n18856 VSS.n57 0.00407143
R28658 VSS.n18734 VSS.n18733 0.00407143
R28659 VSS.n18742 VSS.n113 0.00407143
R28660 VSS.n18796 VSS.n18795 0.00407143
R28661 VSS.n648 VSS.n646 0.00407143
R28662 VSS.n819 VSS.n639 0.00407143
R28663 VSS.n674 VSS.n673 0.00407143
R28664 VSS.n18865 VSS.n18864 0.00407143
R28665 VSS.n821 VSS.n820 0.00407143
R28666 VSS.n675 VSS.n672 0.00407143
R28667 VSS.n790 VSS.n789 0.00407143
R28668 VSS.n1307 VSS.n1305 0.00407143
R28669 VSS.n17933 VSS.n1298 0.00407143
R28670 VSS.n1333 VSS.n1332 0.00407143
R28671 VSS.n17870 VSS.n17869 0.00407143
R28672 VSS.n17935 VSS.n17934 0.00407143
R28673 VSS.n1334 VSS.n1331 0.00407143
R28674 VSS.n17904 VSS.n17903 0.00407143
R28675 VSS.n17135 VSS.n17134 0.00352143
R28676 VSS.n17144 VSS.n16927 0.00352143
R28677 VSS.n17175 VSS.n17174 0.00352143
R28678 VSS.n17176 VSS.n16901 0.00352143
R28679 VSS.n17207 VSS.n17192 0.00352143
R28680 VSS.n17226 VSS.n16887 0.00352143
R28681 VSS.n17247 VSS.n17246 0.00352143
R28682 VSS.n17271 VSS.n16860 0.00352143
R28683 VSS.n17727 VSS.n17726 0.00352143
R28684 VSS.n17736 VSS.n17341 0.00352143
R28685 VSS.n17767 VSS.n17766 0.00352143
R28686 VSS.n17768 VSS.n17315 0.00352143
R28687 VSS.n17799 VSS.n17784 0.00352143
R28688 VSS.n17818 VSS.n17301 0.00352143
R28689 VSS.n17839 VSS.n17838 0.00352143
R28690 VSS.n17863 VSS.n17274 0.00352143
R28691 VSS.n18329 VSS.n18328 0.00352143
R28692 VSS.n18336 VSS.n18318 0.00352143
R28693 VSS.n18350 VSS.n18337 0.00352143
R28694 VSS.n18504 VSS.n18351 0.00352143
R28695 VSS.n18413 VSS.n18392 0.00352143
R28696 VSS.n18486 VSS.n18414 0.00352143
R28697 VSS.n18470 VSS.n18469 0.00352143
R28698 VSS.n18468 VSS.n18430 0.00352143
R28699 VSS.n9777 VSS.n9776 0.00352143
R28700 VSS.n9786 VSS.n9391 0.00352143
R28701 VSS.n9817 VSS.n9816 0.00352143
R28702 VSS.n9818 VSS.n9365 0.00352143
R28703 VSS.n9849 VSS.n9834 0.00352143
R28704 VSS.n9868 VSS.n9351 0.00352143
R28705 VSS.n9889 VSS.n9888 0.00352143
R28706 VSS.n9914 VSS.n9325 0.00352143
R28707 VSS.n16720 VSS.n16719 0.00352143
R28708 VSS.n16729 VSS.n16333 0.00352143
R28709 VSS.n16760 VSS.n16759 0.00352143
R28710 VSS.n16761 VSS.n16307 0.00352143
R28711 VSS.n16792 VSS.n16777 0.00352143
R28712 VSS.n16811 VSS.n16293 0.00352143
R28713 VSS.n16832 VSS.n16831 0.00352143
R28714 VSS.n16857 VSS.n16267 0.00352143
R28715 VSS.n16127 VSS.n16126 0.00352143
R28716 VSS.n16136 VSS.n1505 0.00352143
R28717 VSS.n16167 VSS.n16166 0.00352143
R28718 VSS.n16168 VSS.n1479 0.00352143
R28719 VSS.n16199 VSS.n16184 0.00352143
R28720 VSS.n16218 VSS.n1465 0.00352143
R28721 VSS.n16239 VSS.n16238 0.00352143
R28722 VSS.n16264 VSS.n1439 0.00352143
R28723 VSS.n2093 VSS.n2092 0.00352143
R28724 VSS.n2100 VSS.n2083 0.00352143
R28725 VSS.n2135 VSS.n2118 0.00352143
R28726 VSS.n2136 VSS.n2131 0.00352143
R28727 VSS.n2255 VSS.n2152 0.00352143
R28728 VSS.n2168 VSS.n2167 0.00352143
R28729 VSS.n2218 VSS.n2169 0.00352143
R28730 VSS.n2221 VSS.n2219 0.00352143
R28731 VSS.n3268 VSS.n3267 0.00352143
R28732 VSS.n3277 VSS.n2882 0.00352143
R28733 VSS.n3308 VSS.n3307 0.00352143
R28734 VSS.n3309 VSS.n2856 0.00352143
R28735 VSS.n3340 VSS.n3325 0.00352143
R28736 VSS.n3359 VSS.n2842 0.00352143
R28737 VSS.n3380 VSS.n3379 0.00352143
R28738 VSS.n3405 VSS.n2816 0.00352143
R28739 VSS.n3860 VSS.n3859 0.00352143
R28740 VSS.n3869 VSS.n3474 0.00352143
R28741 VSS.n3900 VSS.n3899 0.00352143
R28742 VSS.n3901 VSS.n3448 0.00352143
R28743 VSS.n3932 VSS.n3917 0.00352143
R28744 VSS.n3951 VSS.n3434 0.00352143
R28745 VSS.n3972 VSS.n3971 0.00352143
R28746 VSS.n3997 VSS.n3408 0.00352143
R28747 VSS.n4452 VSS.n4451 0.00352143
R28748 VSS.n4461 VSS.n4066 0.00352143
R28749 VSS.n4492 VSS.n4491 0.00352143
R28750 VSS.n4493 VSS.n4040 0.00352143
R28751 VSS.n4524 VSS.n4509 0.00352143
R28752 VSS.n4543 VSS.n4026 0.00352143
R28753 VSS.n4564 VSS.n4563 0.00352143
R28754 VSS.n4589 VSS.n4000 0.00352143
R28755 VSS.n5044 VSS.n5043 0.00352143
R28756 VSS.n5053 VSS.n4658 0.00352143
R28757 VSS.n5084 VSS.n5083 0.00352143
R28758 VSS.n5085 VSS.n4632 0.00352143
R28759 VSS.n5116 VSS.n5101 0.00352143
R28760 VSS.n5135 VSS.n4618 0.00352143
R28761 VSS.n5156 VSS.n5155 0.00352143
R28762 VSS.n5181 VSS.n4592 0.00352143
R28763 VSS.n2689 VSS.n2688 0.00352143
R28764 VSS.n2696 VSS.n2679 0.00352143
R28765 VSS.n2731 VSS.n2714 0.00352143
R28766 VSS.n2732 VSS.n2727 0.00352143
R28767 VSS.n5220 VSS.n2748 0.00352143
R28768 VSS.n2764 VSS.n2763 0.00352143
R28769 VSS.n2814 VSS.n2765 0.00352143
R28770 VSS.n5186 VSS.n2815 0.00352143
R28771 VSS.n5650 VSS.n5649 0.00352143
R28772 VSS.n5657 VSS.n5640 0.00352143
R28773 VSS.n5692 VSS.n5675 0.00352143
R28774 VSS.n5693 VSS.n5688 0.00352143
R28775 VSS.n5793 VSS.n5709 0.00352143
R28776 VSS.n5725 VSS.n5724 0.00352143
R28777 VSS.n5731 VSS.n5726 0.00352143
R28778 VSS.n18887 VSS.n1 0.00352143
R28779 VSS.n6223 VSS.n6222 0.00352143
R28780 VSS.n6230 VSS.n6213 0.00352143
R28781 VSS.n6265 VSS.n6248 0.00352143
R28782 VSS.n6266 VSS.n6261 0.00352143
R28783 VSS.n6385 VSS.n6282 0.00352143
R28784 VSS.n6298 VSS.n6297 0.00352143
R28785 VSS.n6348 VSS.n6299 0.00352143
R28786 VSS.n6351 VSS.n6349 0.00352143
R28787 VSS.n8001 VSS.n8000 0.00352143
R28788 VSS.n8010 VSS.n7615 0.00352143
R28789 VSS.n8041 VSS.n8040 0.00352143
R28790 VSS.n8042 VSS.n7589 0.00352143
R28791 VSS.n8073 VSS.n8058 0.00352143
R28792 VSS.n8092 VSS.n7575 0.00352143
R28793 VSS.n8113 VSS.n8112 0.00352143
R28794 VSS.n8138 VSS.n7549 0.00352143
R28795 VSS.n8593 VSS.n8592 0.00352143
R28796 VSS.n8602 VSS.n8207 0.00352143
R28797 VSS.n8633 VSS.n8632 0.00352143
R28798 VSS.n8634 VSS.n8181 0.00352143
R28799 VSS.n8665 VSS.n8650 0.00352143
R28800 VSS.n8684 VSS.n8167 0.00352143
R28801 VSS.n8705 VSS.n8704 0.00352143
R28802 VSS.n8730 VSS.n8141 0.00352143
R28803 VSS.n9185 VSS.n9184 0.00352143
R28804 VSS.n9194 VSS.n8799 0.00352143
R28805 VSS.n9225 VSS.n9224 0.00352143
R28806 VSS.n9226 VSS.n8773 0.00352143
R28807 VSS.n9257 VSS.n9242 0.00352143
R28808 VSS.n9276 VSS.n8759 0.00352143
R28809 VSS.n9297 VSS.n9296 0.00352143
R28810 VSS.n9322 VSS.n8733 0.00352143
R28811 VSS.n10369 VSS.n10368 0.00352143
R28812 VSS.n10378 VSS.n9983 0.00352143
R28813 VSS.n10409 VSS.n10408 0.00352143
R28814 VSS.n10410 VSS.n9957 0.00352143
R28815 VSS.n10441 VSS.n10426 0.00352143
R28816 VSS.n10460 VSS.n9943 0.00352143
R28817 VSS.n10481 VSS.n10480 0.00352143
R28818 VSS.n10506 VSS.n9917 0.00352143
R28819 VSS.n10961 VSS.n10960 0.00352143
R28820 VSS.n10970 VSS.n10575 0.00352143
R28821 VSS.n11001 VSS.n11000 0.00352143
R28822 VSS.n11002 VSS.n10549 0.00352143
R28823 VSS.n11033 VSS.n11018 0.00352143
R28824 VSS.n11052 VSS.n10535 0.00352143
R28825 VSS.n11073 VSS.n11072 0.00352143
R28826 VSS.n11098 VSS.n10509 0.00352143
R28827 VSS.n11553 VSS.n11552 0.00352143
R28828 VSS.n11562 VSS.n11167 0.00352143
R28829 VSS.n11593 VSS.n11592 0.00352143
R28830 VSS.n11594 VSS.n11141 0.00352143
R28831 VSS.n11625 VSS.n11610 0.00352143
R28832 VSS.n11644 VSS.n11127 0.00352143
R28833 VSS.n11665 VSS.n11664 0.00352143
R28834 VSS.n11690 VSS.n11101 0.00352143
R28835 VSS.n12145 VSS.n12144 0.00352143
R28836 VSS.n12154 VSS.n11759 0.00352143
R28837 VSS.n12185 VSS.n12184 0.00352143
R28838 VSS.n12186 VSS.n11733 0.00352143
R28839 VSS.n12217 VSS.n12202 0.00352143
R28840 VSS.n12236 VSS.n11719 0.00352143
R28841 VSS.n12257 VSS.n12256 0.00352143
R28842 VSS.n12282 VSS.n11693 0.00352143
R28843 VSS.n12737 VSS.n12736 0.00352143
R28844 VSS.n12746 VSS.n12351 0.00352143
R28845 VSS.n12777 VSS.n12776 0.00352143
R28846 VSS.n12778 VSS.n12325 0.00352143
R28847 VSS.n12809 VSS.n12794 0.00352143
R28848 VSS.n12828 VSS.n12311 0.00352143
R28849 VSS.n12849 VSS.n12848 0.00352143
R28850 VSS.n12874 VSS.n12285 0.00352143
R28851 VSS.n13329 VSS.n13328 0.00352143
R28852 VSS.n13338 VSS.n12943 0.00352143
R28853 VSS.n13369 VSS.n13368 0.00352143
R28854 VSS.n13370 VSS.n12917 0.00352143
R28855 VSS.n13401 VSS.n13386 0.00352143
R28856 VSS.n13420 VSS.n12903 0.00352143
R28857 VSS.n13441 VSS.n13440 0.00352143
R28858 VSS.n13466 VSS.n12877 0.00352143
R28859 VSS.n13921 VSS.n13920 0.00352143
R28860 VSS.n13930 VSS.n13535 0.00352143
R28861 VSS.n13961 VSS.n13960 0.00352143
R28862 VSS.n13962 VSS.n13509 0.00352143
R28863 VSS.n13993 VSS.n13978 0.00352143
R28864 VSS.n14012 VSS.n13495 0.00352143
R28865 VSS.n14033 VSS.n14032 0.00352143
R28866 VSS.n14058 VSS.n13469 0.00352143
R28867 VSS.n14513 VSS.n14512 0.00352143
R28868 VSS.n14522 VSS.n14127 0.00352143
R28869 VSS.n14553 VSS.n14552 0.00352143
R28870 VSS.n14554 VSS.n14101 0.00352143
R28871 VSS.n14585 VSS.n14570 0.00352143
R28872 VSS.n14604 VSS.n14087 0.00352143
R28873 VSS.n14625 VSS.n14624 0.00352143
R28874 VSS.n14650 VSS.n14061 0.00352143
R28875 VSS.n15105 VSS.n15104 0.00352143
R28876 VSS.n15114 VSS.n14719 0.00352143
R28877 VSS.n15145 VSS.n15144 0.00352143
R28878 VSS.n15146 VSS.n14693 0.00352143
R28879 VSS.n15177 VSS.n15162 0.00352143
R28880 VSS.n15196 VSS.n14679 0.00352143
R28881 VSS.n15217 VSS.n15216 0.00352143
R28882 VSS.n15242 VSS.n14653 0.00352143
R28883 VSS.n15697 VSS.n15696 0.00352143
R28884 VSS.n15706 VSS.n15311 0.00352143
R28885 VSS.n15737 VSS.n15736 0.00352143
R28886 VSS.n15738 VSS.n15285 0.00352143
R28887 VSS.n15769 VSS.n15754 0.00352143
R28888 VSS.n15788 VSS.n15271 0.00352143
R28889 VSS.n15809 VSS.n15808 0.00352143
R28890 VSS.n15834 VSS.n15245 0.00352143
R28891 VSS.n6829 VSS.n6828 0.00352143
R28892 VSS.n6836 VSS.n6819 0.00352143
R28893 VSS.n6871 VSS.n6854 0.00352143
R28894 VSS.n6872 VSS.n6867 0.00352143
R28895 VSS.n15873 VSS.n6888 0.00352143
R28896 VSS.n6904 VSS.n6903 0.00352143
R28897 VSS.n6954 VSS.n6905 0.00352143
R28898 VSS.n15839 VSS.n6955 0.00352143
R28899 VSS.n7409 VSS.n7408 0.00352143
R28900 VSS.n7418 VSS.n7022 0.00352143
R28901 VSS.n7449 VSS.n7448 0.00352143
R28902 VSS.n7450 VSS.n6996 0.00352143
R28903 VSS.n7481 VSS.n7466 0.00352143
R28904 VSS.n7500 VSS.n6982 0.00352143
R28905 VSS.n7521 VSS.n7520 0.00352143
R28906 VSS.n7546 VSS.n6956 0.00352143
R28907 VSS.n18721 VSS.n18720 0.00352143
R28908 VSS.n18730 VSS.n120 0.00352143
R28909 VSS.n18761 VSS.n18760 0.00352143
R28910 VSS.n18762 VSS.n94 0.00352143
R28911 VSS.n18793 VSS.n18778 0.00352143
R28912 VSS.n18812 VSS.n80 0.00352143
R28913 VSS.n18833 VSS.n18832 0.00352143
R28914 VSS.n18858 VSS.n54 0.00352143
R28915 VSS.n652 VSS.n651 0.00352143
R28916 VSS.n659 VSS.n642 0.00352143
R28917 VSS.n694 VSS.n677 0.00352143
R28918 VSS.n695 VSS.n690 0.00352143
R28919 VSS.n787 VSS.n711 0.00352143
R28920 VSS.n727 VSS.n726 0.00352143
R28921 VSS.n733 VSS.n728 0.00352143
R28922 VSS.n18862 VSS.n52 0.00352143
R28923 VSS.n1311 VSS.n1310 0.00352143
R28924 VSS.n1318 VSS.n1301 0.00352143
R28925 VSS.n1353 VSS.n1336 0.00352143
R28926 VSS.n1354 VSS.n1349 0.00352143
R28927 VSS.n17901 VSS.n1370 0.00352143
R28928 VSS.n1386 VSS.n1385 0.00352143
R28929 VSS.n1436 VSS.n1387 0.00352143
R28930 VSS.n17867 VSS.n1437 0.00352143
R28931 VSS.n1041 VSS.n1033 0.00318571
R28932 VSS.n1050 VSS.n1042 0.00318571
R28933 VSS.n17041 VSS.n16966 0.00318571
R28934 VSS.n17061 VSS.n16961 0.00318571
R28935 VSS.n17539 VSS.n17466 0.00318571
R28936 VSS.n17549 VSS.n17443 0.00318571
R28937 VSS.n17633 VSS.n17380 0.00318571
R28938 VSS.n17653 VSS.n17375 0.00318571
R28939 VSS.n18116 VSS.n258 0.00318571
R28940 VSS.n18126 VSS.n235 0.00318571
R28941 VSS.n18193 VSS.n18185 0.00318571
R28942 VSS.n18201 VSS.n18194 0.00318571
R28943 VSS.n9683 VSS.n9430 0.00318571
R28944 VSS.n9703 VSS.n9425 0.00318571
R28945 VSS.n16521 VSS.n16447 0.00318571
R28946 VSS.n16541 VSS.n16442 0.00318571
R28947 VSS.n16626 VSS.n16372 0.00318571
R28948 VSS.n16646 VSS.n16367 0.00318571
R28949 VSS.n1686 VSS.n1612 0.00318571
R28950 VSS.n1706 VSS.n1607 0.00318571
R28951 VSS.n16033 VSS.n1544 0.00318571
R28952 VSS.n16053 VSS.n1539 0.00318571
R28953 VSS.n1881 VSS.n1808 0.00318571
R28954 VSS.n1891 VSS.n1785 0.00318571
R28955 VSS.n1958 VSS.n1950 0.00318571
R28956 VSS.n1966 VSS.n1959 0.00318571
R28957 VSS.n3080 VSS.n3007 0.00318571
R28958 VSS.n3090 VSS.n2984 0.00318571
R28959 VSS.n3174 VSS.n2921 0.00318571
R28960 VSS.n3194 VSS.n2916 0.00318571
R28961 VSS.n3672 VSS.n3599 0.00318571
R28962 VSS.n3682 VSS.n3576 0.00318571
R28963 VSS.n3766 VSS.n3513 0.00318571
R28964 VSS.n3786 VSS.n3508 0.00318571
R28965 VSS.n4264 VSS.n4191 0.00318571
R28966 VSS.n4274 VSS.n4168 0.00318571
R28967 VSS.n4358 VSS.n4105 0.00318571
R28968 VSS.n4378 VSS.n4100 0.00318571
R28969 VSS.n4856 VSS.n4783 0.00318571
R28970 VSS.n4866 VSS.n4760 0.00318571
R28971 VSS.n4950 VSS.n4697 0.00318571
R28972 VSS.n4970 VSS.n4692 0.00318571
R28973 VSS.n2477 VSS.n2404 0.00318571
R28974 VSS.n2487 VSS.n2381 0.00318571
R28975 VSS.n2554 VSS.n2546 0.00318571
R28976 VSS.n2562 VSS.n2555 0.00318571
R28977 VSS.n5438 VSS.n5365 0.00318571
R28978 VSS.n5448 VSS.n5342 0.00318571
R28979 VSS.n5515 VSS.n5507 0.00318571
R28980 VSS.n5523 VSS.n5516 0.00318571
R28981 VSS.n6011 VSS.n5938 0.00318571
R28982 VSS.n6021 VSS.n5915 0.00318571
R28983 VSS.n6088 VSS.n6080 0.00318571
R28984 VSS.n6096 VSS.n6089 0.00318571
R28985 VSS.n7813 VSS.n7740 0.00318571
R28986 VSS.n7823 VSS.n7717 0.00318571
R28987 VSS.n7907 VSS.n7654 0.00318571
R28988 VSS.n7927 VSS.n7649 0.00318571
R28989 VSS.n8405 VSS.n8332 0.00318571
R28990 VSS.n8415 VSS.n8309 0.00318571
R28991 VSS.n8499 VSS.n8246 0.00318571
R28992 VSS.n8519 VSS.n8241 0.00318571
R28993 VSS.n8997 VSS.n8924 0.00318571
R28994 VSS.n9007 VSS.n8901 0.00318571
R28995 VSS.n9091 VSS.n8838 0.00318571
R28996 VSS.n9111 VSS.n8833 0.00318571
R28997 VSS.n10181 VSS.n10108 0.00318571
R28998 VSS.n10191 VSS.n10085 0.00318571
R28999 VSS.n10275 VSS.n10022 0.00318571
R29000 VSS.n10295 VSS.n10017 0.00318571
R29001 VSS.n10773 VSS.n10700 0.00318571
R29002 VSS.n10783 VSS.n10677 0.00318571
R29003 VSS.n10867 VSS.n10614 0.00318571
R29004 VSS.n10887 VSS.n10609 0.00318571
R29005 VSS.n11365 VSS.n11292 0.00318571
R29006 VSS.n11375 VSS.n11269 0.00318571
R29007 VSS.n11459 VSS.n11206 0.00318571
R29008 VSS.n11479 VSS.n11201 0.00318571
R29009 VSS.n11957 VSS.n11884 0.00318571
R29010 VSS.n11967 VSS.n11861 0.00318571
R29011 VSS.n12051 VSS.n11798 0.00318571
R29012 VSS.n12071 VSS.n11793 0.00318571
R29013 VSS.n12549 VSS.n12476 0.00318571
R29014 VSS.n12559 VSS.n12453 0.00318571
R29015 VSS.n12643 VSS.n12390 0.00318571
R29016 VSS.n12663 VSS.n12385 0.00318571
R29017 VSS.n13141 VSS.n13068 0.00318571
R29018 VSS.n13151 VSS.n13045 0.00318571
R29019 VSS.n13235 VSS.n12982 0.00318571
R29020 VSS.n13255 VSS.n12977 0.00318571
R29021 VSS.n13733 VSS.n13660 0.00318571
R29022 VSS.n13743 VSS.n13637 0.00318571
R29023 VSS.n13827 VSS.n13574 0.00318571
R29024 VSS.n13847 VSS.n13569 0.00318571
R29025 VSS.n14325 VSS.n14252 0.00318571
R29026 VSS.n14335 VSS.n14229 0.00318571
R29027 VSS.n14419 VSS.n14166 0.00318571
R29028 VSS.n14439 VSS.n14161 0.00318571
R29029 VSS.n14917 VSS.n14844 0.00318571
R29030 VSS.n14927 VSS.n14821 0.00318571
R29031 VSS.n15011 VSS.n14758 0.00318571
R29032 VSS.n15031 VSS.n14753 0.00318571
R29033 VSS.n15509 VSS.n15436 0.00318571
R29034 VSS.n15519 VSS.n15413 0.00318571
R29035 VSS.n15603 VSS.n15350 0.00318571
R29036 VSS.n15623 VSS.n15345 0.00318571
R29037 VSS.n6617 VSS.n6544 0.00318571
R29038 VSS.n6627 VSS.n6521 0.00318571
R29039 VSS.n6694 VSS.n6686 0.00318571
R29040 VSS.n6702 VSS.n6695 0.00318571
R29041 VSS.n7210 VSS.n7136 0.00318571
R29042 VSS.n7230 VSS.n7131 0.00318571
R29043 VSS.n7315 VSS.n7061 0.00318571
R29044 VSS.n7335 VSS.n7056 0.00318571
R29045 VSS.n308 VSS.n300 0.00318571
R29046 VSS.n317 VSS.n309 0.00318571
R29047 VSS.n18627 VSS.n159 0.00318571
R29048 VSS.n18647 VSS.n154 0.00318571
R29049 VSS.n474 VSS.n466 0.00318571
R29050 VSS.n483 VSS.n475 0.00318571
R29051 VSS.n514 VSS.n506 0.00318571
R29052 VSS.n522 VSS.n515 0.00318571
R29053 VSS.n1176 VSS.n1168 0.00318571
R29054 VSS.n1184 VSS.n1177 0.00318571
R29055 VSS.n1226 VSS.n1159 0.00317857
R29056 VSS.n17985 VSS.n1165 0.00317857
R29057 VSS.n17970 VSS.n17969 0.00317857
R29058 VSS.n1262 VSS.n1188 0.00317857
R29059 VSS.n17960 VSS.n1189 0.00317857
R29060 VSS.n17955 VSS.n1194 0.00317857
R29061 VSS.n1225 VSS.n1161 0.00317857
R29062 VSS.n17986 VSS.n1163 0.00317857
R29063 VSS.n17971 VSS.n1178 0.00317857
R29064 VSS.n17959 VSS.n1190 0.00317857
R29065 VSS.n17956 VSS.n1192 0.00317857
R29066 VSS.n912 VSS.n457 0.00317857
R29067 VSS.n1008 VSS.n463 0.00317857
R29068 VSS.n999 VSS.n470 0.00317857
R29069 VSS.n946 VSS.n487 0.00317857
R29070 VSS.n983 VSS.n488 0.00317857
R29071 VSS.n978 VSS.n493 0.00317857
R29072 VSS.n17018 VSS.n17017 0.00317857
R29073 VSS.n17024 VSS.n16994 0.00317857
R29074 VSS.n17064 VSS.n16963 0.00317857
R29075 VSS.n17073 VSS.n17072 0.00317857
R29076 VSS.n17089 VSS.n17088 0.00317857
R29077 VSS.n17094 VSS.n16934 0.00317857
R29078 VSS.n1093 VSS.n1024 0.00317857
R29079 VSS.n18034 VSS.n1030 0.00317857
R29080 VSS.n18025 VSS.n1037 0.00317857
R29081 VSS.n1127 VSS.n1054 0.00317857
R29082 VSS.n18009 VSS.n1055 0.00317857
R29083 VSS.n18004 VSS.n1060 0.00317857
R29084 VSS.n1092 VSS.n1026 0.00317857
R29085 VSS.n18035 VSS.n1028 0.00317857
R29086 VSS.n18024 VSS.n18023 0.00317857
R29087 VSS.n18008 VSS.n1056 0.00317857
R29088 VSS.n18005 VSS.n1058 0.00317857
R29089 VSS.n17109 VSS.n17108 0.00317857
R29090 VSS.n17186 VSS.n16903 0.00317857
R29091 VSS.n17198 VSS.n16898 0.00317857
R29092 VSS.n17228 VSS.n16885 0.00317857
R29093 VSS.n17251 VSS.n17250 0.00317857
R29094 VSS.n17269 VSS.n17268 0.00317857
R29095 VSS.n17230 VSS.n17229 0.00317857
R29096 VSS.n17019 VSS.n16998 0.00317857
R29097 VSS.n17023 VSS.n17022 0.00317857
R29098 VSS.n17063 VSS.n16964 0.00317857
R29099 VSS.n17090 VSS.n16946 0.00317857
R29100 VSS.n17095 VSS.n17093 0.00317857
R29101 VSS.n17610 VSS.n17609 0.00317857
R29102 VSS.n17616 VSS.n17408 0.00317857
R29103 VSS.n17656 VSS.n17377 0.00317857
R29104 VSS.n17665 VSS.n17664 0.00317857
R29105 VSS.n17681 VSS.n17680 0.00317857
R29106 VSS.n17686 VSS.n17348 0.00317857
R29107 VSS.n17512 VSS.n17511 0.00317857
R29108 VSS.n17518 VSS.n17488 0.00317857
R29109 VSS.n17543 VSS.n17461 0.00317857
R29110 VSS.n17454 VSS.n17441 0.00317857
R29111 VSS.n17574 VSS.n17430 0.00317857
R29112 VSS.n17580 VSS.n17423 0.00317857
R29113 VSS.n17513 VSS.n17492 0.00317857
R29114 VSS.n17517 VSS.n17516 0.00317857
R29115 VSS.n17545 VSS.n17544 0.00317857
R29116 VSS.n17575 VSS.n17432 0.00317857
R29117 VSS.n17579 VSS.n17578 0.00317857
R29118 VSS.n17701 VSS.n17700 0.00317857
R29119 VSS.n17778 VSS.n17317 0.00317857
R29120 VSS.n17790 VSS.n17312 0.00317857
R29121 VSS.n17820 VSS.n17299 0.00317857
R29122 VSS.n17843 VSS.n17842 0.00317857
R29123 VSS.n17861 VSS.n17860 0.00317857
R29124 VSS.n17822 VSS.n17821 0.00317857
R29125 VSS.n17611 VSS.n17412 0.00317857
R29126 VSS.n17615 VSS.n17614 0.00317857
R29127 VSS.n17655 VSS.n17378 0.00317857
R29128 VSS.n17682 VSS.n17360 0.00317857
R29129 VSS.n17687 VSS.n17685 0.00317857
R29130 VSS.n18089 VSS.n18088 0.00317857
R29131 VSS.n18095 VSS.n280 0.00317857
R29132 VSS.n18120 VSS.n253 0.00317857
R29133 VSS.n246 VSS.n233 0.00317857
R29134 VSS.n18151 VSS.n222 0.00317857
R29135 VSS.n18157 VSS.n215 0.00317857
R29136 VSS.n18243 VSS.n212 0.00317857
R29137 VSS.n18574 VSS.n18182 0.00317857
R29138 VSS.n18559 VSS.n18558 0.00317857
R29139 VSS.n18279 VSS.n18205 0.00317857
R29140 VSS.n18549 VSS.n18206 0.00317857
R29141 VSS.n18544 VSS.n18211 0.00317857
R29142 VSS.n18242 VSS.n18178 0.00317857
R29143 VSS.n18575 VSS.n18180 0.00317857
R29144 VSS.n18560 VSS.n18195 0.00317857
R29145 VSS.n18548 VSS.n18207 0.00317857
R29146 VSS.n18545 VSS.n18209 0.00317857
R29147 VSS.n18325 VSS.n18324 0.00317857
R29148 VSS.n18376 VSS.n18355 0.00317857
R29149 VSS.n18403 VSS.n18402 0.00317857
R29150 VSS.n18483 VSS.n18418 0.00317857
R29151 VSS.n18472 VSS.n18426 0.00317857
R29152 VSS.n18465 VSS.n18464 0.00317857
R29153 VSS.n18484 VSS.n18416 0.00317857
R29154 VSS.n18090 VSS.n284 0.00317857
R29155 VSS.n18094 VSS.n18093 0.00317857
R29156 VSS.n18122 VSS.n18121 0.00317857
R29157 VSS.n18152 VSS.n224 0.00317857
R29158 VSS.n18156 VSS.n18155 0.00317857
R29159 VSS.n9562 VSS.n9561 0.00317857
R29160 VSS.n9568 VSS.n9538 0.00317857
R29161 VSS.n9593 VSS.n9511 0.00317857
R29162 VSS.n9504 VSS.n9491 0.00317857
R29163 VSS.n9624 VSS.n9480 0.00317857
R29164 VSS.n9630 VSS.n9473 0.00317857
R29165 VSS.n9660 VSS.n9659 0.00317857
R29166 VSS.n9666 VSS.n9458 0.00317857
R29167 VSS.n9706 VSS.n9427 0.00317857
R29168 VSS.n9715 VSS.n9714 0.00317857
R29169 VSS.n9731 VSS.n9730 0.00317857
R29170 VSS.n9736 VSS.n9398 0.00317857
R29171 VSS.n9661 VSS.n9462 0.00317857
R29172 VSS.n9665 VSS.n9664 0.00317857
R29173 VSS.n9705 VSS.n9428 0.00317857
R29174 VSS.n9732 VSS.n9410 0.00317857
R29175 VSS.n9737 VSS.n9735 0.00317857
R29176 VSS.n9751 VSS.n9750 0.00317857
R29177 VSS.n9828 VSS.n9367 0.00317857
R29178 VSS.n9840 VSS.n9362 0.00317857
R29179 VSS.n9870 VSS.n9349 0.00317857
R29180 VSS.n9894 VSS.n9893 0.00317857
R29181 VSS.n9912 VSS.n9911 0.00317857
R29182 VSS.n9872 VSS.n9871 0.00317857
R29183 VSS.n9563 VSS.n9542 0.00317857
R29184 VSS.n9567 VSS.n9566 0.00317857
R29185 VSS.n9595 VSS.n9594 0.00317857
R29186 VSS.n9625 VSS.n9482 0.00317857
R29187 VSS.n9629 VSS.n9628 0.00317857
R29188 VSS.n16498 VSS.n16497 0.00317857
R29189 VSS.n16504 VSS.n16475 0.00317857
R29190 VSS.n16537 VSS.n16450 0.00317857
R29191 VSS.n16553 VSS.n16552 0.00317857
R29192 VSS.n16570 VSS.n16569 0.00317857
R29193 VSS.n16575 VSS.n16415 0.00317857
R29194 VSS.n16603 VSS.n16602 0.00317857
R29195 VSS.n16609 VSS.n16400 0.00317857
R29196 VSS.n16649 VSS.n16369 0.00317857
R29197 VSS.n16658 VSS.n16657 0.00317857
R29198 VSS.n16674 VSS.n16673 0.00317857
R29199 VSS.n16679 VSS.n16340 0.00317857
R29200 VSS.n16604 VSS.n16404 0.00317857
R29201 VSS.n16608 VSS.n16607 0.00317857
R29202 VSS.n16648 VSS.n16370 0.00317857
R29203 VSS.n16675 VSS.n16352 0.00317857
R29204 VSS.n16680 VSS.n16678 0.00317857
R29205 VSS.n16694 VSS.n16693 0.00317857
R29206 VSS.n16771 VSS.n16309 0.00317857
R29207 VSS.n16783 VSS.n16304 0.00317857
R29208 VSS.n16813 VSS.n16291 0.00317857
R29209 VSS.n16837 VSS.n16836 0.00317857
R29210 VSS.n16855 VSS.n16854 0.00317857
R29211 VSS.n16815 VSS.n16814 0.00317857
R29212 VSS.n16499 VSS.n16479 0.00317857
R29213 VSS.n16503 VSS.n16502 0.00317857
R29214 VSS.n16538 VSS.n16448 0.00317857
R29215 VSS.n16571 VSS.n16427 0.00317857
R29216 VSS.n16576 VSS.n16574 0.00317857
R29217 VSS.n1663 VSS.n1662 0.00317857
R29218 VSS.n1669 VSS.n1640 0.00317857
R29219 VSS.n1702 VSS.n1615 0.00317857
R29220 VSS.n1718 VSS.n1717 0.00317857
R29221 VSS.n1735 VSS.n1734 0.00317857
R29222 VSS.n1740 VSS.n1580 0.00317857
R29223 VSS.n16010 VSS.n16009 0.00317857
R29224 VSS.n16016 VSS.n1572 0.00317857
R29225 VSS.n16056 VSS.n1541 0.00317857
R29226 VSS.n16065 VSS.n16064 0.00317857
R29227 VSS.n16081 VSS.n16080 0.00317857
R29228 VSS.n16086 VSS.n1512 0.00317857
R29229 VSS.n16011 VSS.n1576 0.00317857
R29230 VSS.n16015 VSS.n16014 0.00317857
R29231 VSS.n16055 VSS.n1542 0.00317857
R29232 VSS.n16082 VSS.n1524 0.00317857
R29233 VSS.n16087 VSS.n16085 0.00317857
R29234 VSS.n16101 VSS.n16100 0.00317857
R29235 VSS.n16178 VSS.n1481 0.00317857
R29236 VSS.n16190 VSS.n1476 0.00317857
R29237 VSS.n16220 VSS.n1463 0.00317857
R29238 VSS.n16244 VSS.n16243 0.00317857
R29239 VSS.n16262 VSS.n16261 0.00317857
R29240 VSS.n16222 VSS.n16221 0.00317857
R29241 VSS.n1664 VSS.n1644 0.00317857
R29242 VSS.n1668 VSS.n1667 0.00317857
R29243 VSS.n1703 VSS.n1613 0.00317857
R29244 VSS.n1736 VSS.n1592 0.00317857
R29245 VSS.n1741 VSS.n1739 0.00317857
R29246 VSS.n1854 VSS.n1853 0.00317857
R29247 VSS.n1860 VSS.n1830 0.00317857
R29248 VSS.n1885 VSS.n1803 0.00317857
R29249 VSS.n1796 VSS.n1783 0.00317857
R29250 VSS.n1916 VSS.n1772 0.00317857
R29251 VSS.n1922 VSS.n1765 0.00317857
R29252 VSS.n2008 VSS.n1762 0.00317857
R29253 VSS.n2339 VSS.n1947 0.00317857
R29254 VSS.n2324 VSS.n2323 0.00317857
R29255 VSS.n2044 VSS.n1970 0.00317857
R29256 VSS.n2314 VSS.n1971 0.00317857
R29257 VSS.n2309 VSS.n1976 0.00317857
R29258 VSS.n2007 VSS.n1943 0.00317857
R29259 VSS.n2340 VSS.n1945 0.00317857
R29260 VSS.n2325 VSS.n1960 0.00317857
R29261 VSS.n2313 VSS.n1972 0.00317857
R29262 VSS.n2310 VSS.n1974 0.00317857
R29263 VSS.n2089 VSS.n2088 0.00317857
R29264 VSS.n2146 VSS.n2133 0.00317857
R29265 VSS.n2180 VSS.n2128 0.00317857
R29266 VSS.n2242 VSS.n2241 0.00317857
R29267 VSS.n2214 VSS.n2213 0.00317857
R29268 VSS.n2223 VSS.n2201 0.00317857
R29269 VSS.n2240 VSS.n2161 0.00317857
R29270 VSS.n1855 VSS.n1834 0.00317857
R29271 VSS.n1859 VSS.n1858 0.00317857
R29272 VSS.n1887 VSS.n1886 0.00317857
R29273 VSS.n1917 VSS.n1774 0.00317857
R29274 VSS.n1921 VSS.n1920 0.00317857
R29275 VSS.n3053 VSS.n3052 0.00317857
R29276 VSS.n3059 VSS.n3029 0.00317857
R29277 VSS.n3084 VSS.n3002 0.00317857
R29278 VSS.n2995 VSS.n2982 0.00317857
R29279 VSS.n3115 VSS.n2971 0.00317857
R29280 VSS.n3121 VSS.n2964 0.00317857
R29281 VSS.n3151 VSS.n3150 0.00317857
R29282 VSS.n3157 VSS.n2949 0.00317857
R29283 VSS.n3197 VSS.n2918 0.00317857
R29284 VSS.n3206 VSS.n3205 0.00317857
R29285 VSS.n3222 VSS.n3221 0.00317857
R29286 VSS.n3227 VSS.n2889 0.00317857
R29287 VSS.n3152 VSS.n2953 0.00317857
R29288 VSS.n3156 VSS.n3155 0.00317857
R29289 VSS.n3196 VSS.n2919 0.00317857
R29290 VSS.n3223 VSS.n2901 0.00317857
R29291 VSS.n3228 VSS.n3226 0.00317857
R29292 VSS.n3242 VSS.n3241 0.00317857
R29293 VSS.n3319 VSS.n2858 0.00317857
R29294 VSS.n3331 VSS.n2853 0.00317857
R29295 VSS.n3361 VSS.n2840 0.00317857
R29296 VSS.n3385 VSS.n3384 0.00317857
R29297 VSS.n3403 VSS.n3402 0.00317857
R29298 VSS.n3363 VSS.n3362 0.00317857
R29299 VSS.n3054 VSS.n3033 0.00317857
R29300 VSS.n3058 VSS.n3057 0.00317857
R29301 VSS.n3086 VSS.n3085 0.00317857
R29302 VSS.n3116 VSS.n2973 0.00317857
R29303 VSS.n3120 VSS.n3119 0.00317857
R29304 VSS.n3645 VSS.n3644 0.00317857
R29305 VSS.n3651 VSS.n3621 0.00317857
R29306 VSS.n3676 VSS.n3594 0.00317857
R29307 VSS.n3587 VSS.n3574 0.00317857
R29308 VSS.n3707 VSS.n3563 0.00317857
R29309 VSS.n3713 VSS.n3556 0.00317857
R29310 VSS.n3743 VSS.n3742 0.00317857
R29311 VSS.n3749 VSS.n3541 0.00317857
R29312 VSS.n3789 VSS.n3510 0.00317857
R29313 VSS.n3798 VSS.n3797 0.00317857
R29314 VSS.n3814 VSS.n3813 0.00317857
R29315 VSS.n3819 VSS.n3481 0.00317857
R29316 VSS.n3744 VSS.n3545 0.00317857
R29317 VSS.n3748 VSS.n3747 0.00317857
R29318 VSS.n3788 VSS.n3511 0.00317857
R29319 VSS.n3815 VSS.n3493 0.00317857
R29320 VSS.n3820 VSS.n3818 0.00317857
R29321 VSS.n3834 VSS.n3833 0.00317857
R29322 VSS.n3911 VSS.n3450 0.00317857
R29323 VSS.n3923 VSS.n3445 0.00317857
R29324 VSS.n3953 VSS.n3432 0.00317857
R29325 VSS.n3977 VSS.n3976 0.00317857
R29326 VSS.n3995 VSS.n3994 0.00317857
R29327 VSS.n3955 VSS.n3954 0.00317857
R29328 VSS.n3646 VSS.n3625 0.00317857
R29329 VSS.n3650 VSS.n3649 0.00317857
R29330 VSS.n3678 VSS.n3677 0.00317857
R29331 VSS.n3708 VSS.n3565 0.00317857
R29332 VSS.n3712 VSS.n3711 0.00317857
R29333 VSS.n4237 VSS.n4236 0.00317857
R29334 VSS.n4243 VSS.n4213 0.00317857
R29335 VSS.n4268 VSS.n4186 0.00317857
R29336 VSS.n4179 VSS.n4166 0.00317857
R29337 VSS.n4299 VSS.n4155 0.00317857
R29338 VSS.n4305 VSS.n4148 0.00317857
R29339 VSS.n4335 VSS.n4334 0.00317857
R29340 VSS.n4341 VSS.n4133 0.00317857
R29341 VSS.n4381 VSS.n4102 0.00317857
R29342 VSS.n4390 VSS.n4389 0.00317857
R29343 VSS.n4406 VSS.n4405 0.00317857
R29344 VSS.n4411 VSS.n4073 0.00317857
R29345 VSS.n4336 VSS.n4137 0.00317857
R29346 VSS.n4340 VSS.n4339 0.00317857
R29347 VSS.n4380 VSS.n4103 0.00317857
R29348 VSS.n4407 VSS.n4085 0.00317857
R29349 VSS.n4412 VSS.n4410 0.00317857
R29350 VSS.n4426 VSS.n4425 0.00317857
R29351 VSS.n4503 VSS.n4042 0.00317857
R29352 VSS.n4515 VSS.n4037 0.00317857
R29353 VSS.n4545 VSS.n4024 0.00317857
R29354 VSS.n4569 VSS.n4568 0.00317857
R29355 VSS.n4587 VSS.n4586 0.00317857
R29356 VSS.n4547 VSS.n4546 0.00317857
R29357 VSS.n4238 VSS.n4217 0.00317857
R29358 VSS.n4242 VSS.n4241 0.00317857
R29359 VSS.n4270 VSS.n4269 0.00317857
R29360 VSS.n4300 VSS.n4157 0.00317857
R29361 VSS.n4304 VSS.n4303 0.00317857
R29362 VSS.n4829 VSS.n4828 0.00317857
R29363 VSS.n4835 VSS.n4805 0.00317857
R29364 VSS.n4860 VSS.n4778 0.00317857
R29365 VSS.n4771 VSS.n4758 0.00317857
R29366 VSS.n4891 VSS.n4747 0.00317857
R29367 VSS.n4897 VSS.n4740 0.00317857
R29368 VSS.n4927 VSS.n4926 0.00317857
R29369 VSS.n4933 VSS.n4725 0.00317857
R29370 VSS.n4973 VSS.n4694 0.00317857
R29371 VSS.n4982 VSS.n4981 0.00317857
R29372 VSS.n4998 VSS.n4997 0.00317857
R29373 VSS.n5003 VSS.n4665 0.00317857
R29374 VSS.n4928 VSS.n4729 0.00317857
R29375 VSS.n4932 VSS.n4931 0.00317857
R29376 VSS.n4972 VSS.n4695 0.00317857
R29377 VSS.n4999 VSS.n4677 0.00317857
R29378 VSS.n5004 VSS.n5002 0.00317857
R29379 VSS.n5018 VSS.n5017 0.00317857
R29380 VSS.n5095 VSS.n4634 0.00317857
R29381 VSS.n5107 VSS.n4629 0.00317857
R29382 VSS.n5137 VSS.n4616 0.00317857
R29383 VSS.n5161 VSS.n5160 0.00317857
R29384 VSS.n5179 VSS.n5178 0.00317857
R29385 VSS.n5139 VSS.n5138 0.00317857
R29386 VSS.n4830 VSS.n4809 0.00317857
R29387 VSS.n4834 VSS.n4833 0.00317857
R29388 VSS.n4862 VSS.n4861 0.00317857
R29389 VSS.n4892 VSS.n4749 0.00317857
R29390 VSS.n4896 VSS.n4895 0.00317857
R29391 VSS.n2450 VSS.n2449 0.00317857
R29392 VSS.n2456 VSS.n2426 0.00317857
R29393 VSS.n2481 VSS.n2399 0.00317857
R29394 VSS.n2392 VSS.n2379 0.00317857
R29395 VSS.n2512 VSS.n2368 0.00317857
R29396 VSS.n2518 VSS.n2361 0.00317857
R29397 VSS.n2604 VSS.n2358 0.00317857
R29398 VSS.n5304 VSS.n2543 0.00317857
R29399 VSS.n5289 VSS.n5288 0.00317857
R29400 VSS.n2640 VSS.n2566 0.00317857
R29401 VSS.n5279 VSS.n2567 0.00317857
R29402 VSS.n5274 VSS.n2572 0.00317857
R29403 VSS.n2603 VSS.n2539 0.00317857
R29404 VSS.n5305 VSS.n2541 0.00317857
R29405 VSS.n5290 VSS.n2556 0.00317857
R29406 VSS.n5278 VSS.n2568 0.00317857
R29407 VSS.n5275 VSS.n2570 0.00317857
R29408 VSS.n2685 VSS.n2684 0.00317857
R29409 VSS.n2742 VSS.n2729 0.00317857
R29410 VSS.n2776 VSS.n2724 0.00317857
R29411 VSS.n5207 VSS.n5206 0.00317857
R29412 VSS.n2810 VSS.n2809 0.00317857
R29413 VSS.n5188 VSS.n2797 0.00317857
R29414 VSS.n5205 VSS.n2757 0.00317857
R29415 VSS.n2451 VSS.n2430 0.00317857
R29416 VSS.n2455 VSS.n2454 0.00317857
R29417 VSS.n2483 VSS.n2482 0.00317857
R29418 VSS.n2513 VSS.n2370 0.00317857
R29419 VSS.n2517 VSS.n2516 0.00317857
R29420 VSS.n5411 VSS.n5410 0.00317857
R29421 VSS.n5417 VSS.n5387 0.00317857
R29422 VSS.n5442 VSS.n5360 0.00317857
R29423 VSS.n5353 VSS.n5340 0.00317857
R29424 VSS.n5473 VSS.n5329 0.00317857
R29425 VSS.n5479 VSS.n5322 0.00317857
R29426 VSS.n5565 VSS.n5319 0.00317857
R29427 VSS.n5877 VSS.n5504 0.00317857
R29428 VSS.n5862 VSS.n5861 0.00317857
R29429 VSS.n5601 VSS.n5527 0.00317857
R29430 VSS.n5852 VSS.n5528 0.00317857
R29431 VSS.n5847 VSS.n5533 0.00317857
R29432 VSS.n5564 VSS.n5500 0.00317857
R29433 VSS.n5878 VSS.n5502 0.00317857
R29434 VSS.n5863 VSS.n5517 0.00317857
R29435 VSS.n5851 VSS.n5529 0.00317857
R29436 VSS.n5848 VSS.n5531 0.00317857
R29437 VSS.n5646 VSS.n5645 0.00317857
R29438 VSS.n5703 VSS.n5690 0.00317857
R29439 VSS.n5750 VSS.n5685 0.00317857
R29440 VSS.n5780 VSS.n5779 0.00317857
R29441 VSS.n5736 VSS.n5735 0.00317857
R29442 VSS.n18885 VSS.n18884 0.00317857
R29443 VSS.n5778 VSS.n5718 0.00317857
R29444 VSS.n5412 VSS.n5391 0.00317857
R29445 VSS.n5416 VSS.n5415 0.00317857
R29446 VSS.n5444 VSS.n5443 0.00317857
R29447 VSS.n5474 VSS.n5331 0.00317857
R29448 VSS.n5478 VSS.n5477 0.00317857
R29449 VSS.n5984 VSS.n5983 0.00317857
R29450 VSS.n5990 VSS.n5960 0.00317857
R29451 VSS.n6015 VSS.n5933 0.00317857
R29452 VSS.n5926 VSS.n5913 0.00317857
R29453 VSS.n6046 VSS.n5902 0.00317857
R29454 VSS.n6052 VSS.n5895 0.00317857
R29455 VSS.n6138 VSS.n5892 0.00317857
R29456 VSS.n6469 VSS.n6077 0.00317857
R29457 VSS.n6454 VSS.n6453 0.00317857
R29458 VSS.n6174 VSS.n6100 0.00317857
R29459 VSS.n6444 VSS.n6101 0.00317857
R29460 VSS.n6439 VSS.n6106 0.00317857
R29461 VSS.n6137 VSS.n6073 0.00317857
R29462 VSS.n6470 VSS.n6075 0.00317857
R29463 VSS.n6455 VSS.n6090 0.00317857
R29464 VSS.n6443 VSS.n6102 0.00317857
R29465 VSS.n6440 VSS.n6104 0.00317857
R29466 VSS.n6219 VSS.n6218 0.00317857
R29467 VSS.n6276 VSS.n6263 0.00317857
R29468 VSS.n6310 VSS.n6258 0.00317857
R29469 VSS.n6372 VSS.n6371 0.00317857
R29470 VSS.n6344 VSS.n6343 0.00317857
R29471 VSS.n6353 VSS.n6331 0.00317857
R29472 VSS.n6370 VSS.n6291 0.00317857
R29473 VSS.n5985 VSS.n5964 0.00317857
R29474 VSS.n5989 VSS.n5988 0.00317857
R29475 VSS.n6017 VSS.n6016 0.00317857
R29476 VSS.n6047 VSS.n5904 0.00317857
R29477 VSS.n6051 VSS.n6050 0.00317857
R29478 VSS.n7786 VSS.n7785 0.00317857
R29479 VSS.n7792 VSS.n7762 0.00317857
R29480 VSS.n7817 VSS.n7735 0.00317857
R29481 VSS.n7728 VSS.n7715 0.00317857
R29482 VSS.n7848 VSS.n7704 0.00317857
R29483 VSS.n7854 VSS.n7697 0.00317857
R29484 VSS.n7884 VSS.n7883 0.00317857
R29485 VSS.n7890 VSS.n7682 0.00317857
R29486 VSS.n7930 VSS.n7651 0.00317857
R29487 VSS.n7939 VSS.n7938 0.00317857
R29488 VSS.n7955 VSS.n7954 0.00317857
R29489 VSS.n7960 VSS.n7622 0.00317857
R29490 VSS.n7885 VSS.n7686 0.00317857
R29491 VSS.n7889 VSS.n7888 0.00317857
R29492 VSS.n7929 VSS.n7652 0.00317857
R29493 VSS.n7956 VSS.n7634 0.00317857
R29494 VSS.n7961 VSS.n7959 0.00317857
R29495 VSS.n7975 VSS.n7974 0.00317857
R29496 VSS.n8052 VSS.n7591 0.00317857
R29497 VSS.n8064 VSS.n7586 0.00317857
R29498 VSS.n8094 VSS.n7573 0.00317857
R29499 VSS.n8118 VSS.n8117 0.00317857
R29500 VSS.n8136 VSS.n8135 0.00317857
R29501 VSS.n8096 VSS.n8095 0.00317857
R29502 VSS.n7787 VSS.n7766 0.00317857
R29503 VSS.n7791 VSS.n7790 0.00317857
R29504 VSS.n7819 VSS.n7818 0.00317857
R29505 VSS.n7849 VSS.n7706 0.00317857
R29506 VSS.n7853 VSS.n7852 0.00317857
R29507 VSS.n8378 VSS.n8377 0.00317857
R29508 VSS.n8384 VSS.n8354 0.00317857
R29509 VSS.n8409 VSS.n8327 0.00317857
R29510 VSS.n8320 VSS.n8307 0.00317857
R29511 VSS.n8440 VSS.n8296 0.00317857
R29512 VSS.n8446 VSS.n8289 0.00317857
R29513 VSS.n8476 VSS.n8475 0.00317857
R29514 VSS.n8482 VSS.n8274 0.00317857
R29515 VSS.n8522 VSS.n8243 0.00317857
R29516 VSS.n8531 VSS.n8530 0.00317857
R29517 VSS.n8547 VSS.n8546 0.00317857
R29518 VSS.n8552 VSS.n8214 0.00317857
R29519 VSS.n8477 VSS.n8278 0.00317857
R29520 VSS.n8481 VSS.n8480 0.00317857
R29521 VSS.n8521 VSS.n8244 0.00317857
R29522 VSS.n8548 VSS.n8226 0.00317857
R29523 VSS.n8553 VSS.n8551 0.00317857
R29524 VSS.n8567 VSS.n8566 0.00317857
R29525 VSS.n8644 VSS.n8183 0.00317857
R29526 VSS.n8656 VSS.n8178 0.00317857
R29527 VSS.n8686 VSS.n8165 0.00317857
R29528 VSS.n8710 VSS.n8709 0.00317857
R29529 VSS.n8728 VSS.n8727 0.00317857
R29530 VSS.n8688 VSS.n8687 0.00317857
R29531 VSS.n8379 VSS.n8358 0.00317857
R29532 VSS.n8383 VSS.n8382 0.00317857
R29533 VSS.n8411 VSS.n8410 0.00317857
R29534 VSS.n8441 VSS.n8298 0.00317857
R29535 VSS.n8445 VSS.n8444 0.00317857
R29536 VSS.n8970 VSS.n8969 0.00317857
R29537 VSS.n8976 VSS.n8946 0.00317857
R29538 VSS.n9001 VSS.n8919 0.00317857
R29539 VSS.n8912 VSS.n8899 0.00317857
R29540 VSS.n9032 VSS.n8888 0.00317857
R29541 VSS.n9038 VSS.n8881 0.00317857
R29542 VSS.n9068 VSS.n9067 0.00317857
R29543 VSS.n9074 VSS.n8866 0.00317857
R29544 VSS.n9114 VSS.n8835 0.00317857
R29545 VSS.n9123 VSS.n9122 0.00317857
R29546 VSS.n9139 VSS.n9138 0.00317857
R29547 VSS.n9144 VSS.n8806 0.00317857
R29548 VSS.n9069 VSS.n8870 0.00317857
R29549 VSS.n9073 VSS.n9072 0.00317857
R29550 VSS.n9113 VSS.n8836 0.00317857
R29551 VSS.n9140 VSS.n8818 0.00317857
R29552 VSS.n9145 VSS.n9143 0.00317857
R29553 VSS.n9159 VSS.n9158 0.00317857
R29554 VSS.n9236 VSS.n8775 0.00317857
R29555 VSS.n9248 VSS.n8770 0.00317857
R29556 VSS.n9278 VSS.n8757 0.00317857
R29557 VSS.n9302 VSS.n9301 0.00317857
R29558 VSS.n9320 VSS.n9319 0.00317857
R29559 VSS.n9280 VSS.n9279 0.00317857
R29560 VSS.n8971 VSS.n8950 0.00317857
R29561 VSS.n8975 VSS.n8974 0.00317857
R29562 VSS.n9003 VSS.n9002 0.00317857
R29563 VSS.n9033 VSS.n8890 0.00317857
R29564 VSS.n9037 VSS.n9036 0.00317857
R29565 VSS.n10154 VSS.n10153 0.00317857
R29566 VSS.n10160 VSS.n10130 0.00317857
R29567 VSS.n10185 VSS.n10103 0.00317857
R29568 VSS.n10096 VSS.n10083 0.00317857
R29569 VSS.n10216 VSS.n10072 0.00317857
R29570 VSS.n10222 VSS.n10065 0.00317857
R29571 VSS.n10252 VSS.n10251 0.00317857
R29572 VSS.n10258 VSS.n10050 0.00317857
R29573 VSS.n10298 VSS.n10019 0.00317857
R29574 VSS.n10307 VSS.n10306 0.00317857
R29575 VSS.n10323 VSS.n10322 0.00317857
R29576 VSS.n10328 VSS.n9990 0.00317857
R29577 VSS.n10253 VSS.n10054 0.00317857
R29578 VSS.n10257 VSS.n10256 0.00317857
R29579 VSS.n10297 VSS.n10020 0.00317857
R29580 VSS.n10324 VSS.n10002 0.00317857
R29581 VSS.n10329 VSS.n10327 0.00317857
R29582 VSS.n10343 VSS.n10342 0.00317857
R29583 VSS.n10420 VSS.n9959 0.00317857
R29584 VSS.n10432 VSS.n9954 0.00317857
R29585 VSS.n10462 VSS.n9941 0.00317857
R29586 VSS.n10486 VSS.n10485 0.00317857
R29587 VSS.n10504 VSS.n10503 0.00317857
R29588 VSS.n10464 VSS.n10463 0.00317857
R29589 VSS.n10155 VSS.n10134 0.00317857
R29590 VSS.n10159 VSS.n10158 0.00317857
R29591 VSS.n10187 VSS.n10186 0.00317857
R29592 VSS.n10217 VSS.n10074 0.00317857
R29593 VSS.n10221 VSS.n10220 0.00317857
R29594 VSS.n10746 VSS.n10745 0.00317857
R29595 VSS.n10752 VSS.n10722 0.00317857
R29596 VSS.n10777 VSS.n10695 0.00317857
R29597 VSS.n10688 VSS.n10675 0.00317857
R29598 VSS.n10808 VSS.n10664 0.00317857
R29599 VSS.n10814 VSS.n10657 0.00317857
R29600 VSS.n10844 VSS.n10843 0.00317857
R29601 VSS.n10850 VSS.n10642 0.00317857
R29602 VSS.n10890 VSS.n10611 0.00317857
R29603 VSS.n10899 VSS.n10898 0.00317857
R29604 VSS.n10915 VSS.n10914 0.00317857
R29605 VSS.n10920 VSS.n10582 0.00317857
R29606 VSS.n10845 VSS.n10646 0.00317857
R29607 VSS.n10849 VSS.n10848 0.00317857
R29608 VSS.n10889 VSS.n10612 0.00317857
R29609 VSS.n10916 VSS.n10594 0.00317857
R29610 VSS.n10921 VSS.n10919 0.00317857
R29611 VSS.n10935 VSS.n10934 0.00317857
R29612 VSS.n11012 VSS.n10551 0.00317857
R29613 VSS.n11024 VSS.n10546 0.00317857
R29614 VSS.n11054 VSS.n10533 0.00317857
R29615 VSS.n11078 VSS.n11077 0.00317857
R29616 VSS.n11096 VSS.n11095 0.00317857
R29617 VSS.n11056 VSS.n11055 0.00317857
R29618 VSS.n10747 VSS.n10726 0.00317857
R29619 VSS.n10751 VSS.n10750 0.00317857
R29620 VSS.n10779 VSS.n10778 0.00317857
R29621 VSS.n10809 VSS.n10666 0.00317857
R29622 VSS.n10813 VSS.n10812 0.00317857
R29623 VSS.n11338 VSS.n11337 0.00317857
R29624 VSS.n11344 VSS.n11314 0.00317857
R29625 VSS.n11369 VSS.n11287 0.00317857
R29626 VSS.n11280 VSS.n11267 0.00317857
R29627 VSS.n11400 VSS.n11256 0.00317857
R29628 VSS.n11406 VSS.n11249 0.00317857
R29629 VSS.n11436 VSS.n11435 0.00317857
R29630 VSS.n11442 VSS.n11234 0.00317857
R29631 VSS.n11482 VSS.n11203 0.00317857
R29632 VSS.n11491 VSS.n11490 0.00317857
R29633 VSS.n11507 VSS.n11506 0.00317857
R29634 VSS.n11512 VSS.n11174 0.00317857
R29635 VSS.n11437 VSS.n11238 0.00317857
R29636 VSS.n11441 VSS.n11440 0.00317857
R29637 VSS.n11481 VSS.n11204 0.00317857
R29638 VSS.n11508 VSS.n11186 0.00317857
R29639 VSS.n11513 VSS.n11511 0.00317857
R29640 VSS.n11527 VSS.n11526 0.00317857
R29641 VSS.n11604 VSS.n11143 0.00317857
R29642 VSS.n11616 VSS.n11138 0.00317857
R29643 VSS.n11646 VSS.n11125 0.00317857
R29644 VSS.n11670 VSS.n11669 0.00317857
R29645 VSS.n11688 VSS.n11687 0.00317857
R29646 VSS.n11648 VSS.n11647 0.00317857
R29647 VSS.n11339 VSS.n11318 0.00317857
R29648 VSS.n11343 VSS.n11342 0.00317857
R29649 VSS.n11371 VSS.n11370 0.00317857
R29650 VSS.n11401 VSS.n11258 0.00317857
R29651 VSS.n11405 VSS.n11404 0.00317857
R29652 VSS.n11930 VSS.n11929 0.00317857
R29653 VSS.n11936 VSS.n11906 0.00317857
R29654 VSS.n11961 VSS.n11879 0.00317857
R29655 VSS.n11872 VSS.n11859 0.00317857
R29656 VSS.n11992 VSS.n11848 0.00317857
R29657 VSS.n11998 VSS.n11841 0.00317857
R29658 VSS.n12028 VSS.n12027 0.00317857
R29659 VSS.n12034 VSS.n11826 0.00317857
R29660 VSS.n12074 VSS.n11795 0.00317857
R29661 VSS.n12083 VSS.n12082 0.00317857
R29662 VSS.n12099 VSS.n12098 0.00317857
R29663 VSS.n12104 VSS.n11766 0.00317857
R29664 VSS.n12029 VSS.n11830 0.00317857
R29665 VSS.n12033 VSS.n12032 0.00317857
R29666 VSS.n12073 VSS.n11796 0.00317857
R29667 VSS.n12100 VSS.n11778 0.00317857
R29668 VSS.n12105 VSS.n12103 0.00317857
R29669 VSS.n12119 VSS.n12118 0.00317857
R29670 VSS.n12196 VSS.n11735 0.00317857
R29671 VSS.n12208 VSS.n11730 0.00317857
R29672 VSS.n12238 VSS.n11717 0.00317857
R29673 VSS.n12262 VSS.n12261 0.00317857
R29674 VSS.n12280 VSS.n12279 0.00317857
R29675 VSS.n12240 VSS.n12239 0.00317857
R29676 VSS.n11931 VSS.n11910 0.00317857
R29677 VSS.n11935 VSS.n11934 0.00317857
R29678 VSS.n11963 VSS.n11962 0.00317857
R29679 VSS.n11993 VSS.n11850 0.00317857
R29680 VSS.n11997 VSS.n11996 0.00317857
R29681 VSS.n12522 VSS.n12521 0.00317857
R29682 VSS.n12528 VSS.n12498 0.00317857
R29683 VSS.n12553 VSS.n12471 0.00317857
R29684 VSS.n12464 VSS.n12451 0.00317857
R29685 VSS.n12584 VSS.n12440 0.00317857
R29686 VSS.n12590 VSS.n12433 0.00317857
R29687 VSS.n12620 VSS.n12619 0.00317857
R29688 VSS.n12626 VSS.n12418 0.00317857
R29689 VSS.n12666 VSS.n12387 0.00317857
R29690 VSS.n12675 VSS.n12674 0.00317857
R29691 VSS.n12691 VSS.n12690 0.00317857
R29692 VSS.n12696 VSS.n12358 0.00317857
R29693 VSS.n12621 VSS.n12422 0.00317857
R29694 VSS.n12625 VSS.n12624 0.00317857
R29695 VSS.n12665 VSS.n12388 0.00317857
R29696 VSS.n12692 VSS.n12370 0.00317857
R29697 VSS.n12697 VSS.n12695 0.00317857
R29698 VSS.n12711 VSS.n12710 0.00317857
R29699 VSS.n12788 VSS.n12327 0.00317857
R29700 VSS.n12800 VSS.n12322 0.00317857
R29701 VSS.n12830 VSS.n12309 0.00317857
R29702 VSS.n12854 VSS.n12853 0.00317857
R29703 VSS.n12872 VSS.n12871 0.00317857
R29704 VSS.n12832 VSS.n12831 0.00317857
R29705 VSS.n12523 VSS.n12502 0.00317857
R29706 VSS.n12527 VSS.n12526 0.00317857
R29707 VSS.n12555 VSS.n12554 0.00317857
R29708 VSS.n12585 VSS.n12442 0.00317857
R29709 VSS.n12589 VSS.n12588 0.00317857
R29710 VSS.n13114 VSS.n13113 0.00317857
R29711 VSS.n13120 VSS.n13090 0.00317857
R29712 VSS.n13145 VSS.n13063 0.00317857
R29713 VSS.n13056 VSS.n13043 0.00317857
R29714 VSS.n13176 VSS.n13032 0.00317857
R29715 VSS.n13182 VSS.n13025 0.00317857
R29716 VSS.n13212 VSS.n13211 0.00317857
R29717 VSS.n13218 VSS.n13010 0.00317857
R29718 VSS.n13258 VSS.n12979 0.00317857
R29719 VSS.n13267 VSS.n13266 0.00317857
R29720 VSS.n13283 VSS.n13282 0.00317857
R29721 VSS.n13288 VSS.n12950 0.00317857
R29722 VSS.n13213 VSS.n13014 0.00317857
R29723 VSS.n13217 VSS.n13216 0.00317857
R29724 VSS.n13257 VSS.n12980 0.00317857
R29725 VSS.n13284 VSS.n12962 0.00317857
R29726 VSS.n13289 VSS.n13287 0.00317857
R29727 VSS.n13303 VSS.n13302 0.00317857
R29728 VSS.n13380 VSS.n12919 0.00317857
R29729 VSS.n13392 VSS.n12914 0.00317857
R29730 VSS.n13422 VSS.n12901 0.00317857
R29731 VSS.n13446 VSS.n13445 0.00317857
R29732 VSS.n13464 VSS.n13463 0.00317857
R29733 VSS.n13424 VSS.n13423 0.00317857
R29734 VSS.n13115 VSS.n13094 0.00317857
R29735 VSS.n13119 VSS.n13118 0.00317857
R29736 VSS.n13147 VSS.n13146 0.00317857
R29737 VSS.n13177 VSS.n13034 0.00317857
R29738 VSS.n13181 VSS.n13180 0.00317857
R29739 VSS.n13706 VSS.n13705 0.00317857
R29740 VSS.n13712 VSS.n13682 0.00317857
R29741 VSS.n13737 VSS.n13655 0.00317857
R29742 VSS.n13648 VSS.n13635 0.00317857
R29743 VSS.n13768 VSS.n13624 0.00317857
R29744 VSS.n13774 VSS.n13617 0.00317857
R29745 VSS.n13804 VSS.n13803 0.00317857
R29746 VSS.n13810 VSS.n13602 0.00317857
R29747 VSS.n13850 VSS.n13571 0.00317857
R29748 VSS.n13859 VSS.n13858 0.00317857
R29749 VSS.n13875 VSS.n13874 0.00317857
R29750 VSS.n13880 VSS.n13542 0.00317857
R29751 VSS.n13805 VSS.n13606 0.00317857
R29752 VSS.n13809 VSS.n13808 0.00317857
R29753 VSS.n13849 VSS.n13572 0.00317857
R29754 VSS.n13876 VSS.n13554 0.00317857
R29755 VSS.n13881 VSS.n13879 0.00317857
R29756 VSS.n13895 VSS.n13894 0.00317857
R29757 VSS.n13972 VSS.n13511 0.00317857
R29758 VSS.n13984 VSS.n13506 0.00317857
R29759 VSS.n14014 VSS.n13493 0.00317857
R29760 VSS.n14038 VSS.n14037 0.00317857
R29761 VSS.n14056 VSS.n14055 0.00317857
R29762 VSS.n14016 VSS.n14015 0.00317857
R29763 VSS.n13707 VSS.n13686 0.00317857
R29764 VSS.n13711 VSS.n13710 0.00317857
R29765 VSS.n13739 VSS.n13738 0.00317857
R29766 VSS.n13769 VSS.n13626 0.00317857
R29767 VSS.n13773 VSS.n13772 0.00317857
R29768 VSS.n14298 VSS.n14297 0.00317857
R29769 VSS.n14304 VSS.n14274 0.00317857
R29770 VSS.n14329 VSS.n14247 0.00317857
R29771 VSS.n14240 VSS.n14227 0.00317857
R29772 VSS.n14360 VSS.n14216 0.00317857
R29773 VSS.n14366 VSS.n14209 0.00317857
R29774 VSS.n14396 VSS.n14395 0.00317857
R29775 VSS.n14402 VSS.n14194 0.00317857
R29776 VSS.n14442 VSS.n14163 0.00317857
R29777 VSS.n14451 VSS.n14450 0.00317857
R29778 VSS.n14467 VSS.n14466 0.00317857
R29779 VSS.n14472 VSS.n14134 0.00317857
R29780 VSS.n14397 VSS.n14198 0.00317857
R29781 VSS.n14401 VSS.n14400 0.00317857
R29782 VSS.n14441 VSS.n14164 0.00317857
R29783 VSS.n14468 VSS.n14146 0.00317857
R29784 VSS.n14473 VSS.n14471 0.00317857
R29785 VSS.n14487 VSS.n14486 0.00317857
R29786 VSS.n14564 VSS.n14103 0.00317857
R29787 VSS.n14576 VSS.n14098 0.00317857
R29788 VSS.n14606 VSS.n14085 0.00317857
R29789 VSS.n14630 VSS.n14629 0.00317857
R29790 VSS.n14648 VSS.n14647 0.00317857
R29791 VSS.n14608 VSS.n14607 0.00317857
R29792 VSS.n14299 VSS.n14278 0.00317857
R29793 VSS.n14303 VSS.n14302 0.00317857
R29794 VSS.n14331 VSS.n14330 0.00317857
R29795 VSS.n14361 VSS.n14218 0.00317857
R29796 VSS.n14365 VSS.n14364 0.00317857
R29797 VSS.n14890 VSS.n14889 0.00317857
R29798 VSS.n14896 VSS.n14866 0.00317857
R29799 VSS.n14921 VSS.n14839 0.00317857
R29800 VSS.n14832 VSS.n14819 0.00317857
R29801 VSS.n14952 VSS.n14808 0.00317857
R29802 VSS.n14958 VSS.n14801 0.00317857
R29803 VSS.n14988 VSS.n14987 0.00317857
R29804 VSS.n14994 VSS.n14786 0.00317857
R29805 VSS.n15034 VSS.n14755 0.00317857
R29806 VSS.n15043 VSS.n15042 0.00317857
R29807 VSS.n15059 VSS.n15058 0.00317857
R29808 VSS.n15064 VSS.n14726 0.00317857
R29809 VSS.n14989 VSS.n14790 0.00317857
R29810 VSS.n14993 VSS.n14992 0.00317857
R29811 VSS.n15033 VSS.n14756 0.00317857
R29812 VSS.n15060 VSS.n14738 0.00317857
R29813 VSS.n15065 VSS.n15063 0.00317857
R29814 VSS.n15079 VSS.n15078 0.00317857
R29815 VSS.n15156 VSS.n14695 0.00317857
R29816 VSS.n15168 VSS.n14690 0.00317857
R29817 VSS.n15198 VSS.n14677 0.00317857
R29818 VSS.n15222 VSS.n15221 0.00317857
R29819 VSS.n15240 VSS.n15239 0.00317857
R29820 VSS.n15200 VSS.n15199 0.00317857
R29821 VSS.n14891 VSS.n14870 0.00317857
R29822 VSS.n14895 VSS.n14894 0.00317857
R29823 VSS.n14923 VSS.n14922 0.00317857
R29824 VSS.n14953 VSS.n14810 0.00317857
R29825 VSS.n14957 VSS.n14956 0.00317857
R29826 VSS.n15482 VSS.n15481 0.00317857
R29827 VSS.n15488 VSS.n15458 0.00317857
R29828 VSS.n15513 VSS.n15431 0.00317857
R29829 VSS.n15424 VSS.n15411 0.00317857
R29830 VSS.n15544 VSS.n15400 0.00317857
R29831 VSS.n15550 VSS.n15393 0.00317857
R29832 VSS.n15580 VSS.n15579 0.00317857
R29833 VSS.n15586 VSS.n15378 0.00317857
R29834 VSS.n15626 VSS.n15347 0.00317857
R29835 VSS.n15635 VSS.n15634 0.00317857
R29836 VSS.n15651 VSS.n15650 0.00317857
R29837 VSS.n15656 VSS.n15318 0.00317857
R29838 VSS.n15581 VSS.n15382 0.00317857
R29839 VSS.n15585 VSS.n15584 0.00317857
R29840 VSS.n15625 VSS.n15348 0.00317857
R29841 VSS.n15652 VSS.n15330 0.00317857
R29842 VSS.n15657 VSS.n15655 0.00317857
R29843 VSS.n15671 VSS.n15670 0.00317857
R29844 VSS.n15748 VSS.n15287 0.00317857
R29845 VSS.n15760 VSS.n15282 0.00317857
R29846 VSS.n15790 VSS.n15269 0.00317857
R29847 VSS.n15814 VSS.n15813 0.00317857
R29848 VSS.n15832 VSS.n15831 0.00317857
R29849 VSS.n15792 VSS.n15791 0.00317857
R29850 VSS.n15483 VSS.n15462 0.00317857
R29851 VSS.n15487 VSS.n15486 0.00317857
R29852 VSS.n15515 VSS.n15514 0.00317857
R29853 VSS.n15545 VSS.n15402 0.00317857
R29854 VSS.n15549 VSS.n15548 0.00317857
R29855 VSS.n6590 VSS.n6589 0.00317857
R29856 VSS.n6596 VSS.n6566 0.00317857
R29857 VSS.n6621 VSS.n6539 0.00317857
R29858 VSS.n6532 VSS.n6519 0.00317857
R29859 VSS.n6652 VSS.n6508 0.00317857
R29860 VSS.n6658 VSS.n6501 0.00317857
R29861 VSS.n6744 VSS.n6498 0.00317857
R29862 VSS.n15957 VSS.n6683 0.00317857
R29863 VSS.n15942 VSS.n15941 0.00317857
R29864 VSS.n6780 VSS.n6706 0.00317857
R29865 VSS.n15932 VSS.n6707 0.00317857
R29866 VSS.n15927 VSS.n6712 0.00317857
R29867 VSS.n6743 VSS.n6679 0.00317857
R29868 VSS.n15958 VSS.n6681 0.00317857
R29869 VSS.n15943 VSS.n6696 0.00317857
R29870 VSS.n15931 VSS.n6708 0.00317857
R29871 VSS.n15928 VSS.n6710 0.00317857
R29872 VSS.n6825 VSS.n6824 0.00317857
R29873 VSS.n6882 VSS.n6869 0.00317857
R29874 VSS.n6916 VSS.n6864 0.00317857
R29875 VSS.n15860 VSS.n15859 0.00317857
R29876 VSS.n6950 VSS.n6949 0.00317857
R29877 VSS.n15841 VSS.n6937 0.00317857
R29878 VSS.n15858 VSS.n6897 0.00317857
R29879 VSS.n6591 VSS.n6570 0.00317857
R29880 VSS.n6595 VSS.n6594 0.00317857
R29881 VSS.n6623 VSS.n6622 0.00317857
R29882 VSS.n6653 VSS.n6510 0.00317857
R29883 VSS.n6657 VSS.n6656 0.00317857
R29884 VSS.n7187 VSS.n7186 0.00317857
R29885 VSS.n7193 VSS.n7164 0.00317857
R29886 VSS.n7226 VSS.n7139 0.00317857
R29887 VSS.n7242 VSS.n7241 0.00317857
R29888 VSS.n7259 VSS.n7258 0.00317857
R29889 VSS.n7264 VSS.n7104 0.00317857
R29890 VSS.n7292 VSS.n7291 0.00317857
R29891 VSS.n7298 VSS.n7089 0.00317857
R29892 VSS.n7338 VSS.n7058 0.00317857
R29893 VSS.n7347 VSS.n7346 0.00317857
R29894 VSS.n7363 VSS.n7362 0.00317857
R29895 VSS.n7368 VSS.n7029 0.00317857
R29896 VSS.n7293 VSS.n7093 0.00317857
R29897 VSS.n7297 VSS.n7296 0.00317857
R29898 VSS.n7337 VSS.n7059 0.00317857
R29899 VSS.n7364 VSS.n7041 0.00317857
R29900 VSS.n7369 VSS.n7367 0.00317857
R29901 VSS.n7383 VSS.n7382 0.00317857
R29902 VSS.n7460 VSS.n6998 0.00317857
R29903 VSS.n7472 VSS.n6993 0.00317857
R29904 VSS.n7502 VSS.n6980 0.00317857
R29905 VSS.n7526 VSS.n7525 0.00317857
R29906 VSS.n7544 VSS.n7543 0.00317857
R29907 VSS.n7504 VSS.n7503 0.00317857
R29908 VSS.n7188 VSS.n7168 0.00317857
R29909 VSS.n7192 VSS.n7191 0.00317857
R29910 VSS.n7227 VSS.n7137 0.00317857
R29911 VSS.n7260 VSS.n7116 0.00317857
R29912 VSS.n7265 VSS.n7263 0.00317857
R29913 VSS.n348 VSS.n291 0.00317857
R29914 VSS.n443 VSS.n297 0.00317857
R29915 VSS.n434 VSS.n304 0.00317857
R29916 VSS.n392 VSS.n321 0.00317857
R29917 VSS.n418 VSS.n322 0.00317857
R29918 VSS.n412 VSS.n195 0.00317857
R29919 VSS.n18604 VSS.n18603 0.00317857
R29920 VSS.n18610 VSS.n187 0.00317857
R29921 VSS.n18650 VSS.n156 0.00317857
R29922 VSS.n18659 VSS.n18658 0.00317857
R29923 VSS.n18675 VSS.n18674 0.00317857
R29924 VSS.n18680 VSS.n127 0.00317857
R29925 VSS.n18605 VSS.n191 0.00317857
R29926 VSS.n18609 VSS.n18608 0.00317857
R29927 VSS.n18649 VSS.n157 0.00317857
R29928 VSS.n18676 VSS.n139 0.00317857
R29929 VSS.n18681 VSS.n18679 0.00317857
R29930 VSS.n18695 VSS.n18694 0.00317857
R29931 VSS.n18772 VSS.n96 0.00317857
R29932 VSS.n18784 VSS.n91 0.00317857
R29933 VSS.n18814 VSS.n78 0.00317857
R29934 VSS.n18838 VSS.n18837 0.00317857
R29935 VSS.n18856 VSS.n18855 0.00317857
R29936 VSS.n18816 VSS.n18815 0.00317857
R29937 VSS.n347 VSS.n293 0.00317857
R29938 VSS.n444 VSS.n295 0.00317857
R29939 VSS.n433 VSS.n432 0.00317857
R29940 VSS.n417 VSS.n323 0.00317857
R29941 VSS.n414 VSS.n413 0.00317857
R29942 VSS.n876 VSS.n498 0.00317857
R29943 VSS.n871 VSS.n503 0.00317857
R29944 VSS.n856 VSS.n855 0.00317857
R29945 VSS.n603 VSS.n526 0.00317857
R29946 VSS.n846 VSS.n527 0.00317857
R29947 VSS.n841 VSS.n532 0.00317857
R29948 VSS.n875 VSS.n499 0.00317857
R29949 VSS.n872 VSS.n501 0.00317857
R29950 VSS.n857 VSS.n516 0.00317857
R29951 VSS.n845 VSS.n528 0.00317857
R29952 VSS.n842 VSS.n530 0.00317857
R29953 VSS.n648 VSS.n647 0.00317857
R29954 VSS.n705 VSS.n692 0.00317857
R29955 VSS.n748 VSS.n687 0.00317857
R29956 VSS.n774 VSS.n773 0.00317857
R29957 VSS.n737 VSS.n736 0.00317857
R29958 VSS.n18864 VSS.n50 0.00317857
R29959 VSS.n772 VSS.n720 0.00317857
R29960 VSS.n911 VSS.n459 0.00317857
R29961 VSS.n1009 VSS.n461 0.00317857
R29962 VSS.n998 VSS.n997 0.00317857
R29963 VSS.n982 VSS.n489 0.00317857
R29964 VSS.n979 VSS.n491 0.00317857
R29965 VSS.n1307 VSS.n1306 0.00317857
R29966 VSS.n1364 VSS.n1351 0.00317857
R29967 VSS.n1398 VSS.n1346 0.00317857
R29968 VSS.n17888 VSS.n17887 0.00317857
R29969 VSS.n1432 VSS.n1431 0.00317857
R29970 VSS.n17869 VSS.n1419 0.00317857
R29971 VSS.n17886 VSS.n1379 0.00317857
R29972 VSS.n9589 VSS.n9516 0.00316667
R29973 VSS.n9599 VSS.n9493 0.00316667
R29974 VSS.n1235 VSS.n1166 0.00228571
R29975 VSS.n1240 VSS.n1235 0.00228571
R29976 VSS.n1236 VSS.n1215 0.00228571
R29977 VSS.n17976 VSS.n1172 0.00228571
R29978 VSS.n1267 VSS.n1266 0.00228571
R29979 VSS.n17975 VSS.n17974 0.00228571
R29980 VSS.n922 VSS.n901 0.00228571
R29981 VSS.n993 VSS.n992 0.00228571
R29982 VSS.n951 VSS.n950 0.00228571
R29983 VSS.n17035 VSS.n16985 0.00228571
R29984 VSS.n17035 VSS.n17034 0.00228571
R29985 VSS.n17046 VSS.n16977 0.00228571
R29986 VSS.n17057 VSS.n16969 0.00228571
R29987 VSS.n17078 VSS.n17077 0.00228571
R29988 VSS.n1103 VSS.n1082 0.00228571
R29989 VSS.n18019 VSS.n18018 0.00228571
R29990 VSS.n1132 VSS.n1131 0.00228571
R29991 VSS.n18020 VSS.n1044 0.00228571
R29992 VSS.n16924 VSS.n16921 0.00228571
R29993 VSS.n17160 VSS.n17159 0.00228571
R29994 VSS.n16911 VSS.n16905 0.00228571
R29995 VSS.n17233 VSS.n16884 0.00228571
R29996 VSS.n17243 VSS.n17242 0.00228571
R29997 VSS.n17058 VSS.n16967 0.00228571
R29998 VSS.n17627 VSS.n17399 0.00228571
R29999 VSS.n17627 VSS.n17626 0.00228571
R30000 VSS.n17638 VSS.n17391 0.00228571
R30001 VSS.n17649 VSS.n17383 0.00228571
R30002 VSS.n17670 VSS.n17669 0.00228571
R30003 VSS.n17533 VSS.n17476 0.00228571
R30004 VSS.n17464 VSS.n17463 0.00228571
R30005 VSS.n17565 VSS.n17447 0.00228571
R30006 VSS.n17551 VSS.n17465 0.00228571
R30007 VSS.n17338 VSS.n17335 0.00228571
R30008 VSS.n17752 VSS.n17751 0.00228571
R30009 VSS.n17325 VSS.n17319 0.00228571
R30010 VSS.n17825 VSS.n17298 0.00228571
R30011 VSS.n17835 VSS.n17834 0.00228571
R30012 VSS.n17650 VSS.n17381 0.00228571
R30013 VSS.n18110 VSS.n268 0.00228571
R30014 VSS.n256 VSS.n255 0.00228571
R30015 VSS.n18142 VSS.n239 0.00228571
R30016 VSS.n18252 VSS.n18183 0.00228571
R30017 VSS.n18257 VSS.n18252 0.00228571
R30018 VSS.n18253 VSS.n18232 0.00228571
R30019 VSS.n18565 VSS.n18189 0.00228571
R30020 VSS.n18284 VSS.n18283 0.00228571
R30021 VSS.n18564 VSS.n18563 0.00228571
R30022 VSS.n18363 VSS.n18316 0.00228571
R30023 VSS.n18513 VSS.n18340 0.00228571
R30024 VSS.n18507 VSS.n18506 0.00228571
R30025 VSS.n18447 VSS.n18443 0.00228571
R30026 VSS.n18422 VSS.n18419 0.00228571
R30027 VSS.n18128 VSS.n257 0.00228571
R30028 VSS.n9583 VSS.n9526 0.00228571
R30029 VSS.n9514 VSS.n9513 0.00228571
R30030 VSS.n9615 VSS.n9497 0.00228571
R30031 VSS.n9677 VSS.n9449 0.00228571
R30032 VSS.n9677 VSS.n9676 0.00228571
R30033 VSS.n9688 VSS.n9441 0.00228571
R30034 VSS.n9699 VSS.n9433 0.00228571
R30035 VSS.n9720 VSS.n9719 0.00228571
R30036 VSS.n9700 VSS.n9431 0.00228571
R30037 VSS.n9388 VSS.n9385 0.00228571
R30038 VSS.n9802 VSS.n9801 0.00228571
R30039 VSS.n9375 VSS.n9369 0.00228571
R30040 VSS.n9875 VSS.n9348 0.00228571
R30041 VSS.n9885 VSS.n9884 0.00228571
R30042 VSS.n9601 VSS.n9515 0.00228571
R30043 VSS.n16526 VSS.n16460 0.00228571
R30044 VSS.n16544 VSS.n16444 0.00228571
R30045 VSS.n16558 VSS.n16557 0.00228571
R30046 VSS.n16620 VSS.n16391 0.00228571
R30047 VSS.n16620 VSS.n16619 0.00228571
R30048 VSS.n16631 VSS.n16383 0.00228571
R30049 VSS.n16642 VSS.n16375 0.00228571
R30050 VSS.n16663 VSS.n16662 0.00228571
R30051 VSS.n16643 VSS.n16373 0.00228571
R30052 VSS.n16330 VSS.n16327 0.00228571
R30053 VSS.n16745 VSS.n16744 0.00228571
R30054 VSS.n16317 VSS.n16311 0.00228571
R30055 VSS.n16818 VSS.n16290 0.00228571
R30056 VSS.n16828 VSS.n16827 0.00228571
R30057 VSS.n16543 VSS.n16445 0.00228571
R30058 VSS.n1691 VSS.n1625 0.00228571
R30059 VSS.n1709 VSS.n1609 0.00228571
R30060 VSS.n1723 VSS.n1722 0.00228571
R30061 VSS.n16027 VSS.n1563 0.00228571
R30062 VSS.n16027 VSS.n16026 0.00228571
R30063 VSS.n16038 VSS.n1555 0.00228571
R30064 VSS.n16049 VSS.n1547 0.00228571
R30065 VSS.n16070 VSS.n16069 0.00228571
R30066 VSS.n16050 VSS.n1545 0.00228571
R30067 VSS.n1502 VSS.n1499 0.00228571
R30068 VSS.n16152 VSS.n16151 0.00228571
R30069 VSS.n1489 VSS.n1483 0.00228571
R30070 VSS.n16225 VSS.n1462 0.00228571
R30071 VSS.n16235 VSS.n16234 0.00228571
R30072 VSS.n1708 VSS.n1610 0.00228571
R30073 VSS.n1875 VSS.n1818 0.00228571
R30074 VSS.n1806 VSS.n1805 0.00228571
R30075 VSS.n1907 VSS.n1789 0.00228571
R30076 VSS.n2017 VSS.n1948 0.00228571
R30077 VSS.n2022 VSS.n2017 0.00228571
R30078 VSS.n2018 VSS.n1997 0.00228571
R30079 VSS.n2330 VSS.n1954 0.00228571
R30080 VSS.n2049 VSS.n2048 0.00228571
R30081 VSS.n2329 VSS.n2328 0.00228571
R30082 VSS.n2287 VSS.n2286 0.00228571
R30083 VSS.n2276 VSS.n2275 0.00228571
R30084 VSS.n2134 VSS.n2120 0.00228571
R30085 VSS.n2162 VSS.n2159 0.00228571
R30086 VSS.n2235 VSS.n2171 0.00228571
R30087 VSS.n1893 VSS.n1807 0.00228571
R30088 VSS.n3074 VSS.n3017 0.00228571
R30089 VSS.n3005 VSS.n3004 0.00228571
R30090 VSS.n3106 VSS.n2988 0.00228571
R30091 VSS.n3168 VSS.n2940 0.00228571
R30092 VSS.n3168 VSS.n3167 0.00228571
R30093 VSS.n3179 VSS.n2932 0.00228571
R30094 VSS.n3190 VSS.n2924 0.00228571
R30095 VSS.n3211 VSS.n3210 0.00228571
R30096 VSS.n3191 VSS.n2922 0.00228571
R30097 VSS.n2879 VSS.n2876 0.00228571
R30098 VSS.n3293 VSS.n3292 0.00228571
R30099 VSS.n2866 VSS.n2860 0.00228571
R30100 VSS.n3366 VSS.n2839 0.00228571
R30101 VSS.n3376 VSS.n3375 0.00228571
R30102 VSS.n3092 VSS.n3006 0.00228571
R30103 VSS.n3666 VSS.n3609 0.00228571
R30104 VSS.n3597 VSS.n3596 0.00228571
R30105 VSS.n3698 VSS.n3580 0.00228571
R30106 VSS.n3760 VSS.n3532 0.00228571
R30107 VSS.n3760 VSS.n3759 0.00228571
R30108 VSS.n3771 VSS.n3524 0.00228571
R30109 VSS.n3782 VSS.n3516 0.00228571
R30110 VSS.n3803 VSS.n3802 0.00228571
R30111 VSS.n3783 VSS.n3514 0.00228571
R30112 VSS.n3471 VSS.n3468 0.00228571
R30113 VSS.n3885 VSS.n3884 0.00228571
R30114 VSS.n3458 VSS.n3452 0.00228571
R30115 VSS.n3958 VSS.n3431 0.00228571
R30116 VSS.n3968 VSS.n3967 0.00228571
R30117 VSS.n3684 VSS.n3598 0.00228571
R30118 VSS.n4258 VSS.n4201 0.00228571
R30119 VSS.n4189 VSS.n4188 0.00228571
R30120 VSS.n4290 VSS.n4172 0.00228571
R30121 VSS.n4352 VSS.n4124 0.00228571
R30122 VSS.n4352 VSS.n4351 0.00228571
R30123 VSS.n4363 VSS.n4116 0.00228571
R30124 VSS.n4374 VSS.n4108 0.00228571
R30125 VSS.n4395 VSS.n4394 0.00228571
R30126 VSS.n4375 VSS.n4106 0.00228571
R30127 VSS.n4063 VSS.n4060 0.00228571
R30128 VSS.n4477 VSS.n4476 0.00228571
R30129 VSS.n4050 VSS.n4044 0.00228571
R30130 VSS.n4550 VSS.n4023 0.00228571
R30131 VSS.n4560 VSS.n4559 0.00228571
R30132 VSS.n4276 VSS.n4190 0.00228571
R30133 VSS.n4850 VSS.n4793 0.00228571
R30134 VSS.n4781 VSS.n4780 0.00228571
R30135 VSS.n4882 VSS.n4764 0.00228571
R30136 VSS.n4944 VSS.n4716 0.00228571
R30137 VSS.n4944 VSS.n4943 0.00228571
R30138 VSS.n4955 VSS.n4708 0.00228571
R30139 VSS.n4966 VSS.n4700 0.00228571
R30140 VSS.n4987 VSS.n4986 0.00228571
R30141 VSS.n4967 VSS.n4698 0.00228571
R30142 VSS.n4655 VSS.n4652 0.00228571
R30143 VSS.n5069 VSS.n5068 0.00228571
R30144 VSS.n4642 VSS.n4636 0.00228571
R30145 VSS.n5142 VSS.n4615 0.00228571
R30146 VSS.n5152 VSS.n5151 0.00228571
R30147 VSS.n4868 VSS.n4782 0.00228571
R30148 VSS.n2471 VSS.n2414 0.00228571
R30149 VSS.n2402 VSS.n2401 0.00228571
R30150 VSS.n2503 VSS.n2385 0.00228571
R30151 VSS.n2613 VSS.n2544 0.00228571
R30152 VSS.n2618 VSS.n2613 0.00228571
R30153 VSS.n2614 VSS.n2593 0.00228571
R30154 VSS.n5295 VSS.n2550 0.00228571
R30155 VSS.n2645 VSS.n2644 0.00228571
R30156 VSS.n5294 VSS.n5293 0.00228571
R30157 VSS.n5252 VSS.n5251 0.00228571
R30158 VSS.n5241 VSS.n5240 0.00228571
R30159 VSS.n2730 VSS.n2716 0.00228571
R30160 VSS.n2758 VSS.n2755 0.00228571
R30161 VSS.n5200 VSS.n2767 0.00228571
R30162 VSS.n2489 VSS.n2403 0.00228571
R30163 VSS.n5432 VSS.n5375 0.00228571
R30164 VSS.n5363 VSS.n5362 0.00228571
R30165 VSS.n5464 VSS.n5346 0.00228571
R30166 VSS.n5574 VSS.n5505 0.00228571
R30167 VSS.n5579 VSS.n5574 0.00228571
R30168 VSS.n5575 VSS.n5554 0.00228571
R30169 VSS.n5868 VSS.n5511 0.00228571
R30170 VSS.n5606 VSS.n5605 0.00228571
R30171 VSS.n5867 VSS.n5866 0.00228571
R30172 VSS.n5825 VSS.n5824 0.00228571
R30173 VSS.n5814 VSS.n5813 0.00228571
R30174 VSS.n5691 VSS.n5677 0.00228571
R30175 VSS.n5719 VSS.n5716 0.00228571
R30176 VSS.n5773 VSS.n5728 0.00228571
R30177 VSS.n5450 VSS.n5364 0.00228571
R30178 VSS.n6005 VSS.n5948 0.00228571
R30179 VSS.n5936 VSS.n5935 0.00228571
R30180 VSS.n6037 VSS.n5919 0.00228571
R30181 VSS.n6147 VSS.n6078 0.00228571
R30182 VSS.n6152 VSS.n6147 0.00228571
R30183 VSS.n6148 VSS.n6127 0.00228571
R30184 VSS.n6460 VSS.n6084 0.00228571
R30185 VSS.n6179 VSS.n6178 0.00228571
R30186 VSS.n6459 VSS.n6458 0.00228571
R30187 VSS.n6417 VSS.n6416 0.00228571
R30188 VSS.n6406 VSS.n6405 0.00228571
R30189 VSS.n6264 VSS.n6250 0.00228571
R30190 VSS.n6292 VSS.n6289 0.00228571
R30191 VSS.n6365 VSS.n6301 0.00228571
R30192 VSS.n6023 VSS.n5937 0.00228571
R30193 VSS.n7807 VSS.n7750 0.00228571
R30194 VSS.n7738 VSS.n7737 0.00228571
R30195 VSS.n7839 VSS.n7721 0.00228571
R30196 VSS.n7901 VSS.n7673 0.00228571
R30197 VSS.n7901 VSS.n7900 0.00228571
R30198 VSS.n7912 VSS.n7665 0.00228571
R30199 VSS.n7923 VSS.n7657 0.00228571
R30200 VSS.n7944 VSS.n7943 0.00228571
R30201 VSS.n7924 VSS.n7655 0.00228571
R30202 VSS.n7612 VSS.n7609 0.00228571
R30203 VSS.n8026 VSS.n8025 0.00228571
R30204 VSS.n7599 VSS.n7593 0.00228571
R30205 VSS.n8099 VSS.n7572 0.00228571
R30206 VSS.n8109 VSS.n8108 0.00228571
R30207 VSS.n7825 VSS.n7739 0.00228571
R30208 VSS.n8399 VSS.n8342 0.00228571
R30209 VSS.n8330 VSS.n8329 0.00228571
R30210 VSS.n8431 VSS.n8313 0.00228571
R30211 VSS.n8493 VSS.n8265 0.00228571
R30212 VSS.n8493 VSS.n8492 0.00228571
R30213 VSS.n8504 VSS.n8257 0.00228571
R30214 VSS.n8515 VSS.n8249 0.00228571
R30215 VSS.n8536 VSS.n8535 0.00228571
R30216 VSS.n8516 VSS.n8247 0.00228571
R30217 VSS.n8204 VSS.n8201 0.00228571
R30218 VSS.n8618 VSS.n8617 0.00228571
R30219 VSS.n8191 VSS.n8185 0.00228571
R30220 VSS.n8691 VSS.n8164 0.00228571
R30221 VSS.n8701 VSS.n8700 0.00228571
R30222 VSS.n8417 VSS.n8331 0.00228571
R30223 VSS.n8991 VSS.n8934 0.00228571
R30224 VSS.n8922 VSS.n8921 0.00228571
R30225 VSS.n9023 VSS.n8905 0.00228571
R30226 VSS.n9085 VSS.n8857 0.00228571
R30227 VSS.n9085 VSS.n9084 0.00228571
R30228 VSS.n9096 VSS.n8849 0.00228571
R30229 VSS.n9107 VSS.n8841 0.00228571
R30230 VSS.n9128 VSS.n9127 0.00228571
R30231 VSS.n9108 VSS.n8839 0.00228571
R30232 VSS.n8796 VSS.n8793 0.00228571
R30233 VSS.n9210 VSS.n9209 0.00228571
R30234 VSS.n8783 VSS.n8777 0.00228571
R30235 VSS.n9283 VSS.n8756 0.00228571
R30236 VSS.n9293 VSS.n9292 0.00228571
R30237 VSS.n9009 VSS.n8923 0.00228571
R30238 VSS.n10175 VSS.n10118 0.00228571
R30239 VSS.n10106 VSS.n10105 0.00228571
R30240 VSS.n10207 VSS.n10089 0.00228571
R30241 VSS.n10269 VSS.n10041 0.00228571
R30242 VSS.n10269 VSS.n10268 0.00228571
R30243 VSS.n10280 VSS.n10033 0.00228571
R30244 VSS.n10291 VSS.n10025 0.00228571
R30245 VSS.n10312 VSS.n10311 0.00228571
R30246 VSS.n10292 VSS.n10023 0.00228571
R30247 VSS.n9980 VSS.n9977 0.00228571
R30248 VSS.n10394 VSS.n10393 0.00228571
R30249 VSS.n9967 VSS.n9961 0.00228571
R30250 VSS.n10467 VSS.n9940 0.00228571
R30251 VSS.n10477 VSS.n10476 0.00228571
R30252 VSS.n10193 VSS.n10107 0.00228571
R30253 VSS.n10767 VSS.n10710 0.00228571
R30254 VSS.n10698 VSS.n10697 0.00228571
R30255 VSS.n10799 VSS.n10681 0.00228571
R30256 VSS.n10861 VSS.n10633 0.00228571
R30257 VSS.n10861 VSS.n10860 0.00228571
R30258 VSS.n10872 VSS.n10625 0.00228571
R30259 VSS.n10883 VSS.n10617 0.00228571
R30260 VSS.n10904 VSS.n10903 0.00228571
R30261 VSS.n10884 VSS.n10615 0.00228571
R30262 VSS.n10572 VSS.n10569 0.00228571
R30263 VSS.n10986 VSS.n10985 0.00228571
R30264 VSS.n10559 VSS.n10553 0.00228571
R30265 VSS.n11059 VSS.n10532 0.00228571
R30266 VSS.n11069 VSS.n11068 0.00228571
R30267 VSS.n10785 VSS.n10699 0.00228571
R30268 VSS.n11359 VSS.n11302 0.00228571
R30269 VSS.n11290 VSS.n11289 0.00228571
R30270 VSS.n11391 VSS.n11273 0.00228571
R30271 VSS.n11453 VSS.n11225 0.00228571
R30272 VSS.n11453 VSS.n11452 0.00228571
R30273 VSS.n11464 VSS.n11217 0.00228571
R30274 VSS.n11475 VSS.n11209 0.00228571
R30275 VSS.n11496 VSS.n11495 0.00228571
R30276 VSS.n11476 VSS.n11207 0.00228571
R30277 VSS.n11164 VSS.n11161 0.00228571
R30278 VSS.n11578 VSS.n11577 0.00228571
R30279 VSS.n11151 VSS.n11145 0.00228571
R30280 VSS.n11651 VSS.n11124 0.00228571
R30281 VSS.n11661 VSS.n11660 0.00228571
R30282 VSS.n11377 VSS.n11291 0.00228571
R30283 VSS.n11951 VSS.n11894 0.00228571
R30284 VSS.n11882 VSS.n11881 0.00228571
R30285 VSS.n11983 VSS.n11865 0.00228571
R30286 VSS.n12045 VSS.n11817 0.00228571
R30287 VSS.n12045 VSS.n12044 0.00228571
R30288 VSS.n12056 VSS.n11809 0.00228571
R30289 VSS.n12067 VSS.n11801 0.00228571
R30290 VSS.n12088 VSS.n12087 0.00228571
R30291 VSS.n12068 VSS.n11799 0.00228571
R30292 VSS.n11756 VSS.n11753 0.00228571
R30293 VSS.n12170 VSS.n12169 0.00228571
R30294 VSS.n11743 VSS.n11737 0.00228571
R30295 VSS.n12243 VSS.n11716 0.00228571
R30296 VSS.n12253 VSS.n12252 0.00228571
R30297 VSS.n11969 VSS.n11883 0.00228571
R30298 VSS.n12543 VSS.n12486 0.00228571
R30299 VSS.n12474 VSS.n12473 0.00228571
R30300 VSS.n12575 VSS.n12457 0.00228571
R30301 VSS.n12637 VSS.n12409 0.00228571
R30302 VSS.n12637 VSS.n12636 0.00228571
R30303 VSS.n12648 VSS.n12401 0.00228571
R30304 VSS.n12659 VSS.n12393 0.00228571
R30305 VSS.n12680 VSS.n12679 0.00228571
R30306 VSS.n12660 VSS.n12391 0.00228571
R30307 VSS.n12348 VSS.n12345 0.00228571
R30308 VSS.n12762 VSS.n12761 0.00228571
R30309 VSS.n12335 VSS.n12329 0.00228571
R30310 VSS.n12835 VSS.n12308 0.00228571
R30311 VSS.n12845 VSS.n12844 0.00228571
R30312 VSS.n12561 VSS.n12475 0.00228571
R30313 VSS.n13135 VSS.n13078 0.00228571
R30314 VSS.n13066 VSS.n13065 0.00228571
R30315 VSS.n13167 VSS.n13049 0.00228571
R30316 VSS.n13229 VSS.n13001 0.00228571
R30317 VSS.n13229 VSS.n13228 0.00228571
R30318 VSS.n13240 VSS.n12993 0.00228571
R30319 VSS.n13251 VSS.n12985 0.00228571
R30320 VSS.n13272 VSS.n13271 0.00228571
R30321 VSS.n13252 VSS.n12983 0.00228571
R30322 VSS.n12940 VSS.n12937 0.00228571
R30323 VSS.n13354 VSS.n13353 0.00228571
R30324 VSS.n12927 VSS.n12921 0.00228571
R30325 VSS.n13427 VSS.n12900 0.00228571
R30326 VSS.n13437 VSS.n13436 0.00228571
R30327 VSS.n13153 VSS.n13067 0.00228571
R30328 VSS.n13727 VSS.n13670 0.00228571
R30329 VSS.n13658 VSS.n13657 0.00228571
R30330 VSS.n13759 VSS.n13641 0.00228571
R30331 VSS.n13821 VSS.n13593 0.00228571
R30332 VSS.n13821 VSS.n13820 0.00228571
R30333 VSS.n13832 VSS.n13585 0.00228571
R30334 VSS.n13843 VSS.n13577 0.00228571
R30335 VSS.n13864 VSS.n13863 0.00228571
R30336 VSS.n13844 VSS.n13575 0.00228571
R30337 VSS.n13532 VSS.n13529 0.00228571
R30338 VSS.n13946 VSS.n13945 0.00228571
R30339 VSS.n13519 VSS.n13513 0.00228571
R30340 VSS.n14019 VSS.n13492 0.00228571
R30341 VSS.n14029 VSS.n14028 0.00228571
R30342 VSS.n13745 VSS.n13659 0.00228571
R30343 VSS.n14319 VSS.n14262 0.00228571
R30344 VSS.n14250 VSS.n14249 0.00228571
R30345 VSS.n14351 VSS.n14233 0.00228571
R30346 VSS.n14413 VSS.n14185 0.00228571
R30347 VSS.n14413 VSS.n14412 0.00228571
R30348 VSS.n14424 VSS.n14177 0.00228571
R30349 VSS.n14435 VSS.n14169 0.00228571
R30350 VSS.n14456 VSS.n14455 0.00228571
R30351 VSS.n14436 VSS.n14167 0.00228571
R30352 VSS.n14124 VSS.n14121 0.00228571
R30353 VSS.n14538 VSS.n14537 0.00228571
R30354 VSS.n14111 VSS.n14105 0.00228571
R30355 VSS.n14611 VSS.n14084 0.00228571
R30356 VSS.n14621 VSS.n14620 0.00228571
R30357 VSS.n14337 VSS.n14251 0.00228571
R30358 VSS.n14911 VSS.n14854 0.00228571
R30359 VSS.n14842 VSS.n14841 0.00228571
R30360 VSS.n14943 VSS.n14825 0.00228571
R30361 VSS.n15005 VSS.n14777 0.00228571
R30362 VSS.n15005 VSS.n15004 0.00228571
R30363 VSS.n15016 VSS.n14769 0.00228571
R30364 VSS.n15027 VSS.n14761 0.00228571
R30365 VSS.n15048 VSS.n15047 0.00228571
R30366 VSS.n15028 VSS.n14759 0.00228571
R30367 VSS.n14716 VSS.n14713 0.00228571
R30368 VSS.n15130 VSS.n15129 0.00228571
R30369 VSS.n14703 VSS.n14697 0.00228571
R30370 VSS.n15203 VSS.n14676 0.00228571
R30371 VSS.n15213 VSS.n15212 0.00228571
R30372 VSS.n14929 VSS.n14843 0.00228571
R30373 VSS.n15503 VSS.n15446 0.00228571
R30374 VSS.n15434 VSS.n15433 0.00228571
R30375 VSS.n15535 VSS.n15417 0.00228571
R30376 VSS.n15597 VSS.n15369 0.00228571
R30377 VSS.n15597 VSS.n15596 0.00228571
R30378 VSS.n15608 VSS.n15361 0.00228571
R30379 VSS.n15619 VSS.n15353 0.00228571
R30380 VSS.n15640 VSS.n15639 0.00228571
R30381 VSS.n15620 VSS.n15351 0.00228571
R30382 VSS.n15308 VSS.n15305 0.00228571
R30383 VSS.n15722 VSS.n15721 0.00228571
R30384 VSS.n15295 VSS.n15289 0.00228571
R30385 VSS.n15795 VSS.n15268 0.00228571
R30386 VSS.n15805 VSS.n15804 0.00228571
R30387 VSS.n15521 VSS.n15435 0.00228571
R30388 VSS.n6611 VSS.n6554 0.00228571
R30389 VSS.n6542 VSS.n6541 0.00228571
R30390 VSS.n6643 VSS.n6525 0.00228571
R30391 VSS.n6753 VSS.n6684 0.00228571
R30392 VSS.n6758 VSS.n6753 0.00228571
R30393 VSS.n6754 VSS.n6733 0.00228571
R30394 VSS.n15948 VSS.n6690 0.00228571
R30395 VSS.n6785 VSS.n6784 0.00228571
R30396 VSS.n15947 VSS.n15946 0.00228571
R30397 VSS.n15905 VSS.n15904 0.00228571
R30398 VSS.n15894 VSS.n15893 0.00228571
R30399 VSS.n6870 VSS.n6856 0.00228571
R30400 VSS.n6898 VSS.n6895 0.00228571
R30401 VSS.n15853 VSS.n6907 0.00228571
R30402 VSS.n6629 VSS.n6543 0.00228571
R30403 VSS.n7215 VSS.n7149 0.00228571
R30404 VSS.n7233 VSS.n7133 0.00228571
R30405 VSS.n7247 VSS.n7246 0.00228571
R30406 VSS.n7309 VSS.n7080 0.00228571
R30407 VSS.n7309 VSS.n7308 0.00228571
R30408 VSS.n7320 VSS.n7072 0.00228571
R30409 VSS.n7331 VSS.n7064 0.00228571
R30410 VSS.n7352 VSS.n7351 0.00228571
R30411 VSS.n7332 VSS.n7062 0.00228571
R30412 VSS.n7019 VSS.n7016 0.00228571
R30413 VSS.n7434 VSS.n7433 0.00228571
R30414 VSS.n7006 VSS.n7000 0.00228571
R30415 VSS.n7507 VSS.n6979 0.00228571
R30416 VSS.n7517 VSS.n7516 0.00228571
R30417 VSS.n7232 VSS.n7134 0.00228571
R30418 VSS.n370 VSS.n369 0.00228571
R30419 VSS.n428 VSS.n427 0.00228571
R30420 VSS.n388 VSS.n387 0.00228571
R30421 VSS.n18621 VSS.n178 0.00228571
R30422 VSS.n18621 VSS.n18620 0.00228571
R30423 VSS.n18632 VSS.n170 0.00228571
R30424 VSS.n18643 VSS.n162 0.00228571
R30425 VSS.n18664 VSS.n18663 0.00228571
R30426 VSS.n18644 VSS.n160 0.00228571
R30427 VSS.n117 VSS.n114 0.00228571
R30428 VSS.n18746 VSS.n18745 0.00228571
R30429 VSS.n104 VSS.n98 0.00228571
R30430 VSS.n18819 VSS.n77 0.00228571
R30431 VSS.n18829 VSS.n18828 0.00228571
R30432 VSS.n429 VSS.n311 0.00228571
R30433 VSS.n576 VSS.n504 0.00228571
R30434 VSS.n581 VSS.n576 0.00228571
R30435 VSS.n577 VSS.n553 0.00228571
R30436 VSS.n862 VSS.n510 0.00228571
R30437 VSS.n608 VSS.n607 0.00228571
R30438 VSS.n861 VSS.n860 0.00228571
R30439 VSS.n819 VSS.n818 0.00228571
R30440 VSS.n808 VSS.n807 0.00228571
R30441 VSS.n693 VSS.n679 0.00228571
R30442 VSS.n721 VSS.n718 0.00228571
R30443 VSS.n767 VSS.n730 0.00228571
R30444 VSS.n994 VSS.n477 0.00228571
R30445 VSS.n17933 VSS.n17932 0.00228571
R30446 VSS.n17922 VSS.n17921 0.00228571
R30447 VSS.n1352 VSS.n1338 0.00228571
R30448 VSS.n1380 VSS.n1377 0.00228571
R30449 VSS.n17881 VSS.n1389 0.00228571
R30450 VSS.n18038 VSS.n18037 0.00217857
R30451 VSS.n18036 VSS.n1027 0.00217857
R30452 VSS.n18007 VSS.n1051 0.00217857
R30453 VSS.n18006 VSS.n1057 0.00217857
R30454 VSS.n17020 VSS.n16996 0.00217857
R30455 VSS.n17021 VSS.n16982 0.00217857
R30456 VSS.n17091 VSS.n16944 0.00217857
R30457 VSS.n17092 VSS.n16932 0.00217857
R30458 VSS.n17514 VSS.n17490 0.00217857
R30459 VSS.n17515 VSS.n17470 0.00217857
R30460 VSS.n17576 VSS.n17439 0.00217857
R30461 VSS.n17577 VSS.n17421 0.00217857
R30462 VSS.n17612 VSS.n17410 0.00217857
R30463 VSS.n17613 VSS.n17396 0.00217857
R30464 VSS.n17683 VSS.n17358 0.00217857
R30465 VSS.n17684 VSS.n17346 0.00217857
R30466 VSS.n18091 VSS.n282 0.00217857
R30467 VSS.n18092 VSS.n262 0.00217857
R30468 VSS.n18153 VSS.n231 0.00217857
R30469 VSS.n18154 VSS.n213 0.00217857
R30470 VSS.n18578 VSS.n18577 0.00217857
R30471 VSS.n18576 VSS.n18179 0.00217857
R30472 VSS.n18547 VSS.n18202 0.00217857
R30473 VSS.n18546 VSS.n18208 0.00217857
R30474 VSS.n9662 VSS.n9460 0.00217857
R30475 VSS.n9663 VSS.n9446 0.00217857
R30476 VSS.n9733 VSS.n9408 0.00217857
R30477 VSS.n9734 VSS.n9396 0.00217857
R30478 VSS.n16500 VSS.n16477 0.00217857
R30479 VSS.n16501 VSS.n16465 0.00217857
R30480 VSS.n16572 VSS.n16425 0.00217857
R30481 VSS.n16573 VSS.n16413 0.00217857
R30482 VSS.n16605 VSS.n16402 0.00217857
R30483 VSS.n16606 VSS.n16388 0.00217857
R30484 VSS.n16676 VSS.n16350 0.00217857
R30485 VSS.n16677 VSS.n16338 0.00217857
R30486 VSS.n1665 VSS.n1642 0.00217857
R30487 VSS.n1666 VSS.n1630 0.00217857
R30488 VSS.n1737 VSS.n1590 0.00217857
R30489 VSS.n1738 VSS.n1578 0.00217857
R30490 VSS.n16012 VSS.n1574 0.00217857
R30491 VSS.n16013 VSS.n1560 0.00217857
R30492 VSS.n16083 VSS.n1522 0.00217857
R30493 VSS.n16084 VSS.n1510 0.00217857
R30494 VSS.n1856 VSS.n1832 0.00217857
R30495 VSS.n1857 VSS.n1812 0.00217857
R30496 VSS.n1918 VSS.n1781 0.00217857
R30497 VSS.n1919 VSS.n1763 0.00217857
R30498 VSS.n2343 VSS.n2342 0.00217857
R30499 VSS.n2341 VSS.n1944 0.00217857
R30500 VSS.n2312 VSS.n1967 0.00217857
R30501 VSS.n2311 VSS.n1973 0.00217857
R30502 VSS.n3055 VSS.n3031 0.00217857
R30503 VSS.n3056 VSS.n3011 0.00217857
R30504 VSS.n3117 VSS.n2980 0.00217857
R30505 VSS.n3118 VSS.n2962 0.00217857
R30506 VSS.n3153 VSS.n2951 0.00217857
R30507 VSS.n3154 VSS.n2937 0.00217857
R30508 VSS.n3224 VSS.n2899 0.00217857
R30509 VSS.n3225 VSS.n2887 0.00217857
R30510 VSS.n3647 VSS.n3623 0.00217857
R30511 VSS.n3648 VSS.n3603 0.00217857
R30512 VSS.n3709 VSS.n3572 0.00217857
R30513 VSS.n3710 VSS.n3554 0.00217857
R30514 VSS.n3745 VSS.n3543 0.00217857
R30515 VSS.n3746 VSS.n3529 0.00217857
R30516 VSS.n3816 VSS.n3491 0.00217857
R30517 VSS.n3817 VSS.n3479 0.00217857
R30518 VSS.n4239 VSS.n4215 0.00217857
R30519 VSS.n4240 VSS.n4195 0.00217857
R30520 VSS.n4301 VSS.n4164 0.00217857
R30521 VSS.n4302 VSS.n4146 0.00217857
R30522 VSS.n4337 VSS.n4135 0.00217857
R30523 VSS.n4338 VSS.n4121 0.00217857
R30524 VSS.n4408 VSS.n4083 0.00217857
R30525 VSS.n4409 VSS.n4071 0.00217857
R30526 VSS.n4831 VSS.n4807 0.00217857
R30527 VSS.n4832 VSS.n4787 0.00217857
R30528 VSS.n4893 VSS.n4756 0.00217857
R30529 VSS.n4894 VSS.n4738 0.00217857
R30530 VSS.n4929 VSS.n4727 0.00217857
R30531 VSS.n4930 VSS.n4713 0.00217857
R30532 VSS.n5000 VSS.n4675 0.00217857
R30533 VSS.n5001 VSS.n4663 0.00217857
R30534 VSS.n2452 VSS.n2428 0.00217857
R30535 VSS.n2453 VSS.n2408 0.00217857
R30536 VSS.n2514 VSS.n2377 0.00217857
R30537 VSS.n2515 VSS.n2359 0.00217857
R30538 VSS.n5308 VSS.n5307 0.00217857
R30539 VSS.n5306 VSS.n2540 0.00217857
R30540 VSS.n5277 VSS.n2563 0.00217857
R30541 VSS.n5276 VSS.n2569 0.00217857
R30542 VSS.n5413 VSS.n5389 0.00217857
R30543 VSS.n5414 VSS.n5369 0.00217857
R30544 VSS.n5475 VSS.n5338 0.00217857
R30545 VSS.n5476 VSS.n5320 0.00217857
R30546 VSS.n5881 VSS.n5880 0.00217857
R30547 VSS.n5879 VSS.n5501 0.00217857
R30548 VSS.n5850 VSS.n5524 0.00217857
R30549 VSS.n5849 VSS.n5530 0.00217857
R30550 VSS.n5986 VSS.n5962 0.00217857
R30551 VSS.n5987 VSS.n5942 0.00217857
R30552 VSS.n6048 VSS.n5911 0.00217857
R30553 VSS.n6049 VSS.n5893 0.00217857
R30554 VSS.n6473 VSS.n6472 0.00217857
R30555 VSS.n6471 VSS.n6074 0.00217857
R30556 VSS.n6442 VSS.n6097 0.00217857
R30557 VSS.n6441 VSS.n6103 0.00217857
R30558 VSS.n7788 VSS.n7764 0.00217857
R30559 VSS.n7789 VSS.n7744 0.00217857
R30560 VSS.n7850 VSS.n7713 0.00217857
R30561 VSS.n7851 VSS.n7695 0.00217857
R30562 VSS.n7886 VSS.n7684 0.00217857
R30563 VSS.n7887 VSS.n7670 0.00217857
R30564 VSS.n7957 VSS.n7632 0.00217857
R30565 VSS.n7958 VSS.n7620 0.00217857
R30566 VSS.n8380 VSS.n8356 0.00217857
R30567 VSS.n8381 VSS.n8336 0.00217857
R30568 VSS.n8442 VSS.n8305 0.00217857
R30569 VSS.n8443 VSS.n8287 0.00217857
R30570 VSS.n8478 VSS.n8276 0.00217857
R30571 VSS.n8479 VSS.n8262 0.00217857
R30572 VSS.n8549 VSS.n8224 0.00217857
R30573 VSS.n8550 VSS.n8212 0.00217857
R30574 VSS.n8972 VSS.n8948 0.00217857
R30575 VSS.n8973 VSS.n8928 0.00217857
R30576 VSS.n9034 VSS.n8897 0.00217857
R30577 VSS.n9035 VSS.n8879 0.00217857
R30578 VSS.n9070 VSS.n8868 0.00217857
R30579 VSS.n9071 VSS.n8854 0.00217857
R30580 VSS.n9141 VSS.n8816 0.00217857
R30581 VSS.n9142 VSS.n8804 0.00217857
R30582 VSS.n10156 VSS.n10132 0.00217857
R30583 VSS.n10157 VSS.n10112 0.00217857
R30584 VSS.n10218 VSS.n10081 0.00217857
R30585 VSS.n10219 VSS.n10063 0.00217857
R30586 VSS.n10254 VSS.n10052 0.00217857
R30587 VSS.n10255 VSS.n10038 0.00217857
R30588 VSS.n10325 VSS.n10000 0.00217857
R30589 VSS.n10326 VSS.n9988 0.00217857
R30590 VSS.n10748 VSS.n10724 0.00217857
R30591 VSS.n10749 VSS.n10704 0.00217857
R30592 VSS.n10810 VSS.n10673 0.00217857
R30593 VSS.n10811 VSS.n10655 0.00217857
R30594 VSS.n10846 VSS.n10644 0.00217857
R30595 VSS.n10847 VSS.n10630 0.00217857
R30596 VSS.n10917 VSS.n10592 0.00217857
R30597 VSS.n10918 VSS.n10580 0.00217857
R30598 VSS.n11340 VSS.n11316 0.00217857
R30599 VSS.n11341 VSS.n11296 0.00217857
R30600 VSS.n11402 VSS.n11265 0.00217857
R30601 VSS.n11403 VSS.n11247 0.00217857
R30602 VSS.n11438 VSS.n11236 0.00217857
R30603 VSS.n11439 VSS.n11222 0.00217857
R30604 VSS.n11509 VSS.n11184 0.00217857
R30605 VSS.n11510 VSS.n11172 0.00217857
R30606 VSS.n11932 VSS.n11908 0.00217857
R30607 VSS.n11933 VSS.n11888 0.00217857
R30608 VSS.n11994 VSS.n11857 0.00217857
R30609 VSS.n11995 VSS.n11839 0.00217857
R30610 VSS.n12030 VSS.n11828 0.00217857
R30611 VSS.n12031 VSS.n11814 0.00217857
R30612 VSS.n12101 VSS.n11776 0.00217857
R30613 VSS.n12102 VSS.n11764 0.00217857
R30614 VSS.n12524 VSS.n12500 0.00217857
R30615 VSS.n12525 VSS.n12480 0.00217857
R30616 VSS.n12586 VSS.n12449 0.00217857
R30617 VSS.n12587 VSS.n12431 0.00217857
R30618 VSS.n12622 VSS.n12420 0.00217857
R30619 VSS.n12623 VSS.n12406 0.00217857
R30620 VSS.n12693 VSS.n12368 0.00217857
R30621 VSS.n12694 VSS.n12356 0.00217857
R30622 VSS.n13116 VSS.n13092 0.00217857
R30623 VSS.n13117 VSS.n13072 0.00217857
R30624 VSS.n13178 VSS.n13041 0.00217857
R30625 VSS.n13179 VSS.n13023 0.00217857
R30626 VSS.n13214 VSS.n13012 0.00217857
R30627 VSS.n13215 VSS.n12998 0.00217857
R30628 VSS.n13285 VSS.n12960 0.00217857
R30629 VSS.n13286 VSS.n12948 0.00217857
R30630 VSS.n13708 VSS.n13684 0.00217857
R30631 VSS.n13709 VSS.n13664 0.00217857
R30632 VSS.n13770 VSS.n13633 0.00217857
R30633 VSS.n13771 VSS.n13615 0.00217857
R30634 VSS.n13806 VSS.n13604 0.00217857
R30635 VSS.n13807 VSS.n13590 0.00217857
R30636 VSS.n13877 VSS.n13552 0.00217857
R30637 VSS.n13878 VSS.n13540 0.00217857
R30638 VSS.n14300 VSS.n14276 0.00217857
R30639 VSS.n14301 VSS.n14256 0.00217857
R30640 VSS.n14362 VSS.n14225 0.00217857
R30641 VSS.n14363 VSS.n14207 0.00217857
R30642 VSS.n14398 VSS.n14196 0.00217857
R30643 VSS.n14399 VSS.n14182 0.00217857
R30644 VSS.n14469 VSS.n14144 0.00217857
R30645 VSS.n14470 VSS.n14132 0.00217857
R30646 VSS.n14892 VSS.n14868 0.00217857
R30647 VSS.n14893 VSS.n14848 0.00217857
R30648 VSS.n14954 VSS.n14817 0.00217857
R30649 VSS.n14955 VSS.n14799 0.00217857
R30650 VSS.n14990 VSS.n14788 0.00217857
R30651 VSS.n14991 VSS.n14774 0.00217857
R30652 VSS.n15061 VSS.n14736 0.00217857
R30653 VSS.n15062 VSS.n14724 0.00217857
R30654 VSS.n15484 VSS.n15460 0.00217857
R30655 VSS.n15485 VSS.n15440 0.00217857
R30656 VSS.n15546 VSS.n15409 0.00217857
R30657 VSS.n15547 VSS.n15391 0.00217857
R30658 VSS.n15582 VSS.n15380 0.00217857
R30659 VSS.n15583 VSS.n15366 0.00217857
R30660 VSS.n15653 VSS.n15328 0.00217857
R30661 VSS.n15654 VSS.n15316 0.00217857
R30662 VSS.n6592 VSS.n6568 0.00217857
R30663 VSS.n6593 VSS.n6548 0.00217857
R30664 VSS.n6654 VSS.n6517 0.00217857
R30665 VSS.n6655 VSS.n6499 0.00217857
R30666 VSS.n15961 VSS.n15960 0.00217857
R30667 VSS.n15959 VSS.n6680 0.00217857
R30668 VSS.n15930 VSS.n6703 0.00217857
R30669 VSS.n15929 VSS.n6709 0.00217857
R30670 VSS.n7189 VSS.n7166 0.00217857
R30671 VSS.n7190 VSS.n7154 0.00217857
R30672 VSS.n7261 VSS.n7114 0.00217857
R30673 VSS.n7262 VSS.n7102 0.00217857
R30674 VSS.n7294 VSS.n7091 0.00217857
R30675 VSS.n7295 VSS.n7077 0.00217857
R30676 VSS.n7365 VSS.n7039 0.00217857
R30677 VSS.n7366 VSS.n7027 0.00217857
R30678 VSS.n447 VSS.n446 0.00217857
R30679 VSS.n445 VSS.n294 0.00217857
R30680 VSS.n416 VSS.n318 0.00217857
R30681 VSS.n415 VSS.n193 0.00217857
R30682 VSS.n18606 VSS.n189 0.00217857
R30683 VSS.n18607 VSS.n175 0.00217857
R30684 VSS.n18677 VSS.n137 0.00217857
R30685 VSS.n18678 VSS.n125 0.00217857
R30686 VSS.n1012 VSS.n1011 0.00217857
R30687 VSS.n1010 VSS.n460 0.00217857
R30688 VSS.n981 VSS.n484 0.00217857
R30689 VSS.n980 VSS.n490 0.00217857
R30690 VSS.n874 VSS.n495 0.00217857
R30691 VSS.n873 VSS.n500 0.00217857
R30692 VSS.n844 VSS.n523 0.00217857
R30693 VSS.n843 VSS.n529 0.00217857
R30694 VSS.n17989 VSS.n17988 0.00217857
R30695 VSS.n17987 VSS.n1162 0.00217857
R30696 VSS.n17958 VSS.n1185 0.00217857
R30697 VSS.n17957 VSS.n1191 0.00217857
R30698 VSS.n9564 VSS.n9540 0.00216667
R30699 VSS.n9565 VSS.n9520 0.00216667
R30700 VSS.n9626 VSS.n9489 0.00216667
R30701 VSS.n9627 VSS.n9471 0.00216667
R30702 VSS.n1276 VSS.n1205 0.00139286
R30703 VSS.n1282 VSS.n1202 0.00139286
R30704 VSS.n895 VSS.n478 0.00139286
R30705 VSS.n961 VSS.n890 0.00139286
R30706 VSS.n967 VSS.n887 0.00139286
R30707 VSS.n17087 VSS.n16950 0.00139286
R30708 VSS.n17099 VSS.n16941 0.00139286
R30709 VSS.n1076 VSS.n1045 0.00139286
R30710 VSS.n1142 VSS.n1071 0.00139286
R30711 VSS.n1148 VSS.n1068 0.00139286
R30712 VSS.n1043 VSS.n1040 0.00139286
R30713 VSS.n17201 VSS.n17196 0.00139286
R30714 VSS.n17205 VSS.n17204 0.00139286
R30715 VSS.n17197 VSS.n16900 0.00139286
R30716 VSS.n17206 VSS.n17195 0.00139286
R30717 VSS.n17679 VSS.n17364 0.00139286
R30718 VSS.n17691 VSS.n17355 0.00139286
R30719 VSS.n17554 VSS.n17553 0.00139286
R30720 VSS.n17587 VSS.n17586 0.00139286
R30721 VSS.n17438 VSS.n17434 0.00139286
R30722 VSS.n17552 VSS.n17462 0.00139286
R30723 VSS.n17793 VSS.n17788 0.00139286
R30724 VSS.n17797 VSS.n17796 0.00139286
R30725 VSS.n17789 VSS.n17314 0.00139286
R30726 VSS.n17798 VSS.n17787 0.00139286
R30727 VSS.n18131 VSS.n18130 0.00139286
R30728 VSS.n18164 VSS.n18163 0.00139286
R30729 VSS.n230 VSS.n226 0.00139286
R30730 VSS.n18293 VSS.n18222 0.00139286
R30731 VSS.n18299 VSS.n18219 0.00139286
R30732 VSS.n18406 VSS.n18394 0.00139286
R30733 VSS.n18409 VSS.n18388 0.00139286
R30734 VSS.n18397 VSS.n18395 0.00139286
R30735 VSS.n18411 VSS.n18410 0.00139286
R30736 VSS.n18129 VSS.n254 0.00139286
R30737 VSS.n9604 VSS.n9603 0.00139286
R30738 VSS.n9637 VSS.n9636 0.00139286
R30739 VSS.n9488 VSS.n9484 0.00139286
R30740 VSS.n9729 VSS.n9414 0.00139286
R30741 VSS.n9741 VSS.n9405 0.00139286
R30742 VSS.n9843 VSS.n9838 0.00139286
R30743 VSS.n9847 VSS.n9846 0.00139286
R30744 VSS.n9839 VSS.n9364 0.00139286
R30745 VSS.n9848 VSS.n9837 0.00139286
R30746 VSS.n9602 VSS.n9512 0.00139286
R30747 VSS.n16536 VSS.n16452 0.00139286
R30748 VSS.n16568 VSS.n16431 0.00139286
R30749 VSS.n16580 VSS.n16422 0.00139286
R30750 VSS.n16672 VSS.n16356 0.00139286
R30751 VSS.n16684 VSS.n16347 0.00139286
R30752 VSS.n16786 VSS.n16781 0.00139286
R30753 VSS.n16790 VSS.n16789 0.00139286
R30754 VSS.n16782 VSS.n16306 0.00139286
R30755 VSS.n16791 VSS.n16780 0.00139286
R30756 VSS.n16451 VSS.n16449 0.00139286
R30757 VSS.n1701 VSS.n1617 0.00139286
R30758 VSS.n1733 VSS.n1596 0.00139286
R30759 VSS.n1745 VSS.n1587 0.00139286
R30760 VSS.n16079 VSS.n1528 0.00139286
R30761 VSS.n16091 VSS.n1519 0.00139286
R30762 VSS.n16193 VSS.n16188 0.00139286
R30763 VSS.n16197 VSS.n16196 0.00139286
R30764 VSS.n16189 VSS.n1478 0.00139286
R30765 VSS.n16198 VSS.n16187 0.00139286
R30766 VSS.n1616 VSS.n1614 0.00139286
R30767 VSS.n1896 VSS.n1895 0.00139286
R30768 VSS.n1929 VSS.n1928 0.00139286
R30769 VSS.n1780 VSS.n1776 0.00139286
R30770 VSS.n2058 VSS.n1987 0.00139286
R30771 VSS.n2064 VSS.n1984 0.00139286
R30772 VSS.n2183 VSS.n2181 0.00139286
R30773 VSS.n2253 VSS.n2252 0.00139286
R30774 VSS.n2182 VSS.n2130 0.00139286
R30775 VSS.n2254 VSS.n2154 0.00139286
R30776 VSS.n1894 VSS.n1804 0.00139286
R30777 VSS.n3095 VSS.n3094 0.00139286
R30778 VSS.n3128 VSS.n3127 0.00139286
R30779 VSS.n2979 VSS.n2975 0.00139286
R30780 VSS.n3220 VSS.n2905 0.00139286
R30781 VSS.n3232 VSS.n2896 0.00139286
R30782 VSS.n3334 VSS.n3329 0.00139286
R30783 VSS.n3338 VSS.n3337 0.00139286
R30784 VSS.n3330 VSS.n2855 0.00139286
R30785 VSS.n3339 VSS.n3328 0.00139286
R30786 VSS.n3093 VSS.n3003 0.00139286
R30787 VSS.n3687 VSS.n3686 0.00139286
R30788 VSS.n3720 VSS.n3719 0.00139286
R30789 VSS.n3571 VSS.n3567 0.00139286
R30790 VSS.n3812 VSS.n3497 0.00139286
R30791 VSS.n3824 VSS.n3488 0.00139286
R30792 VSS.n3926 VSS.n3921 0.00139286
R30793 VSS.n3930 VSS.n3929 0.00139286
R30794 VSS.n3922 VSS.n3447 0.00139286
R30795 VSS.n3931 VSS.n3920 0.00139286
R30796 VSS.n3685 VSS.n3595 0.00139286
R30797 VSS.n4279 VSS.n4278 0.00139286
R30798 VSS.n4312 VSS.n4311 0.00139286
R30799 VSS.n4163 VSS.n4159 0.00139286
R30800 VSS.n4404 VSS.n4089 0.00139286
R30801 VSS.n4416 VSS.n4080 0.00139286
R30802 VSS.n4518 VSS.n4513 0.00139286
R30803 VSS.n4522 VSS.n4521 0.00139286
R30804 VSS.n4514 VSS.n4039 0.00139286
R30805 VSS.n4523 VSS.n4512 0.00139286
R30806 VSS.n4277 VSS.n4187 0.00139286
R30807 VSS.n4871 VSS.n4870 0.00139286
R30808 VSS.n4904 VSS.n4903 0.00139286
R30809 VSS.n4755 VSS.n4751 0.00139286
R30810 VSS.n4996 VSS.n4681 0.00139286
R30811 VSS.n5008 VSS.n4672 0.00139286
R30812 VSS.n5110 VSS.n5105 0.00139286
R30813 VSS.n5114 VSS.n5113 0.00139286
R30814 VSS.n5106 VSS.n4631 0.00139286
R30815 VSS.n5115 VSS.n5104 0.00139286
R30816 VSS.n4869 VSS.n4779 0.00139286
R30817 VSS.n2492 VSS.n2491 0.00139286
R30818 VSS.n2525 VSS.n2524 0.00139286
R30819 VSS.n2376 VSS.n2372 0.00139286
R30820 VSS.n2654 VSS.n2583 0.00139286
R30821 VSS.n2660 VSS.n2580 0.00139286
R30822 VSS.n2779 VSS.n2777 0.00139286
R30823 VSS.n5218 VSS.n5217 0.00139286
R30824 VSS.n2778 VSS.n2726 0.00139286
R30825 VSS.n5219 VSS.n2750 0.00139286
R30826 VSS.n2490 VSS.n2400 0.00139286
R30827 VSS.n5453 VSS.n5452 0.00139286
R30828 VSS.n5486 VSS.n5485 0.00139286
R30829 VSS.n5337 VSS.n5333 0.00139286
R30830 VSS.n5615 VSS.n5544 0.00139286
R30831 VSS.n5621 VSS.n5541 0.00139286
R30832 VSS.n5753 VSS.n5751 0.00139286
R30833 VSS.n5791 VSS.n5790 0.00139286
R30834 VSS.n5752 VSS.n5687 0.00139286
R30835 VSS.n5792 VSS.n5711 0.00139286
R30836 VSS.n5451 VSS.n5361 0.00139286
R30837 VSS.n6026 VSS.n6025 0.00139286
R30838 VSS.n6059 VSS.n6058 0.00139286
R30839 VSS.n5910 VSS.n5906 0.00139286
R30840 VSS.n6188 VSS.n6117 0.00139286
R30841 VSS.n6194 VSS.n6114 0.00139286
R30842 VSS.n6313 VSS.n6311 0.00139286
R30843 VSS.n6383 VSS.n6382 0.00139286
R30844 VSS.n6312 VSS.n6260 0.00139286
R30845 VSS.n6384 VSS.n6284 0.00139286
R30846 VSS.n6024 VSS.n5934 0.00139286
R30847 VSS.n7828 VSS.n7827 0.00139286
R30848 VSS.n7861 VSS.n7860 0.00139286
R30849 VSS.n7712 VSS.n7708 0.00139286
R30850 VSS.n7953 VSS.n7638 0.00139286
R30851 VSS.n7965 VSS.n7629 0.00139286
R30852 VSS.n8067 VSS.n8062 0.00139286
R30853 VSS.n8071 VSS.n8070 0.00139286
R30854 VSS.n8063 VSS.n7588 0.00139286
R30855 VSS.n8072 VSS.n8061 0.00139286
R30856 VSS.n7826 VSS.n7736 0.00139286
R30857 VSS.n8420 VSS.n8419 0.00139286
R30858 VSS.n8453 VSS.n8452 0.00139286
R30859 VSS.n8304 VSS.n8300 0.00139286
R30860 VSS.n8545 VSS.n8230 0.00139286
R30861 VSS.n8557 VSS.n8221 0.00139286
R30862 VSS.n8659 VSS.n8654 0.00139286
R30863 VSS.n8663 VSS.n8662 0.00139286
R30864 VSS.n8655 VSS.n8180 0.00139286
R30865 VSS.n8664 VSS.n8653 0.00139286
R30866 VSS.n8418 VSS.n8328 0.00139286
R30867 VSS.n9012 VSS.n9011 0.00139286
R30868 VSS.n9045 VSS.n9044 0.00139286
R30869 VSS.n8896 VSS.n8892 0.00139286
R30870 VSS.n9137 VSS.n8822 0.00139286
R30871 VSS.n9149 VSS.n8813 0.00139286
R30872 VSS.n9251 VSS.n9246 0.00139286
R30873 VSS.n9255 VSS.n9254 0.00139286
R30874 VSS.n9247 VSS.n8772 0.00139286
R30875 VSS.n9256 VSS.n9245 0.00139286
R30876 VSS.n9010 VSS.n8920 0.00139286
R30877 VSS.n10196 VSS.n10195 0.00139286
R30878 VSS.n10229 VSS.n10228 0.00139286
R30879 VSS.n10080 VSS.n10076 0.00139286
R30880 VSS.n10321 VSS.n10006 0.00139286
R30881 VSS.n10333 VSS.n9997 0.00139286
R30882 VSS.n10435 VSS.n10430 0.00139286
R30883 VSS.n10439 VSS.n10438 0.00139286
R30884 VSS.n10431 VSS.n9956 0.00139286
R30885 VSS.n10440 VSS.n10429 0.00139286
R30886 VSS.n10194 VSS.n10104 0.00139286
R30887 VSS.n10788 VSS.n10787 0.00139286
R30888 VSS.n10821 VSS.n10820 0.00139286
R30889 VSS.n10672 VSS.n10668 0.00139286
R30890 VSS.n10913 VSS.n10598 0.00139286
R30891 VSS.n10925 VSS.n10589 0.00139286
R30892 VSS.n11027 VSS.n11022 0.00139286
R30893 VSS.n11031 VSS.n11030 0.00139286
R30894 VSS.n11023 VSS.n10548 0.00139286
R30895 VSS.n11032 VSS.n11021 0.00139286
R30896 VSS.n10786 VSS.n10696 0.00139286
R30897 VSS.n11380 VSS.n11379 0.00139286
R30898 VSS.n11413 VSS.n11412 0.00139286
R30899 VSS.n11264 VSS.n11260 0.00139286
R30900 VSS.n11505 VSS.n11190 0.00139286
R30901 VSS.n11517 VSS.n11181 0.00139286
R30902 VSS.n11619 VSS.n11614 0.00139286
R30903 VSS.n11623 VSS.n11622 0.00139286
R30904 VSS.n11615 VSS.n11140 0.00139286
R30905 VSS.n11624 VSS.n11613 0.00139286
R30906 VSS.n11378 VSS.n11288 0.00139286
R30907 VSS.n11972 VSS.n11971 0.00139286
R30908 VSS.n12005 VSS.n12004 0.00139286
R30909 VSS.n11856 VSS.n11852 0.00139286
R30910 VSS.n12097 VSS.n11782 0.00139286
R30911 VSS.n12109 VSS.n11773 0.00139286
R30912 VSS.n12211 VSS.n12206 0.00139286
R30913 VSS.n12215 VSS.n12214 0.00139286
R30914 VSS.n12207 VSS.n11732 0.00139286
R30915 VSS.n12216 VSS.n12205 0.00139286
R30916 VSS.n11970 VSS.n11880 0.00139286
R30917 VSS.n12564 VSS.n12563 0.00139286
R30918 VSS.n12597 VSS.n12596 0.00139286
R30919 VSS.n12448 VSS.n12444 0.00139286
R30920 VSS.n12689 VSS.n12374 0.00139286
R30921 VSS.n12701 VSS.n12365 0.00139286
R30922 VSS.n12803 VSS.n12798 0.00139286
R30923 VSS.n12807 VSS.n12806 0.00139286
R30924 VSS.n12799 VSS.n12324 0.00139286
R30925 VSS.n12808 VSS.n12797 0.00139286
R30926 VSS.n12562 VSS.n12472 0.00139286
R30927 VSS.n13156 VSS.n13155 0.00139286
R30928 VSS.n13189 VSS.n13188 0.00139286
R30929 VSS.n13040 VSS.n13036 0.00139286
R30930 VSS.n13281 VSS.n12966 0.00139286
R30931 VSS.n13293 VSS.n12957 0.00139286
R30932 VSS.n13395 VSS.n13390 0.00139286
R30933 VSS.n13399 VSS.n13398 0.00139286
R30934 VSS.n13391 VSS.n12916 0.00139286
R30935 VSS.n13400 VSS.n13389 0.00139286
R30936 VSS.n13154 VSS.n13064 0.00139286
R30937 VSS.n13748 VSS.n13747 0.00139286
R30938 VSS.n13781 VSS.n13780 0.00139286
R30939 VSS.n13632 VSS.n13628 0.00139286
R30940 VSS.n13873 VSS.n13558 0.00139286
R30941 VSS.n13885 VSS.n13549 0.00139286
R30942 VSS.n13987 VSS.n13982 0.00139286
R30943 VSS.n13991 VSS.n13990 0.00139286
R30944 VSS.n13983 VSS.n13508 0.00139286
R30945 VSS.n13992 VSS.n13981 0.00139286
R30946 VSS.n13746 VSS.n13656 0.00139286
R30947 VSS.n14340 VSS.n14339 0.00139286
R30948 VSS.n14373 VSS.n14372 0.00139286
R30949 VSS.n14224 VSS.n14220 0.00139286
R30950 VSS.n14465 VSS.n14150 0.00139286
R30951 VSS.n14477 VSS.n14141 0.00139286
R30952 VSS.n14579 VSS.n14574 0.00139286
R30953 VSS.n14583 VSS.n14582 0.00139286
R30954 VSS.n14575 VSS.n14100 0.00139286
R30955 VSS.n14584 VSS.n14573 0.00139286
R30956 VSS.n14338 VSS.n14248 0.00139286
R30957 VSS.n14932 VSS.n14931 0.00139286
R30958 VSS.n14965 VSS.n14964 0.00139286
R30959 VSS.n14816 VSS.n14812 0.00139286
R30960 VSS.n15057 VSS.n14742 0.00139286
R30961 VSS.n15069 VSS.n14733 0.00139286
R30962 VSS.n15171 VSS.n15166 0.00139286
R30963 VSS.n15175 VSS.n15174 0.00139286
R30964 VSS.n15167 VSS.n14692 0.00139286
R30965 VSS.n15176 VSS.n15165 0.00139286
R30966 VSS.n14930 VSS.n14840 0.00139286
R30967 VSS.n15524 VSS.n15523 0.00139286
R30968 VSS.n15557 VSS.n15556 0.00139286
R30969 VSS.n15408 VSS.n15404 0.00139286
R30970 VSS.n15649 VSS.n15334 0.00139286
R30971 VSS.n15661 VSS.n15325 0.00139286
R30972 VSS.n15763 VSS.n15758 0.00139286
R30973 VSS.n15767 VSS.n15766 0.00139286
R30974 VSS.n15759 VSS.n15284 0.00139286
R30975 VSS.n15768 VSS.n15757 0.00139286
R30976 VSS.n15522 VSS.n15432 0.00139286
R30977 VSS.n6632 VSS.n6631 0.00139286
R30978 VSS.n6665 VSS.n6664 0.00139286
R30979 VSS.n6516 VSS.n6512 0.00139286
R30980 VSS.n6794 VSS.n6723 0.00139286
R30981 VSS.n6800 VSS.n6720 0.00139286
R30982 VSS.n6919 VSS.n6917 0.00139286
R30983 VSS.n15871 VSS.n15870 0.00139286
R30984 VSS.n6918 VSS.n6866 0.00139286
R30985 VSS.n15872 VSS.n6890 0.00139286
R30986 VSS.n6630 VSS.n6540 0.00139286
R30987 VSS.n7225 VSS.n7141 0.00139286
R30988 VSS.n7257 VSS.n7120 0.00139286
R30989 VSS.n7269 VSS.n7111 0.00139286
R30990 VSS.n7361 VSS.n7045 0.00139286
R30991 VSS.n7373 VSS.n7036 0.00139286
R30992 VSS.n7475 VSS.n7470 0.00139286
R30993 VSS.n7479 VSS.n7478 0.00139286
R30994 VSS.n7471 VSS.n6995 0.00139286
R30995 VSS.n7480 VSS.n7469 0.00139286
R30996 VSS.n7140 VSS.n7138 0.00139286
R30997 VSS.n378 VSS.n312 0.00139286
R30998 VSS.n395 VSS.n327 0.00139286
R30999 VSS.n406 VSS.n325 0.00139286
R31000 VSS.n18673 VSS.n143 0.00139286
R31001 VSS.n18685 VSS.n134 0.00139286
R31002 VSS.n18787 VSS.n18782 0.00139286
R31003 VSS.n18791 VSS.n18790 0.00139286
R31004 VSS.n18783 VSS.n93 0.00139286
R31005 VSS.n18792 VSS.n18781 0.00139286
R31006 VSS.n310 VSS.n307 0.00139286
R31007 VSS.n617 VSS.n543 0.00139286
R31008 VSS.n623 VSS.n540 0.00139286
R31009 VSS.n751 VSS.n749 0.00139286
R31010 VSS.n785 VSS.n784 0.00139286
R31011 VSS.n750 VSS.n689 0.00139286
R31012 VSS.n786 VSS.n713 0.00139286
R31013 VSS.n476 VSS.n473 0.00139286
R31014 VSS.n1401 VSS.n1399 0.00139286
R31015 VSS.n17899 VSS.n17898 0.00139286
R31016 VSS.n1400 VSS.n1348 0.00139286
R31017 VSS.n17900 VSS.n1372 0.00139286
R31018 VSS.n17865 VSS.n17864 0.00054824
R31019 VSS.n17273 VSS.n17272 0.00054824
R31020 VSS.n16859 VSS.n16858 0.00054824
R31021 VSS.n16266 VSS.n16265 0.00054824
R31022 VSS.n2220 VSS.n1438 0.00054824
R31023 VSS.n3407 VSS.n3406 0.00054824
R31024 VSS.n3999 VSS.n3998 0.00054824
R31025 VSS.n4591 VSS.n4590 0.00054824
R31026 VSS.n5183 VSS.n5182 0.00054824
R31027 VSS.n5185 VSS.n5184 0.00054824
R31028 VSS.n18889 VSS.n18888 0.00054824
R31029 VSS.n6350 VSS.n0 0.00054824
R31030 VSS.n8140 VSS.n8139 0.00054824
R31031 VSS.n8732 VSS.n8731 0.00054824
R31032 VSS.n9324 VSS.n9323 0.00054824
R31033 VSS.n9916 VSS.n9915 0.00054824
R31034 VSS.n10508 VSS.n10507 0.00054824
R31035 VSS.n11100 VSS.n11099 0.00054824
R31036 VSS.n11692 VSS.n11691 0.00054824
R31037 VSS.n12284 VSS.n12283 0.00054824
R31038 VSS.n12876 VSS.n12875 0.00054824
R31039 VSS.n13468 VSS.n13467 0.00054824
R31040 VSS.n14060 VSS.n14059 0.00054824
R31041 VSS.n14652 VSS.n14651 0.00054824
R31042 VSS.n15244 VSS.n15243 0.00054824
R31043 VSS.n15836 VSS.n15835 0.00054824
R31044 VSS.n15838 VSS.n15837 0.00054824
R31045 VSS.n7548 VSS.n7547 0.00054824
R31046 VSS.n18429 VSS.n53 0.00054824
R31047 VSS.n18860 VSS.n18859 0.00054824
R31048 D0_BUF.n15 D0_BUF.n0 400.238
R31049 D0_BUF.n3 D0_BUF.n2 292.5
R31050 D0_BUF.n17 D0_BUF.n16 153.333
R31051 D0_BUF D0_BUF.n17 105.785
R31052 D0_BUF.n0 D0_BUF.t2 83.8685
R31053 D0_BUF.n16 D0_BUF.t5 80.9765
R31054 D0_BUF.n16 D0_BUF.t3 57.8405
R31055 D0_BUF.n0 D0_BUF.t4 54.9485
R31056 D0_BUF.n5 D0_BUF.t1 47.274
R31057 D0_BUF.n2 D0_BUF.t0 27.6955
R31058 D0_BUF.n17 D0_BUF.n15 23.9595
R31059 D0_BUF.n11 D0_BUF.n3 13.177
R31060 D0_BUF.n8 D0_BUF.n3 13.177
R31061 D0_BUF.n11 D0_BUF.n10 9.3005
R31062 D0_BUF.n9 D0_BUF.n8 9.3005
R31063 D0_BUF.n6 D0_BUF.n5 9.3005
R31064 D0_BUF.n7 D0_BUF.n4 9.3005
R31065 D0_BUF.n12 D0_BUF.n1 9.3005
R31066 D0_BUF.n14 D0_BUF.n13 9.3005
R31067 D0_BUF.n13 D0_BUF.n2 9.02061
R31068 D0_BUF.n6 D0_BUF.n2 9.0206
R31069 D0_BUF.n13 D0_BUF.n12 6.02403
R31070 D0_BUF.n7 D0_BUF.n6 6.02403
R31071 D0_BUF.n15 D0_BUF 5.08342
R31072 D0_BUF D0_BUF.n14 2.37139
R31073 D0_BUF.n12 D0_BUF.n11 0.376971
R31074 D0_BUF.n8 D0_BUF.n7 0.376971
R31075 D0_BUF.n10 D0_BUF.n9 0.190717
R31076 D0_BUF.n14 D0_BUF.n1 0.0439783
R31077 D0_BUF.n5 D0_BUF.n4 0.0439783
R31078 D0_BUF.n10 D0_BUF.n1 0.00321739
R31079 D0_BUF.n9 D0_BUF.n4 0.00321739
R31080 VCC.n426 VCC.t184 4282.54
R31081 VCC.n978 VCC.t345 4282.54
R31082 VCC.n1536 VCC.t436 4282.54
R31083 VCC.n2087 VCC.t110 4282.54
R31084 VCC.n2645 VCC.t375 4282.54
R31085 VCC.n3196 VCC.t153 4282.54
R31086 VCC.n3754 VCC.t40 4282.54
R31087 VCC.n4305 VCC.t458 4282.54
R31088 VCC.n4863 VCC.t3 4282.54
R31089 VCC.n5414 VCC.t438 4282.54
R31090 VCC.n5972 VCC.t258 4282.54
R31091 VCC.n6523 VCC.t56 4282.54
R31092 VCC.n7081 VCC.t166 4282.54
R31093 VCC.n7632 VCC.t379 4282.54
R31094 VCC.n8190 VCC.t445 4282.54
R31095 VCC.n8741 VCC.t405 4282.54
R31096 VCC.n9299 VCC.t492 4282.54
R31097 VCC.n9850 VCC.t358 4282.54
R31098 VCC.n10407 VCC.t30 4282.54
R31099 VCC.n10957 VCC.t16 4282.54
R31100 VCC.n11514 VCC.t503 4282.54
R31101 VCC.n12064 VCC.t396 4282.54
R31102 VCC.n12621 VCC.t269 4282.54
R31103 VCC.n13171 VCC.t137 4282.54
R31104 VCC.n13728 VCC.t573 4282.54
R31105 VCC.n14278 VCC.t474 4282.54
R31106 VCC.n14835 VCC.t509 4282.54
R31107 VCC.n15385 VCC.t60 4282.54
R31108 VCC.n15942 VCC.t176 4282.54
R31109 VCC.n16492 VCC.t563 4282.54
R31110 VCC.n17049 VCC.t627 4282.54
R31111 VCC.n17412 VCC.t450 4282.54
R31112 VCC.t191 VCC.t187 1149.1
R31113 VCC.t338 VCC.t342 1149.1
R31114 VCC.t288 VCC.t437 1149.1
R31115 VCC.t430 VCC.t113 1149.1
R31116 VCC.t292 VCC.t374 1149.1
R31117 VCC.t591 VCC.t154 1149.1
R31118 VCC.t576 VCC.t37 1149.1
R31119 VCC.t317 VCC.t457 1149.1
R31120 VCC.t535 VCC.t2 1149.1
R31121 VCC.t326 VCC.t439 1149.1
R31122 VCC.t27 VCC.t255 1149.1
R31123 VCC.t304 VCC.t55 1149.1
R31124 VCC.t227 VCC.t167 1149.1
R31125 VCC.t584 VCC.t378 1149.1
R31126 VCC.t281 VCC.t448 1149.1
R31127 VCC.t35 VCC.t404 1149.1
R31128 VCC.t540 VCC.t493 1149.1
R31129 VCC.t499 VCC.t355 1149.1
R31130 VCC.t239 VCC.t29 1149.1
R31131 VCC.t614 VCC.t13 1149.1
R31132 VCC.t119 VCC.t500 1149.1
R31133 VCC.t217 VCC.t395 1149.1
R31134 VCC.t180 VCC.t266 1149.1
R31135 VCC.t513 VCC.t136 1149.1
R31136 VCC.t604 VCC.t570 1149.1
R31137 VCC.t464 VCC.t471 1149.1
R31138 VCC.t76 VCC.t510 1149.1
R31139 VCC.t556 VCC.t57 1149.1
R31140 VCC.t490 VCC.t173 1149.1
R31141 VCC.t594 VCC.t564 1149.1
R31142 VCC.t124 VCC.t626 1149.1
R31143 VCC.t200 VCC.t449 1149.1
R31144 VCC.t184 VCC.t191 978.443
R31145 VCC.t345 VCC.t338 978.443
R31146 VCC.t436 VCC.t288 978.443
R31147 VCC.t110 VCC.t430 978.443
R31148 VCC.t375 VCC.t292 978.443
R31149 VCC.t153 VCC.t591 978.443
R31150 VCC.t40 VCC.t576 978.443
R31151 VCC.t458 VCC.t317 978.443
R31152 VCC.t3 VCC.t535 978.443
R31153 VCC.t438 VCC.t326 978.443
R31154 VCC.t258 VCC.t27 978.443
R31155 VCC.t56 VCC.t304 978.443
R31156 VCC.t166 VCC.t227 978.443
R31157 VCC.t379 VCC.t584 978.443
R31158 VCC.t445 VCC.t281 978.443
R31159 VCC.t405 VCC.t35 978.443
R31160 VCC.t492 VCC.t540 978.443
R31161 VCC.t358 VCC.t499 978.443
R31162 VCC.t30 VCC.t239 978.443
R31163 VCC.t16 VCC.t614 978.443
R31164 VCC.t503 VCC.t119 978.443
R31165 VCC.t396 VCC.t217 978.443
R31166 VCC.t269 VCC.t180 978.443
R31167 VCC.t137 VCC.t513 978.443
R31168 VCC.t573 VCC.t604 978.443
R31169 VCC.t474 VCC.t464 978.443
R31170 VCC.t509 VCC.t76 978.443
R31171 VCC.t60 VCC.t556 978.443
R31172 VCC.t176 VCC.t490 978.443
R31173 VCC.t563 VCC.t594 978.443
R31174 VCC.t627 VCC.t124 978.443
R31175 VCC.t450 VCC.t200 978.443
R31176 VCC.t187 VCC.t188 972.755
R31177 VCC.t342 VCC.t335 972.755
R31178 VCC.t437 VCC.t285 972.755
R31179 VCC.t113 VCC.t427 972.755
R31180 VCC.t374 VCC.t289 972.755
R31181 VCC.t154 VCC.t588 972.755
R31182 VCC.t37 VCC.t577 972.755
R31183 VCC.t457 VCC.t314 972.755
R31184 VCC.t2 VCC.t536 972.755
R31185 VCC.t439 VCC.t323 972.755
R31186 VCC.t255 VCC.t28 972.755
R31187 VCC.t55 VCC.t305 972.755
R31188 VCC.t167 VCC.t224 972.755
R31189 VCC.t378 VCC.t581 972.755
R31190 VCC.t448 VCC.t278 972.755
R31191 VCC.t404 VCC.t36 972.755
R31192 VCC.t493 VCC.t537 972.755
R31193 VCC.t355 VCC.t496 972.755
R31194 VCC.t29 VCC.t240 972.755
R31195 VCC.t13 VCC.t611 972.755
R31196 VCC.t500 VCC.t120 972.755
R31197 VCC.t395 VCC.t214 972.755
R31198 VCC.t266 VCC.t177 972.755
R31199 VCC.t136 VCC.t514 972.755
R31200 VCC.t570 VCC.t605 972.755
R31201 VCC.t471 VCC.t461 972.755
R31202 VCC.t510 VCC.t73 972.755
R31203 VCC.t57 VCC.t557 972.755
R31204 VCC.t173 VCC.t487 972.755
R31205 VCC.t564 VCC.t595 972.755
R31206 VCC.t626 VCC.t121 972.755
R31207 VCC.t449 VCC.t201 972.755
R31208 VCC.t188 VCC.n425 723.087
R31209 VCC.t335 VCC.n977 723.087
R31210 VCC.t285 VCC.n1535 723.087
R31211 VCC.t427 VCC.n2086 723.087
R31212 VCC.t289 VCC.n2644 723.087
R31213 VCC.t588 VCC.n3195 723.087
R31214 VCC.t577 VCC.n3753 723.087
R31215 VCC.t314 VCC.n4304 723.087
R31216 VCC.t536 VCC.n4862 723.087
R31217 VCC.t323 VCC.n5413 723.087
R31218 VCC.t28 VCC.n5971 723.087
R31219 VCC.t305 VCC.n6522 723.087
R31220 VCC.t224 VCC.n7080 723.087
R31221 VCC.t581 VCC.n7631 723.087
R31222 VCC.t278 VCC.n8189 723.087
R31223 VCC.t36 VCC.n8740 723.087
R31224 VCC.t537 VCC.n9298 723.087
R31225 VCC.t496 VCC.n9849 723.087
R31226 VCC.t240 VCC.n10406 723.087
R31227 VCC.t611 VCC.n10956 723.087
R31228 VCC.t120 VCC.n11513 723.087
R31229 VCC.t214 VCC.n12063 723.087
R31230 VCC.t177 VCC.n12620 723.087
R31231 VCC.t514 VCC.n13170 723.087
R31232 VCC.t605 VCC.n13727 723.087
R31233 VCC.t461 VCC.n14277 723.087
R31234 VCC.t73 VCC.n14834 723.087
R31235 VCC.t557 VCC.n15384 723.087
R31236 VCC.t487 VCC.n15941 723.087
R31237 VCC.t595 VCC.n16491 723.087
R31238 VCC.t121 VCC.n17048 723.087
R31239 VCC.t201 VCC.n17411 723.087
R31240 VCC.t465 VCC.t231 571.485
R31241 VCC.t130 VCC.t569 571.485
R31242 VCC.t470 VCC.t386 571.485
R31243 VCC.t66 VCC.t389 571.485
R31244 VCC.t383 VCC.t298 571.485
R31245 VCC.t431 VCC.t484 571.485
R31246 VCC.t271 VCC.t17 571.485
R31247 VCC.t411 VCC.t555 571.485
R31248 VCC.t181 VCC.t478 571.485
R31249 VCC.t401 VCC.t140 571.485
R31250 VCC.t197 VCC.t598 571.485
R31251 VCC.t523 VCC.t329 571.485
R31252 VCC.t165 VCC.t160 571.485
R31253 VCC.t364 VCC.t6 571.485
R31254 VCC.t259 VCC.t550 571.485
R31255 VCC.t41 VCC.t157 571.485
R31256 VCC.t172 VCC.t442 571.485
R31257 VCC.t620 VCC.t414 571.485
R31258 VCC.t299 VCC.t349 571.485
R31259 VCC.t223 VCC.t103 571.485
R31260 VCC.t243 VCC.t249 571.485
R31261 VCC.t530 VCC.t623 571.485
R31262 VCC.t615 VCC.t334 571.485
R31263 VCC.t394 VCC.t147 571.485
R31264 VCC.t517 VCC.t204 571.485
R31265 VCC.t631 VCC.t234 571.485
R31266 VCC.t274 VCC.t603 571.485
R31267 VCC.t100 VCC.t95 571.485
R31268 VCC.t63 VCC.t127 571.485
R31269 VCC.t107 VCC.t104 571.485
R31270 VCC.t82 VCC.t477 571.485
R31271 VCC.t491 VCC.t85 571.485
R31272 VCC.t89 VCC.t277 571.485
R31273 VCC.t426 VCC.t421 571.485
R31274 VCC.t150 VCC.t320 571.485
R31275 VCC.t69 VCC.t481 571.485
R31276 VCC.t77 VCC.t541 571.485
R31277 VCC.t382 VCC.t49 571.485
R31278 VCC.t94 VCC.t24 571.485
R31279 VCC.t417 VCC.t218 571.485
R31280 VCC.t544 VCC.t451 571.485
R31281 VCC.t194 VCC.t230 571.485
R31282 VCC.t116 VCC.t504 571.485
R31283 VCC.t361 VCC.t86 571.485
R31284 VCC.t72 VCC.t549 571.485
R31285 VCC.t265 VCC.t260 571.485
R31286 VCC.t270 VCC.t562 571.485
R31287 VCC.t293 VCC.t211 571.485
R31288 VCC.t313 VCC.t308 571.485
R31289 VCC.t205 VCC.t630 571.485
R31290 VCC.t252 VCC.t210 571.485
R31291 VCC.t282 VCC.t585 571.485
R31292 VCC.t454 VCC.t133 571.485
R31293 VCC.t524 VCC.t352 571.485
R31294 VCC.t303 VCC.t52 571.485
R31295 VCC.t146 VCC.t339 571.485
R31296 VCC.t244 VCC.t7 571.485
R31297 VCC.t406 VCC.t529 571.485
R31298 VCC.t143 VCC.t418 571.485
R31299 VCC.t44 VCC.t520 571.485
R31300 VCC.t580 VCC.t346 571.485
R31301 VCC.t302 VCC.t610 571.485
R31302 VCC.t12 VCC.t371 571.485
R31303 VCC.n122 VCC.t130 544.823
R31304 VCC.n674 VCC.t66 544.823
R31305 VCC.n1231 VCC.t383 544.823
R31306 VCC.n1783 VCC.t411 544.823
R31307 VCC.n2340 VCC.t181 544.823
R31308 VCC.n2892 VCC.t523 544.823
R31309 VCC.n3449 VCC.t165 544.823
R31310 VCC.n4001 VCC.t41 544.823
R31311 VCC.n4558 VCC.t172 544.823
R31312 VCC.n5110 VCC.t223 544.823
R31313 VCC.n5667 VCC.t243 544.823
R31314 VCC.n6219 VCC.t394 544.823
R31315 VCC.n6776 VCC.t517 544.823
R31316 VCC.n7328 VCC.t100 544.823
R31317 VCC.n7885 VCC.t63 544.823
R31318 VCC.n8437 VCC.t82 544.823
R31319 VCC.n8994 VCC.t89 544.823
R31320 VCC.n9546 VCC.t69 544.823
R31321 VCC.n10102 VCC.t77 544.823
R31322 VCC.n10653 VCC.t417 544.823
R31323 VCC.n11209 VCC.t544 544.823
R31324 VCC.n11760 VCC.t361 544.823
R31325 VCC.n12316 VCC.t72 544.823
R31326 VCC.n12867 VCC.t293 544.823
R31327 VCC.n13423 VCC.t313 544.823
R31328 VCC.n13974 VCC.t282 544.823
R31329 VCC.n14530 VCC.t454 544.823
R31330 VCC.n15081 VCC.t146 544.823
R31331 VCC.n15637 VCC.t244 544.823
R31332 VCC.n16188 VCC.t44 544.823
R31333 VCC.n16744 VCC.t580 544.823
R31334 VCC.n17295 VCC.t12 544.823
R31335 VCC.n209 VCC.t465 542.996
R31336 VCC.n761 VCC.t470 542.996
R31337 VCC.n1319 VCC.t431 542.996
R31338 VCC.n1870 VCC.t271 542.996
R31339 VCC.n2428 VCC.t401 542.996
R31340 VCC.n2979 VCC.t197 542.996
R31341 VCC.n3537 VCC.t364 542.996
R31342 VCC.n4088 VCC.t259 542.996
R31343 VCC.n4646 VCC.t620 542.996
R31344 VCC.n5197 VCC.t299 542.996
R31345 VCC.n5755 VCC.t530 542.996
R31346 VCC.n6306 VCC.t615 542.996
R31347 VCC.n6864 VCC.t631 542.996
R31348 VCC.n7415 VCC.t274 542.996
R31349 VCC.n7973 VCC.t107 542.996
R31350 VCC.n8524 VCC.t491 542.996
R31351 VCC.n9082 VCC.t426 542.996
R31352 VCC.n9633 VCC.t150 542.996
R31353 VCC.n10190 VCC.t382 542.996
R31354 VCC.n10740 VCC.t94 542.996
R31355 VCC.n11297 VCC.t194 542.996
R31356 VCC.n11847 VCC.t116 542.996
R31357 VCC.n12404 VCC.t265 542.996
R31358 VCC.n12954 VCC.t270 542.996
R31359 VCC.n13511 VCC.t205 542.996
R31360 VCC.n14061 VCC.t252 542.996
R31361 VCC.n14618 VCC.t524 542.996
R31362 VCC.n15168 VCC.t303 542.996
R31363 VCC.n15725 VCC.t406 542.996
R31364 VCC.n16275 VCC.t143 542.996
R31365 VCC.n16832 VCC.t302 542.996
R31366 VCC.n209 VCC.n194 187.349
R31367 VCC.n123 VCC.n122 187.349
R31368 VCC.n426 VCC.n79 187.349
R31369 VCC.n761 VCC.n746 187.349
R31370 VCC.n675 VCC.n674 187.349
R31371 VCC.n978 VCC.n631 187.349
R31372 VCC.n1232 VCC.n1231 187.349
R31373 VCC.n1536 VCC.n1188 187.349
R31374 VCC.n1319 VCC.n1304 187.349
R31375 VCC.n1870 VCC.n1855 187.349
R31376 VCC.n1784 VCC.n1783 187.349
R31377 VCC.n2087 VCC.n1740 187.349
R31378 VCC.n2341 VCC.n2340 187.349
R31379 VCC.n2645 VCC.n2297 187.349
R31380 VCC.n2428 VCC.n2413 187.349
R31381 VCC.n2979 VCC.n2964 187.349
R31382 VCC.n2893 VCC.n2892 187.349
R31383 VCC.n3196 VCC.n2849 187.349
R31384 VCC.n3450 VCC.n3449 187.349
R31385 VCC.n3754 VCC.n3406 187.349
R31386 VCC.n3537 VCC.n3522 187.349
R31387 VCC.n4088 VCC.n4073 187.349
R31388 VCC.n4002 VCC.n4001 187.349
R31389 VCC.n4305 VCC.n3958 187.349
R31390 VCC.n4559 VCC.n4558 187.349
R31391 VCC.n4863 VCC.n4515 187.349
R31392 VCC.n4646 VCC.n4631 187.349
R31393 VCC.n5197 VCC.n5182 187.349
R31394 VCC.n5111 VCC.n5110 187.349
R31395 VCC.n5414 VCC.n5067 187.349
R31396 VCC.n5668 VCC.n5667 187.349
R31397 VCC.n5972 VCC.n5624 187.349
R31398 VCC.n5755 VCC.n5740 187.349
R31399 VCC.n6306 VCC.n6291 187.349
R31400 VCC.n6220 VCC.n6219 187.349
R31401 VCC.n6523 VCC.n6176 187.349
R31402 VCC.n6777 VCC.n6776 187.349
R31403 VCC.n7081 VCC.n6733 187.349
R31404 VCC.n6864 VCC.n6849 187.349
R31405 VCC.n7415 VCC.n7400 187.349
R31406 VCC.n7329 VCC.n7328 187.349
R31407 VCC.n7632 VCC.n7285 187.349
R31408 VCC.n7886 VCC.n7885 187.349
R31409 VCC.n8190 VCC.n7842 187.349
R31410 VCC.n7973 VCC.n7958 187.349
R31411 VCC.n8438 VCC.n8437 187.349
R31412 VCC.n8741 VCC.n8394 187.349
R31413 VCC.n8524 VCC.n8509 187.349
R31414 VCC.n8995 VCC.n8994 187.349
R31415 VCC.n9299 VCC.n8951 187.349
R31416 VCC.n9082 VCC.n9067 187.349
R31417 VCC.n9633 VCC.n9618 187.349
R31418 VCC.n9547 VCC.n9546 187.349
R31419 VCC.n9850 VCC.n9503 187.349
R31420 VCC.n10103 VCC.n10102 187.349
R31421 VCC.n10407 VCC.n10059 187.349
R31422 VCC.n10190 VCC.n10175 187.349
R31423 VCC.n10740 VCC.n10725 187.349
R31424 VCC.n10654 VCC.n10653 187.349
R31425 VCC.n10957 VCC.n10610 187.349
R31426 VCC.n11210 VCC.n11209 187.349
R31427 VCC.n11514 VCC.n11166 187.349
R31428 VCC.n11297 VCC.n11282 187.349
R31429 VCC.n11847 VCC.n11832 187.349
R31430 VCC.n11761 VCC.n11760 187.349
R31431 VCC.n12064 VCC.n11717 187.349
R31432 VCC.n12317 VCC.n12316 187.349
R31433 VCC.n12621 VCC.n12273 187.349
R31434 VCC.n12404 VCC.n12389 187.349
R31435 VCC.n12954 VCC.n12939 187.349
R31436 VCC.n12868 VCC.n12867 187.349
R31437 VCC.n13171 VCC.n12824 187.349
R31438 VCC.n13424 VCC.n13423 187.349
R31439 VCC.n13728 VCC.n13380 187.349
R31440 VCC.n13511 VCC.n13496 187.349
R31441 VCC.n14061 VCC.n14046 187.349
R31442 VCC.n13975 VCC.n13974 187.349
R31443 VCC.n14278 VCC.n13931 187.349
R31444 VCC.n14531 VCC.n14530 187.349
R31445 VCC.n14835 VCC.n14487 187.349
R31446 VCC.n14618 VCC.n14603 187.349
R31447 VCC.n15168 VCC.n15153 187.349
R31448 VCC.n15082 VCC.n15081 187.349
R31449 VCC.n15385 VCC.n15038 187.349
R31450 VCC.n15638 VCC.n15637 187.349
R31451 VCC.n15942 VCC.n15594 187.349
R31452 VCC.n15725 VCC.n15710 187.349
R31453 VCC.n16275 VCC.n16260 187.349
R31454 VCC.n16189 VCC.n16188 187.349
R31455 VCC.n16492 VCC.n16145 187.349
R31456 VCC.n16745 VCC.n16744 187.349
R31457 VCC.n17049 VCC.n16701 187.349
R31458 VCC.n16832 VCC.n16817 187.349
R31459 VCC.n17296 VCC.n17295 187.349
R31460 VCC.n17412 VCC.n17252 187.349
R31461 VCC.n231 VCC.n230 185
R31462 VCC.n230 VCC.n229 185
R31463 VCC.n270 VCC.n269 185
R31464 VCC.n269 VCC.n268 185
R31465 VCC.n286 VCC.n140 185
R31466 VCC.n290 VCC.n140 185
R31467 VCC.n292 VCC.n141 185
R31468 VCC.n292 VCC.n291 185
R31469 VCC.n271 VCC.n143 185
R31470 VCC.n143 VCC.n142 185
R31471 VCC.n210 VCC.n208 185
R31472 VCC.n183 VCC.n182 185
R31473 VCC.n182 VCC.n181 185
R31474 VCC.n225 VCC.n224 185
R31475 VCC.n226 VCC.n225 185
R31476 VCC.n180 VCC.n178 185
R31477 VCC.n228 VCC.n180 185
R31478 VCC.n359 VCC.n358 185
R31479 VCC.n360 VCC.n359 185
R31480 VCC.n92 VCC.n91 185
R31481 VCC.n395 VCC.n92 185
R31482 VCC.n416 VCC.n415 185
R31483 VCC.n417 VCC.n416 185
R31484 VCC.n414 VCC.n80 185
R31485 VCC.n418 VCC.n80 185
R31486 VCC.n398 VCC.n397 185
R31487 VCC.n397 VCC.n396 185
R31488 VCC.n427 VCC.n81 185
R31489 VCC.n121 VCC.n120 185
R31490 VCC.n119 VCC.n118 185
R31491 VCC.n336 VCC.n119 185
R31492 VCC.n339 VCC.n338 185
R31493 VCC.n338 VCC.n337 185
R31494 VCC.n107 VCC.n106 185
R31495 VCC.n361 VCC.n107 185
R31496 VCC.n546 VCC.n545 185
R31497 VCC.n547 VCC.n546 185
R31498 VCC.n421 VCC.n56 185
R31499 VCC.n419 VCC.n56 185
R31500 VCC.n493 VCC.n39 185
R31501 VCC.n494 VCC.n493 185
R31502 VCC.n21 VCC.n20 185
R31503 VCC.n526 VCC.n21 185
R31504 VCC.n529 VCC.n528 185
R31505 VCC.n528 VCC.n527 185
R31506 VCC.n24 VCC.n23 185
R31507 VCC.n23 VCC.n22 185
R31508 VCC.n498 VCC.n497 185
R31509 VCC.n497 VCC.n496 185
R31510 VCC.n492 VCC.n491 185
R31511 VCC.n492 VCC.n41 185
R31512 VCC.n475 VCC.n474 185
R31513 VCC.n474 VCC.n473 185
R31514 VCC.n55 VCC.n54 185
R31515 VCC.n471 VCC.n55 185
R31516 VCC.n423 VCC.n422 185
R31517 VCC.n423 VCC.n420 185
R31518 VCC.n4 VCC.n3 185
R31519 VCC.n783 VCC.n782 185
R31520 VCC.n782 VCC.n781 185
R31521 VCC.n822 VCC.n821 185
R31522 VCC.n821 VCC.n820 185
R31523 VCC.n838 VCC.n692 185
R31524 VCC.n842 VCC.n692 185
R31525 VCC.n844 VCC.n693 185
R31526 VCC.n844 VCC.n843 185
R31527 VCC.n823 VCC.n695 185
R31528 VCC.n695 VCC.n694 185
R31529 VCC.n762 VCC.n760 185
R31530 VCC.n735 VCC.n734 185
R31531 VCC.n734 VCC.n733 185
R31532 VCC.n777 VCC.n776 185
R31533 VCC.n778 VCC.n777 185
R31534 VCC.n732 VCC.n730 185
R31535 VCC.n780 VCC.n732 185
R31536 VCC.n911 VCC.n910 185
R31537 VCC.n912 VCC.n911 185
R31538 VCC.n644 VCC.n643 185
R31539 VCC.n947 VCC.n644 185
R31540 VCC.n968 VCC.n967 185
R31541 VCC.n969 VCC.n968 185
R31542 VCC.n966 VCC.n632 185
R31543 VCC.n970 VCC.n632 185
R31544 VCC.n950 VCC.n949 185
R31545 VCC.n949 VCC.n948 185
R31546 VCC.n979 VCC.n633 185
R31547 VCC.n673 VCC.n672 185
R31548 VCC.n671 VCC.n670 185
R31549 VCC.n888 VCC.n671 185
R31550 VCC.n891 VCC.n890 185
R31551 VCC.n890 VCC.n889 185
R31552 VCC.n659 VCC.n658 185
R31553 VCC.n913 VCC.n659 185
R31554 VCC.n973 VCC.n608 185
R31555 VCC.n971 VCC.n608 185
R31556 VCC.n607 VCC.n606 185
R31557 VCC.n1023 VCC.n607 185
R31558 VCC.n1044 VCC.n1043 185
R31559 VCC.n1044 VCC.n593 185
R31560 VCC.n576 VCC.n575 185
R31561 VCC.n575 VCC.n574 185
R31562 VCC.n1081 VCC.n1080 185
R31563 VCC.n1080 VCC.n1079 185
R31564 VCC.n1100 VCC.n1099 185
R31565 VCC.n1101 VCC.n1100 185
R31566 VCC.n1050 VCC.n1049 185
R31567 VCC.n1049 VCC.n1048 185
R31568 VCC.n1027 VCC.n1026 185
R31569 VCC.n1026 VCC.n1025 185
R31570 VCC.n1045 VCC.n591 185
R31571 VCC.n1046 VCC.n1045 185
R31572 VCC.n573 VCC.n572 185
R31573 VCC.n1078 VCC.n573 185
R31574 VCC.n558 VCC.n557 185
R31575 VCC.n975 VCC.n974 185
R31576 VCC.n975 VCC.n972 185
R31577 VCC.n1531 VCC.n1530 185
R31578 VCC.n1530 VCC.n1529 185
R31579 VCC.n1579 VCC.n1578 185
R31580 VCC.n1580 VCC.n1579 185
R31581 VCC.n1162 VCC.n1160 185
R31582 VCC.n1584 VCC.n1162 185
R31583 VCC.n1142 VCC.n1135 185
R31584 VCC.n1620 VCC.n1142 185
R31585 VCC.n1650 VCC.n1649 185
R31586 VCC.n1651 VCC.n1650 185
R31587 VCC.n1654 VCC.n1112 185
R31588 VCC.n1654 VCC.n1653 185
R31589 VCC.n1116 VCC.n1115 185
R31590 VCC.n1115 VCC.n1114 185
R31591 VCC.n1618 VCC.n1617 185
R31592 VCC.n1619 VCC.n1618 185
R31593 VCC.n1582 VCC.n1145 185
R31594 VCC.n1583 VCC.n1582 185
R31595 VCC.n1161 VCC.n1159 185
R31596 VCC.n1581 VCC.n1161 185
R31597 VCC.n1656 VCC.n1655 185
R31598 VCC.n1533 VCC.n1532 185
R31599 VCC.n1533 VCC.n1528 185
R31600 VCC.n1448 VCC.n1447 185
R31601 VCC.n1447 VCC.n1446 185
R31602 VCC.n1216 VCC.n1215 185
R31603 VCC.n1470 VCC.n1216 185
R31604 VCC.n1201 VCC.n1200 185
R31605 VCC.n1504 VCC.n1201 185
R31606 VCC.n1525 VCC.n1524 185
R31607 VCC.n1526 VCC.n1525 185
R31608 VCC.n1523 VCC.n1189 185
R31609 VCC.n1527 VCC.n1189 185
R31610 VCC.n1468 VCC.n1467 185
R31611 VCC.n1469 VCC.n1468 185
R31612 VCC.n1228 VCC.n1227 185
R31613 VCC.n1445 VCC.n1228 185
R31614 VCC.n1507 VCC.n1506 185
R31615 VCC.n1506 VCC.n1505 185
R31616 VCC.n1537 VCC.n1190 185
R31617 VCC.n1230 VCC.n1229 185
R31618 VCC.n1335 VCC.n1334 185
R31619 VCC.n1336 VCC.n1335 185
R31620 VCC.n1290 VCC.n1288 185
R31621 VCC.n1338 VCC.n1290 185
R31622 VCC.n1380 VCC.n1379 185
R31623 VCC.n1379 VCC.n1378 185
R31624 VCC.n1396 VCC.n1250 185
R31625 VCC.n1400 VCC.n1250 185
R31626 VCC.n1402 VCC.n1251 185
R31627 VCC.n1402 VCC.n1401 185
R31628 VCC.n1341 VCC.n1340 185
R31629 VCC.n1340 VCC.n1339 185
R31630 VCC.n1293 VCC.n1292 185
R31631 VCC.n1292 VCC.n1291 185
R31632 VCC.n1381 VCC.n1253 185
R31633 VCC.n1253 VCC.n1252 185
R31634 VCC.n1320 VCC.n1318 185
R31635 VCC.n1892 VCC.n1891 185
R31636 VCC.n1891 VCC.n1890 185
R31637 VCC.n1931 VCC.n1930 185
R31638 VCC.n1930 VCC.n1929 185
R31639 VCC.n1947 VCC.n1801 185
R31640 VCC.n1951 VCC.n1801 185
R31641 VCC.n1953 VCC.n1802 185
R31642 VCC.n1953 VCC.n1952 185
R31643 VCC.n1932 VCC.n1804 185
R31644 VCC.n1804 VCC.n1803 185
R31645 VCC.n1871 VCC.n1869 185
R31646 VCC.n1844 VCC.n1843 185
R31647 VCC.n1843 VCC.n1842 185
R31648 VCC.n1886 VCC.n1885 185
R31649 VCC.n1887 VCC.n1886 185
R31650 VCC.n1841 VCC.n1839 185
R31651 VCC.n1889 VCC.n1841 185
R31652 VCC.n2020 VCC.n2019 185
R31653 VCC.n2021 VCC.n2020 185
R31654 VCC.n1753 VCC.n1752 185
R31655 VCC.n2056 VCC.n1753 185
R31656 VCC.n2077 VCC.n2076 185
R31657 VCC.n2078 VCC.n2077 185
R31658 VCC.n2075 VCC.n1741 185
R31659 VCC.n2079 VCC.n1741 185
R31660 VCC.n2059 VCC.n2058 185
R31661 VCC.n2058 VCC.n2057 185
R31662 VCC.n2088 VCC.n1742 185
R31663 VCC.n1782 VCC.n1781 185
R31664 VCC.n1780 VCC.n1779 185
R31665 VCC.n1997 VCC.n1780 185
R31666 VCC.n2000 VCC.n1999 185
R31667 VCC.n1999 VCC.n1998 185
R31668 VCC.n1768 VCC.n1767 185
R31669 VCC.n2022 VCC.n1768 185
R31670 VCC.n2082 VCC.n1717 185
R31671 VCC.n2080 VCC.n1717 185
R31672 VCC.n1716 VCC.n1715 185
R31673 VCC.n2132 VCC.n1716 185
R31674 VCC.n2153 VCC.n2152 185
R31675 VCC.n2153 VCC.n1702 185
R31676 VCC.n1685 VCC.n1684 185
R31677 VCC.n1684 VCC.n1683 185
R31678 VCC.n2190 VCC.n2189 185
R31679 VCC.n2189 VCC.n2188 185
R31680 VCC.n2209 VCC.n2208 185
R31681 VCC.n2210 VCC.n2209 185
R31682 VCC.n2159 VCC.n2158 185
R31683 VCC.n2158 VCC.n2157 185
R31684 VCC.n2136 VCC.n2135 185
R31685 VCC.n2135 VCC.n2134 185
R31686 VCC.n2154 VCC.n1700 185
R31687 VCC.n2155 VCC.n2154 185
R31688 VCC.n1682 VCC.n1681 185
R31689 VCC.n2187 VCC.n1682 185
R31690 VCC.n1667 VCC.n1666 185
R31691 VCC.n2084 VCC.n2083 185
R31692 VCC.n2084 VCC.n2081 185
R31693 VCC.n2640 VCC.n2639 185
R31694 VCC.n2639 VCC.n2638 185
R31695 VCC.n2688 VCC.n2687 185
R31696 VCC.n2689 VCC.n2688 185
R31697 VCC.n2271 VCC.n2269 185
R31698 VCC.n2693 VCC.n2271 185
R31699 VCC.n2251 VCC.n2244 185
R31700 VCC.n2729 VCC.n2251 185
R31701 VCC.n2759 VCC.n2758 185
R31702 VCC.n2760 VCC.n2759 185
R31703 VCC.n2763 VCC.n2221 185
R31704 VCC.n2763 VCC.n2762 185
R31705 VCC.n2225 VCC.n2224 185
R31706 VCC.n2224 VCC.n2223 185
R31707 VCC.n2727 VCC.n2726 185
R31708 VCC.n2728 VCC.n2727 185
R31709 VCC.n2691 VCC.n2254 185
R31710 VCC.n2692 VCC.n2691 185
R31711 VCC.n2270 VCC.n2268 185
R31712 VCC.n2690 VCC.n2270 185
R31713 VCC.n2765 VCC.n2764 185
R31714 VCC.n2642 VCC.n2641 185
R31715 VCC.n2642 VCC.n2637 185
R31716 VCC.n2557 VCC.n2556 185
R31717 VCC.n2556 VCC.n2555 185
R31718 VCC.n2325 VCC.n2324 185
R31719 VCC.n2579 VCC.n2325 185
R31720 VCC.n2310 VCC.n2309 185
R31721 VCC.n2613 VCC.n2310 185
R31722 VCC.n2634 VCC.n2633 185
R31723 VCC.n2635 VCC.n2634 185
R31724 VCC.n2632 VCC.n2298 185
R31725 VCC.n2636 VCC.n2298 185
R31726 VCC.n2577 VCC.n2576 185
R31727 VCC.n2578 VCC.n2577 185
R31728 VCC.n2337 VCC.n2336 185
R31729 VCC.n2554 VCC.n2337 185
R31730 VCC.n2616 VCC.n2615 185
R31731 VCC.n2615 VCC.n2614 185
R31732 VCC.n2646 VCC.n2299 185
R31733 VCC.n2339 VCC.n2338 185
R31734 VCC.n2444 VCC.n2443 185
R31735 VCC.n2445 VCC.n2444 185
R31736 VCC.n2399 VCC.n2397 185
R31737 VCC.n2447 VCC.n2399 185
R31738 VCC.n2489 VCC.n2488 185
R31739 VCC.n2488 VCC.n2487 185
R31740 VCC.n2505 VCC.n2359 185
R31741 VCC.n2509 VCC.n2359 185
R31742 VCC.n2511 VCC.n2360 185
R31743 VCC.n2511 VCC.n2510 185
R31744 VCC.n2450 VCC.n2449 185
R31745 VCC.n2449 VCC.n2448 185
R31746 VCC.n2402 VCC.n2401 185
R31747 VCC.n2401 VCC.n2400 185
R31748 VCC.n2490 VCC.n2362 185
R31749 VCC.n2362 VCC.n2361 185
R31750 VCC.n2429 VCC.n2427 185
R31751 VCC.n3001 VCC.n3000 185
R31752 VCC.n3000 VCC.n2999 185
R31753 VCC.n3040 VCC.n3039 185
R31754 VCC.n3039 VCC.n3038 185
R31755 VCC.n3056 VCC.n2910 185
R31756 VCC.n3060 VCC.n2910 185
R31757 VCC.n3062 VCC.n2911 185
R31758 VCC.n3062 VCC.n3061 185
R31759 VCC.n3041 VCC.n2913 185
R31760 VCC.n2913 VCC.n2912 185
R31761 VCC.n2980 VCC.n2978 185
R31762 VCC.n2953 VCC.n2952 185
R31763 VCC.n2952 VCC.n2951 185
R31764 VCC.n2995 VCC.n2994 185
R31765 VCC.n2996 VCC.n2995 185
R31766 VCC.n2950 VCC.n2948 185
R31767 VCC.n2998 VCC.n2950 185
R31768 VCC.n3129 VCC.n3128 185
R31769 VCC.n3130 VCC.n3129 185
R31770 VCC.n2862 VCC.n2861 185
R31771 VCC.n3165 VCC.n2862 185
R31772 VCC.n3186 VCC.n3185 185
R31773 VCC.n3187 VCC.n3186 185
R31774 VCC.n3184 VCC.n2850 185
R31775 VCC.n3188 VCC.n2850 185
R31776 VCC.n3168 VCC.n3167 185
R31777 VCC.n3167 VCC.n3166 185
R31778 VCC.n3197 VCC.n2851 185
R31779 VCC.n2891 VCC.n2890 185
R31780 VCC.n2889 VCC.n2888 185
R31781 VCC.n3106 VCC.n2889 185
R31782 VCC.n3109 VCC.n3108 185
R31783 VCC.n3108 VCC.n3107 185
R31784 VCC.n2877 VCC.n2876 185
R31785 VCC.n3131 VCC.n2877 185
R31786 VCC.n3191 VCC.n2826 185
R31787 VCC.n3189 VCC.n2826 185
R31788 VCC.n2825 VCC.n2824 185
R31789 VCC.n3241 VCC.n2825 185
R31790 VCC.n3262 VCC.n3261 185
R31791 VCC.n3262 VCC.n2811 185
R31792 VCC.n2794 VCC.n2793 185
R31793 VCC.n2793 VCC.n2792 185
R31794 VCC.n3299 VCC.n3298 185
R31795 VCC.n3298 VCC.n3297 185
R31796 VCC.n3318 VCC.n3317 185
R31797 VCC.n3319 VCC.n3318 185
R31798 VCC.n3268 VCC.n3267 185
R31799 VCC.n3267 VCC.n3266 185
R31800 VCC.n3245 VCC.n3244 185
R31801 VCC.n3244 VCC.n3243 185
R31802 VCC.n3263 VCC.n2809 185
R31803 VCC.n3264 VCC.n3263 185
R31804 VCC.n2791 VCC.n2790 185
R31805 VCC.n3296 VCC.n2791 185
R31806 VCC.n2776 VCC.n2775 185
R31807 VCC.n3193 VCC.n3192 185
R31808 VCC.n3193 VCC.n3190 185
R31809 VCC.n3749 VCC.n3748 185
R31810 VCC.n3748 VCC.n3747 185
R31811 VCC.n3797 VCC.n3796 185
R31812 VCC.n3798 VCC.n3797 185
R31813 VCC.n3380 VCC.n3378 185
R31814 VCC.n3802 VCC.n3380 185
R31815 VCC.n3360 VCC.n3353 185
R31816 VCC.n3838 VCC.n3360 185
R31817 VCC.n3868 VCC.n3867 185
R31818 VCC.n3869 VCC.n3868 185
R31819 VCC.n3872 VCC.n3330 185
R31820 VCC.n3872 VCC.n3871 185
R31821 VCC.n3334 VCC.n3333 185
R31822 VCC.n3333 VCC.n3332 185
R31823 VCC.n3836 VCC.n3835 185
R31824 VCC.n3837 VCC.n3836 185
R31825 VCC.n3800 VCC.n3363 185
R31826 VCC.n3801 VCC.n3800 185
R31827 VCC.n3379 VCC.n3377 185
R31828 VCC.n3799 VCC.n3379 185
R31829 VCC.n3874 VCC.n3873 185
R31830 VCC.n3751 VCC.n3750 185
R31831 VCC.n3751 VCC.n3746 185
R31832 VCC.n3666 VCC.n3665 185
R31833 VCC.n3665 VCC.n3664 185
R31834 VCC.n3434 VCC.n3433 185
R31835 VCC.n3688 VCC.n3434 185
R31836 VCC.n3419 VCC.n3418 185
R31837 VCC.n3722 VCC.n3419 185
R31838 VCC.n3743 VCC.n3742 185
R31839 VCC.n3744 VCC.n3743 185
R31840 VCC.n3741 VCC.n3407 185
R31841 VCC.n3745 VCC.n3407 185
R31842 VCC.n3686 VCC.n3685 185
R31843 VCC.n3687 VCC.n3686 185
R31844 VCC.n3446 VCC.n3445 185
R31845 VCC.n3663 VCC.n3446 185
R31846 VCC.n3725 VCC.n3724 185
R31847 VCC.n3724 VCC.n3723 185
R31848 VCC.n3755 VCC.n3408 185
R31849 VCC.n3448 VCC.n3447 185
R31850 VCC.n3553 VCC.n3552 185
R31851 VCC.n3554 VCC.n3553 185
R31852 VCC.n3508 VCC.n3506 185
R31853 VCC.n3556 VCC.n3508 185
R31854 VCC.n3598 VCC.n3597 185
R31855 VCC.n3597 VCC.n3596 185
R31856 VCC.n3614 VCC.n3468 185
R31857 VCC.n3618 VCC.n3468 185
R31858 VCC.n3620 VCC.n3469 185
R31859 VCC.n3620 VCC.n3619 185
R31860 VCC.n3559 VCC.n3558 185
R31861 VCC.n3558 VCC.n3557 185
R31862 VCC.n3511 VCC.n3510 185
R31863 VCC.n3510 VCC.n3509 185
R31864 VCC.n3599 VCC.n3471 185
R31865 VCC.n3471 VCC.n3470 185
R31866 VCC.n3538 VCC.n3536 185
R31867 VCC.n4110 VCC.n4109 185
R31868 VCC.n4109 VCC.n4108 185
R31869 VCC.n4149 VCC.n4148 185
R31870 VCC.n4148 VCC.n4147 185
R31871 VCC.n4165 VCC.n4019 185
R31872 VCC.n4169 VCC.n4019 185
R31873 VCC.n4171 VCC.n4020 185
R31874 VCC.n4171 VCC.n4170 185
R31875 VCC.n4150 VCC.n4022 185
R31876 VCC.n4022 VCC.n4021 185
R31877 VCC.n4089 VCC.n4087 185
R31878 VCC.n4062 VCC.n4061 185
R31879 VCC.n4061 VCC.n4060 185
R31880 VCC.n4104 VCC.n4103 185
R31881 VCC.n4105 VCC.n4104 185
R31882 VCC.n4059 VCC.n4057 185
R31883 VCC.n4107 VCC.n4059 185
R31884 VCC.n4238 VCC.n4237 185
R31885 VCC.n4239 VCC.n4238 185
R31886 VCC.n3971 VCC.n3970 185
R31887 VCC.n4274 VCC.n3971 185
R31888 VCC.n4295 VCC.n4294 185
R31889 VCC.n4296 VCC.n4295 185
R31890 VCC.n4293 VCC.n3959 185
R31891 VCC.n4297 VCC.n3959 185
R31892 VCC.n4277 VCC.n4276 185
R31893 VCC.n4276 VCC.n4275 185
R31894 VCC.n4306 VCC.n3960 185
R31895 VCC.n4000 VCC.n3999 185
R31896 VCC.n3998 VCC.n3997 185
R31897 VCC.n4215 VCC.n3998 185
R31898 VCC.n4218 VCC.n4217 185
R31899 VCC.n4217 VCC.n4216 185
R31900 VCC.n3986 VCC.n3985 185
R31901 VCC.n4240 VCC.n3986 185
R31902 VCC.n4300 VCC.n3935 185
R31903 VCC.n4298 VCC.n3935 185
R31904 VCC.n3934 VCC.n3933 185
R31905 VCC.n4350 VCC.n3934 185
R31906 VCC.n4371 VCC.n4370 185
R31907 VCC.n4371 VCC.n3920 185
R31908 VCC.n3903 VCC.n3902 185
R31909 VCC.n3902 VCC.n3901 185
R31910 VCC.n4408 VCC.n4407 185
R31911 VCC.n4407 VCC.n4406 185
R31912 VCC.n4427 VCC.n4426 185
R31913 VCC.n4428 VCC.n4427 185
R31914 VCC.n4377 VCC.n4376 185
R31915 VCC.n4376 VCC.n4375 185
R31916 VCC.n4354 VCC.n4353 185
R31917 VCC.n4353 VCC.n4352 185
R31918 VCC.n4372 VCC.n3918 185
R31919 VCC.n4373 VCC.n4372 185
R31920 VCC.n3900 VCC.n3899 185
R31921 VCC.n4405 VCC.n3900 185
R31922 VCC.n3885 VCC.n3884 185
R31923 VCC.n4302 VCC.n4301 185
R31924 VCC.n4302 VCC.n4299 185
R31925 VCC.n4858 VCC.n4857 185
R31926 VCC.n4857 VCC.n4856 185
R31927 VCC.n4906 VCC.n4905 185
R31928 VCC.n4907 VCC.n4906 185
R31929 VCC.n4489 VCC.n4487 185
R31930 VCC.n4911 VCC.n4489 185
R31931 VCC.n4469 VCC.n4462 185
R31932 VCC.n4947 VCC.n4469 185
R31933 VCC.n4977 VCC.n4976 185
R31934 VCC.n4978 VCC.n4977 185
R31935 VCC.n4981 VCC.n4439 185
R31936 VCC.n4981 VCC.n4980 185
R31937 VCC.n4443 VCC.n4442 185
R31938 VCC.n4442 VCC.n4441 185
R31939 VCC.n4945 VCC.n4944 185
R31940 VCC.n4946 VCC.n4945 185
R31941 VCC.n4909 VCC.n4472 185
R31942 VCC.n4910 VCC.n4909 185
R31943 VCC.n4488 VCC.n4486 185
R31944 VCC.n4908 VCC.n4488 185
R31945 VCC.n4983 VCC.n4982 185
R31946 VCC.n4860 VCC.n4859 185
R31947 VCC.n4860 VCC.n4855 185
R31948 VCC.n4775 VCC.n4774 185
R31949 VCC.n4774 VCC.n4773 185
R31950 VCC.n4543 VCC.n4542 185
R31951 VCC.n4797 VCC.n4543 185
R31952 VCC.n4528 VCC.n4527 185
R31953 VCC.n4831 VCC.n4528 185
R31954 VCC.n4852 VCC.n4851 185
R31955 VCC.n4853 VCC.n4852 185
R31956 VCC.n4850 VCC.n4516 185
R31957 VCC.n4854 VCC.n4516 185
R31958 VCC.n4795 VCC.n4794 185
R31959 VCC.n4796 VCC.n4795 185
R31960 VCC.n4555 VCC.n4554 185
R31961 VCC.n4772 VCC.n4555 185
R31962 VCC.n4834 VCC.n4833 185
R31963 VCC.n4833 VCC.n4832 185
R31964 VCC.n4864 VCC.n4517 185
R31965 VCC.n4557 VCC.n4556 185
R31966 VCC.n4662 VCC.n4661 185
R31967 VCC.n4663 VCC.n4662 185
R31968 VCC.n4617 VCC.n4615 185
R31969 VCC.n4665 VCC.n4617 185
R31970 VCC.n4707 VCC.n4706 185
R31971 VCC.n4706 VCC.n4705 185
R31972 VCC.n4723 VCC.n4577 185
R31973 VCC.n4727 VCC.n4577 185
R31974 VCC.n4729 VCC.n4578 185
R31975 VCC.n4729 VCC.n4728 185
R31976 VCC.n4668 VCC.n4667 185
R31977 VCC.n4667 VCC.n4666 185
R31978 VCC.n4620 VCC.n4619 185
R31979 VCC.n4619 VCC.n4618 185
R31980 VCC.n4708 VCC.n4580 185
R31981 VCC.n4580 VCC.n4579 185
R31982 VCC.n4647 VCC.n4645 185
R31983 VCC.n5219 VCC.n5218 185
R31984 VCC.n5218 VCC.n5217 185
R31985 VCC.n5258 VCC.n5257 185
R31986 VCC.n5257 VCC.n5256 185
R31987 VCC.n5274 VCC.n5128 185
R31988 VCC.n5278 VCC.n5128 185
R31989 VCC.n5280 VCC.n5129 185
R31990 VCC.n5280 VCC.n5279 185
R31991 VCC.n5259 VCC.n5131 185
R31992 VCC.n5131 VCC.n5130 185
R31993 VCC.n5198 VCC.n5196 185
R31994 VCC.n5171 VCC.n5170 185
R31995 VCC.n5170 VCC.n5169 185
R31996 VCC.n5213 VCC.n5212 185
R31997 VCC.n5214 VCC.n5213 185
R31998 VCC.n5168 VCC.n5166 185
R31999 VCC.n5216 VCC.n5168 185
R32000 VCC.n5347 VCC.n5346 185
R32001 VCC.n5348 VCC.n5347 185
R32002 VCC.n5080 VCC.n5079 185
R32003 VCC.n5383 VCC.n5080 185
R32004 VCC.n5404 VCC.n5403 185
R32005 VCC.n5405 VCC.n5404 185
R32006 VCC.n5402 VCC.n5068 185
R32007 VCC.n5406 VCC.n5068 185
R32008 VCC.n5386 VCC.n5385 185
R32009 VCC.n5385 VCC.n5384 185
R32010 VCC.n5415 VCC.n5069 185
R32011 VCC.n5109 VCC.n5108 185
R32012 VCC.n5107 VCC.n5106 185
R32013 VCC.n5324 VCC.n5107 185
R32014 VCC.n5327 VCC.n5326 185
R32015 VCC.n5326 VCC.n5325 185
R32016 VCC.n5095 VCC.n5094 185
R32017 VCC.n5349 VCC.n5095 185
R32018 VCC.n5409 VCC.n5044 185
R32019 VCC.n5407 VCC.n5044 185
R32020 VCC.n5043 VCC.n5042 185
R32021 VCC.n5459 VCC.n5043 185
R32022 VCC.n5480 VCC.n5479 185
R32023 VCC.n5480 VCC.n5029 185
R32024 VCC.n5012 VCC.n5011 185
R32025 VCC.n5011 VCC.n5010 185
R32026 VCC.n5517 VCC.n5516 185
R32027 VCC.n5516 VCC.n5515 185
R32028 VCC.n5536 VCC.n5535 185
R32029 VCC.n5537 VCC.n5536 185
R32030 VCC.n5486 VCC.n5485 185
R32031 VCC.n5485 VCC.n5484 185
R32032 VCC.n5463 VCC.n5462 185
R32033 VCC.n5462 VCC.n5461 185
R32034 VCC.n5481 VCC.n5027 185
R32035 VCC.n5482 VCC.n5481 185
R32036 VCC.n5009 VCC.n5008 185
R32037 VCC.n5514 VCC.n5009 185
R32038 VCC.n4994 VCC.n4993 185
R32039 VCC.n5411 VCC.n5410 185
R32040 VCC.n5411 VCC.n5408 185
R32041 VCC.n5967 VCC.n5966 185
R32042 VCC.n5966 VCC.n5965 185
R32043 VCC.n6015 VCC.n6014 185
R32044 VCC.n6016 VCC.n6015 185
R32045 VCC.n5598 VCC.n5596 185
R32046 VCC.n6020 VCC.n5598 185
R32047 VCC.n5578 VCC.n5571 185
R32048 VCC.n6056 VCC.n5578 185
R32049 VCC.n6086 VCC.n6085 185
R32050 VCC.n6087 VCC.n6086 185
R32051 VCC.n6090 VCC.n5548 185
R32052 VCC.n6090 VCC.n6089 185
R32053 VCC.n5552 VCC.n5551 185
R32054 VCC.n5551 VCC.n5550 185
R32055 VCC.n6054 VCC.n6053 185
R32056 VCC.n6055 VCC.n6054 185
R32057 VCC.n6018 VCC.n5581 185
R32058 VCC.n6019 VCC.n6018 185
R32059 VCC.n5597 VCC.n5595 185
R32060 VCC.n6017 VCC.n5597 185
R32061 VCC.n6092 VCC.n6091 185
R32062 VCC.n5969 VCC.n5968 185
R32063 VCC.n5969 VCC.n5964 185
R32064 VCC.n5884 VCC.n5883 185
R32065 VCC.n5883 VCC.n5882 185
R32066 VCC.n5652 VCC.n5651 185
R32067 VCC.n5906 VCC.n5652 185
R32068 VCC.n5637 VCC.n5636 185
R32069 VCC.n5940 VCC.n5637 185
R32070 VCC.n5961 VCC.n5960 185
R32071 VCC.n5962 VCC.n5961 185
R32072 VCC.n5959 VCC.n5625 185
R32073 VCC.n5963 VCC.n5625 185
R32074 VCC.n5904 VCC.n5903 185
R32075 VCC.n5905 VCC.n5904 185
R32076 VCC.n5664 VCC.n5663 185
R32077 VCC.n5881 VCC.n5664 185
R32078 VCC.n5943 VCC.n5942 185
R32079 VCC.n5942 VCC.n5941 185
R32080 VCC.n5973 VCC.n5626 185
R32081 VCC.n5666 VCC.n5665 185
R32082 VCC.n5771 VCC.n5770 185
R32083 VCC.n5772 VCC.n5771 185
R32084 VCC.n5726 VCC.n5724 185
R32085 VCC.n5774 VCC.n5726 185
R32086 VCC.n5816 VCC.n5815 185
R32087 VCC.n5815 VCC.n5814 185
R32088 VCC.n5832 VCC.n5686 185
R32089 VCC.n5836 VCC.n5686 185
R32090 VCC.n5838 VCC.n5687 185
R32091 VCC.n5838 VCC.n5837 185
R32092 VCC.n5777 VCC.n5776 185
R32093 VCC.n5776 VCC.n5775 185
R32094 VCC.n5729 VCC.n5728 185
R32095 VCC.n5728 VCC.n5727 185
R32096 VCC.n5817 VCC.n5689 185
R32097 VCC.n5689 VCC.n5688 185
R32098 VCC.n5756 VCC.n5754 185
R32099 VCC.n6328 VCC.n6327 185
R32100 VCC.n6327 VCC.n6326 185
R32101 VCC.n6367 VCC.n6366 185
R32102 VCC.n6366 VCC.n6365 185
R32103 VCC.n6383 VCC.n6237 185
R32104 VCC.n6387 VCC.n6237 185
R32105 VCC.n6389 VCC.n6238 185
R32106 VCC.n6389 VCC.n6388 185
R32107 VCC.n6368 VCC.n6240 185
R32108 VCC.n6240 VCC.n6239 185
R32109 VCC.n6307 VCC.n6305 185
R32110 VCC.n6280 VCC.n6279 185
R32111 VCC.n6279 VCC.n6278 185
R32112 VCC.n6322 VCC.n6321 185
R32113 VCC.n6323 VCC.n6322 185
R32114 VCC.n6277 VCC.n6275 185
R32115 VCC.n6325 VCC.n6277 185
R32116 VCC.n6456 VCC.n6455 185
R32117 VCC.n6457 VCC.n6456 185
R32118 VCC.n6189 VCC.n6188 185
R32119 VCC.n6492 VCC.n6189 185
R32120 VCC.n6513 VCC.n6512 185
R32121 VCC.n6514 VCC.n6513 185
R32122 VCC.n6511 VCC.n6177 185
R32123 VCC.n6515 VCC.n6177 185
R32124 VCC.n6495 VCC.n6494 185
R32125 VCC.n6494 VCC.n6493 185
R32126 VCC.n6524 VCC.n6178 185
R32127 VCC.n6218 VCC.n6217 185
R32128 VCC.n6216 VCC.n6215 185
R32129 VCC.n6433 VCC.n6216 185
R32130 VCC.n6436 VCC.n6435 185
R32131 VCC.n6435 VCC.n6434 185
R32132 VCC.n6204 VCC.n6203 185
R32133 VCC.n6458 VCC.n6204 185
R32134 VCC.n6518 VCC.n6153 185
R32135 VCC.n6516 VCC.n6153 185
R32136 VCC.n6152 VCC.n6151 185
R32137 VCC.n6568 VCC.n6152 185
R32138 VCC.n6589 VCC.n6588 185
R32139 VCC.n6589 VCC.n6138 185
R32140 VCC.n6121 VCC.n6120 185
R32141 VCC.n6120 VCC.n6119 185
R32142 VCC.n6626 VCC.n6625 185
R32143 VCC.n6625 VCC.n6624 185
R32144 VCC.n6645 VCC.n6644 185
R32145 VCC.n6646 VCC.n6645 185
R32146 VCC.n6595 VCC.n6594 185
R32147 VCC.n6594 VCC.n6593 185
R32148 VCC.n6572 VCC.n6571 185
R32149 VCC.n6571 VCC.n6570 185
R32150 VCC.n6590 VCC.n6136 185
R32151 VCC.n6591 VCC.n6590 185
R32152 VCC.n6118 VCC.n6117 185
R32153 VCC.n6623 VCC.n6118 185
R32154 VCC.n6103 VCC.n6102 185
R32155 VCC.n6520 VCC.n6519 185
R32156 VCC.n6520 VCC.n6517 185
R32157 VCC.n7076 VCC.n7075 185
R32158 VCC.n7075 VCC.n7074 185
R32159 VCC.n7124 VCC.n7123 185
R32160 VCC.n7125 VCC.n7124 185
R32161 VCC.n6707 VCC.n6705 185
R32162 VCC.n7129 VCC.n6707 185
R32163 VCC.n6687 VCC.n6680 185
R32164 VCC.n7165 VCC.n6687 185
R32165 VCC.n7195 VCC.n7194 185
R32166 VCC.n7196 VCC.n7195 185
R32167 VCC.n7199 VCC.n6657 185
R32168 VCC.n7199 VCC.n7198 185
R32169 VCC.n6661 VCC.n6660 185
R32170 VCC.n6660 VCC.n6659 185
R32171 VCC.n7163 VCC.n7162 185
R32172 VCC.n7164 VCC.n7163 185
R32173 VCC.n7127 VCC.n6690 185
R32174 VCC.n7128 VCC.n7127 185
R32175 VCC.n6706 VCC.n6704 185
R32176 VCC.n7126 VCC.n6706 185
R32177 VCC.n7201 VCC.n7200 185
R32178 VCC.n7078 VCC.n7077 185
R32179 VCC.n7078 VCC.n7073 185
R32180 VCC.n6993 VCC.n6992 185
R32181 VCC.n6992 VCC.n6991 185
R32182 VCC.n6761 VCC.n6760 185
R32183 VCC.n7015 VCC.n6761 185
R32184 VCC.n6746 VCC.n6745 185
R32185 VCC.n7049 VCC.n6746 185
R32186 VCC.n7070 VCC.n7069 185
R32187 VCC.n7071 VCC.n7070 185
R32188 VCC.n7068 VCC.n6734 185
R32189 VCC.n7072 VCC.n6734 185
R32190 VCC.n7013 VCC.n7012 185
R32191 VCC.n7014 VCC.n7013 185
R32192 VCC.n6773 VCC.n6772 185
R32193 VCC.n6990 VCC.n6773 185
R32194 VCC.n7052 VCC.n7051 185
R32195 VCC.n7051 VCC.n7050 185
R32196 VCC.n7082 VCC.n6735 185
R32197 VCC.n6775 VCC.n6774 185
R32198 VCC.n6880 VCC.n6879 185
R32199 VCC.n6881 VCC.n6880 185
R32200 VCC.n6835 VCC.n6833 185
R32201 VCC.n6883 VCC.n6835 185
R32202 VCC.n6925 VCC.n6924 185
R32203 VCC.n6924 VCC.n6923 185
R32204 VCC.n6941 VCC.n6795 185
R32205 VCC.n6945 VCC.n6795 185
R32206 VCC.n6947 VCC.n6796 185
R32207 VCC.n6947 VCC.n6946 185
R32208 VCC.n6886 VCC.n6885 185
R32209 VCC.n6885 VCC.n6884 185
R32210 VCC.n6838 VCC.n6837 185
R32211 VCC.n6837 VCC.n6836 185
R32212 VCC.n6926 VCC.n6798 185
R32213 VCC.n6798 VCC.n6797 185
R32214 VCC.n6865 VCC.n6863 185
R32215 VCC.n7437 VCC.n7436 185
R32216 VCC.n7436 VCC.n7435 185
R32217 VCC.n7476 VCC.n7475 185
R32218 VCC.n7475 VCC.n7474 185
R32219 VCC.n7492 VCC.n7346 185
R32220 VCC.n7496 VCC.n7346 185
R32221 VCC.n7498 VCC.n7347 185
R32222 VCC.n7498 VCC.n7497 185
R32223 VCC.n7477 VCC.n7349 185
R32224 VCC.n7349 VCC.n7348 185
R32225 VCC.n7416 VCC.n7414 185
R32226 VCC.n7389 VCC.n7388 185
R32227 VCC.n7388 VCC.n7387 185
R32228 VCC.n7431 VCC.n7430 185
R32229 VCC.n7432 VCC.n7431 185
R32230 VCC.n7386 VCC.n7384 185
R32231 VCC.n7434 VCC.n7386 185
R32232 VCC.n7565 VCC.n7564 185
R32233 VCC.n7566 VCC.n7565 185
R32234 VCC.n7298 VCC.n7297 185
R32235 VCC.n7601 VCC.n7298 185
R32236 VCC.n7622 VCC.n7621 185
R32237 VCC.n7623 VCC.n7622 185
R32238 VCC.n7620 VCC.n7286 185
R32239 VCC.n7624 VCC.n7286 185
R32240 VCC.n7604 VCC.n7603 185
R32241 VCC.n7603 VCC.n7602 185
R32242 VCC.n7633 VCC.n7287 185
R32243 VCC.n7327 VCC.n7326 185
R32244 VCC.n7325 VCC.n7324 185
R32245 VCC.n7542 VCC.n7325 185
R32246 VCC.n7545 VCC.n7544 185
R32247 VCC.n7544 VCC.n7543 185
R32248 VCC.n7313 VCC.n7312 185
R32249 VCC.n7567 VCC.n7313 185
R32250 VCC.n7627 VCC.n7262 185
R32251 VCC.n7625 VCC.n7262 185
R32252 VCC.n7261 VCC.n7260 185
R32253 VCC.n7677 VCC.n7261 185
R32254 VCC.n7698 VCC.n7697 185
R32255 VCC.n7698 VCC.n7247 185
R32256 VCC.n7230 VCC.n7229 185
R32257 VCC.n7229 VCC.n7228 185
R32258 VCC.n7735 VCC.n7734 185
R32259 VCC.n7734 VCC.n7733 185
R32260 VCC.n7754 VCC.n7753 185
R32261 VCC.n7755 VCC.n7754 185
R32262 VCC.n7704 VCC.n7703 185
R32263 VCC.n7703 VCC.n7702 185
R32264 VCC.n7681 VCC.n7680 185
R32265 VCC.n7680 VCC.n7679 185
R32266 VCC.n7699 VCC.n7245 185
R32267 VCC.n7700 VCC.n7699 185
R32268 VCC.n7227 VCC.n7226 185
R32269 VCC.n7732 VCC.n7227 185
R32270 VCC.n7212 VCC.n7211 185
R32271 VCC.n7629 VCC.n7628 185
R32272 VCC.n7629 VCC.n7626 185
R32273 VCC.n8185 VCC.n8184 185
R32274 VCC.n8184 VCC.n8183 185
R32275 VCC.n8233 VCC.n8232 185
R32276 VCC.n8234 VCC.n8233 185
R32277 VCC.n7816 VCC.n7814 185
R32278 VCC.n8238 VCC.n7816 185
R32279 VCC.n7796 VCC.n7789 185
R32280 VCC.n8274 VCC.n7796 185
R32281 VCC.n8304 VCC.n8303 185
R32282 VCC.n8305 VCC.n8304 185
R32283 VCC.n8308 VCC.n7766 185
R32284 VCC.n8308 VCC.n8307 185
R32285 VCC.n7770 VCC.n7769 185
R32286 VCC.n7769 VCC.n7768 185
R32287 VCC.n8272 VCC.n8271 185
R32288 VCC.n8273 VCC.n8272 185
R32289 VCC.n8236 VCC.n7799 185
R32290 VCC.n8237 VCC.n8236 185
R32291 VCC.n7815 VCC.n7813 185
R32292 VCC.n8235 VCC.n7815 185
R32293 VCC.n8310 VCC.n8309 185
R32294 VCC.n8187 VCC.n8186 185
R32295 VCC.n8187 VCC.n8182 185
R32296 VCC.n8102 VCC.n8101 185
R32297 VCC.n8101 VCC.n8100 185
R32298 VCC.n7870 VCC.n7869 185
R32299 VCC.n8124 VCC.n7870 185
R32300 VCC.n7855 VCC.n7854 185
R32301 VCC.n8158 VCC.n7855 185
R32302 VCC.n8179 VCC.n8178 185
R32303 VCC.n8180 VCC.n8179 185
R32304 VCC.n8177 VCC.n7843 185
R32305 VCC.n8181 VCC.n7843 185
R32306 VCC.n8122 VCC.n8121 185
R32307 VCC.n8123 VCC.n8122 185
R32308 VCC.n7882 VCC.n7881 185
R32309 VCC.n8099 VCC.n7882 185
R32310 VCC.n8161 VCC.n8160 185
R32311 VCC.n8160 VCC.n8159 185
R32312 VCC.n8191 VCC.n7844 185
R32313 VCC.n7884 VCC.n7883 185
R32314 VCC.n7989 VCC.n7988 185
R32315 VCC.n7990 VCC.n7989 185
R32316 VCC.n7944 VCC.n7942 185
R32317 VCC.n7992 VCC.n7944 185
R32318 VCC.n8034 VCC.n8033 185
R32319 VCC.n8033 VCC.n8032 185
R32320 VCC.n8050 VCC.n7904 185
R32321 VCC.n8054 VCC.n7904 185
R32322 VCC.n8056 VCC.n7905 185
R32323 VCC.n8056 VCC.n8055 185
R32324 VCC.n7995 VCC.n7994 185
R32325 VCC.n7994 VCC.n7993 185
R32326 VCC.n7947 VCC.n7946 185
R32327 VCC.n7946 VCC.n7945 185
R32328 VCC.n8035 VCC.n7907 185
R32329 VCC.n7907 VCC.n7906 185
R32330 VCC.n7974 VCC.n7972 185
R32331 VCC.n8674 VCC.n8673 185
R32332 VCC.n8675 VCC.n8674 185
R32333 VCC.n8407 VCC.n8406 185
R32334 VCC.n8710 VCC.n8407 185
R32335 VCC.n8731 VCC.n8730 185
R32336 VCC.n8732 VCC.n8731 185
R32337 VCC.n8729 VCC.n8395 185
R32338 VCC.n8733 VCC.n8395 185
R32339 VCC.n8713 VCC.n8712 185
R32340 VCC.n8712 VCC.n8711 185
R32341 VCC.n8742 VCC.n8396 185
R32342 VCC.n8436 VCC.n8435 185
R32343 VCC.n8434 VCC.n8433 185
R32344 VCC.n8651 VCC.n8434 185
R32345 VCC.n8654 VCC.n8653 185
R32346 VCC.n8653 VCC.n8652 185
R32347 VCC.n8422 VCC.n8421 185
R32348 VCC.n8676 VCC.n8422 185
R32349 VCC.n8736 VCC.n8371 185
R32350 VCC.n8734 VCC.n8371 185
R32351 VCC.n8370 VCC.n8369 185
R32352 VCC.n8786 VCC.n8370 185
R32353 VCC.n8807 VCC.n8806 185
R32354 VCC.n8807 VCC.n8356 185
R32355 VCC.n8339 VCC.n8338 185
R32356 VCC.n8338 VCC.n8337 185
R32357 VCC.n8844 VCC.n8843 185
R32358 VCC.n8843 VCC.n8842 185
R32359 VCC.n8863 VCC.n8862 185
R32360 VCC.n8864 VCC.n8863 185
R32361 VCC.n8813 VCC.n8812 185
R32362 VCC.n8812 VCC.n8811 185
R32363 VCC.n8790 VCC.n8789 185
R32364 VCC.n8789 VCC.n8788 185
R32365 VCC.n8808 VCC.n8354 185
R32366 VCC.n8809 VCC.n8808 185
R32367 VCC.n8336 VCC.n8335 185
R32368 VCC.n8841 VCC.n8336 185
R32369 VCC.n8321 VCC.n8320 185
R32370 VCC.n8738 VCC.n8737 185
R32371 VCC.n8738 VCC.n8735 185
R32372 VCC.n8540 VCC.n8539 185
R32373 VCC.n8541 VCC.n8540 185
R32374 VCC.n8495 VCC.n8493 185
R32375 VCC.n8543 VCC.n8495 185
R32376 VCC.n8585 VCC.n8584 185
R32377 VCC.n8584 VCC.n8583 185
R32378 VCC.n8601 VCC.n8455 185
R32379 VCC.n8605 VCC.n8455 185
R32380 VCC.n8607 VCC.n8456 185
R32381 VCC.n8607 VCC.n8606 185
R32382 VCC.n8546 VCC.n8545 185
R32383 VCC.n8545 VCC.n8544 185
R32384 VCC.n8498 VCC.n8497 185
R32385 VCC.n8497 VCC.n8496 185
R32386 VCC.n8586 VCC.n8458 185
R32387 VCC.n8458 VCC.n8457 185
R32388 VCC.n8525 VCC.n8523 185
R32389 VCC.n9294 VCC.n9293 185
R32390 VCC.n9293 VCC.n9292 185
R32391 VCC.n9342 VCC.n9341 185
R32392 VCC.n9343 VCC.n9342 185
R32393 VCC.n8925 VCC.n8923 185
R32394 VCC.n9347 VCC.n8925 185
R32395 VCC.n8905 VCC.n8898 185
R32396 VCC.n9383 VCC.n8905 185
R32397 VCC.n9413 VCC.n9412 185
R32398 VCC.n9414 VCC.n9413 185
R32399 VCC.n9417 VCC.n8875 185
R32400 VCC.n9417 VCC.n9416 185
R32401 VCC.n8879 VCC.n8878 185
R32402 VCC.n8878 VCC.n8877 185
R32403 VCC.n9381 VCC.n9380 185
R32404 VCC.n9382 VCC.n9381 185
R32405 VCC.n9345 VCC.n8908 185
R32406 VCC.n9346 VCC.n9345 185
R32407 VCC.n8924 VCC.n8922 185
R32408 VCC.n9344 VCC.n8924 185
R32409 VCC.n9419 VCC.n9418 185
R32410 VCC.n9296 VCC.n9295 185
R32411 VCC.n9296 VCC.n9291 185
R32412 VCC.n9211 VCC.n9210 185
R32413 VCC.n9210 VCC.n9209 185
R32414 VCC.n8979 VCC.n8978 185
R32415 VCC.n9233 VCC.n8979 185
R32416 VCC.n8964 VCC.n8963 185
R32417 VCC.n9267 VCC.n8964 185
R32418 VCC.n9288 VCC.n9287 185
R32419 VCC.n9289 VCC.n9288 185
R32420 VCC.n9286 VCC.n8952 185
R32421 VCC.n9290 VCC.n8952 185
R32422 VCC.n9231 VCC.n9230 185
R32423 VCC.n9232 VCC.n9231 185
R32424 VCC.n8991 VCC.n8990 185
R32425 VCC.n9208 VCC.n8991 185
R32426 VCC.n9270 VCC.n9269 185
R32427 VCC.n9269 VCC.n9268 185
R32428 VCC.n9300 VCC.n8953 185
R32429 VCC.n8993 VCC.n8992 185
R32430 VCC.n9098 VCC.n9097 185
R32431 VCC.n9099 VCC.n9098 185
R32432 VCC.n9053 VCC.n9051 185
R32433 VCC.n9101 VCC.n9053 185
R32434 VCC.n9143 VCC.n9142 185
R32435 VCC.n9142 VCC.n9141 185
R32436 VCC.n9159 VCC.n9013 185
R32437 VCC.n9163 VCC.n9013 185
R32438 VCC.n9165 VCC.n9014 185
R32439 VCC.n9165 VCC.n9164 185
R32440 VCC.n9104 VCC.n9103 185
R32441 VCC.n9103 VCC.n9102 185
R32442 VCC.n9056 VCC.n9055 185
R32443 VCC.n9055 VCC.n9054 185
R32444 VCC.n9144 VCC.n9016 185
R32445 VCC.n9016 VCC.n9015 185
R32446 VCC.n9083 VCC.n9081 185
R32447 VCC.n9655 VCC.n9654 185
R32448 VCC.n9654 VCC.n9653 185
R32449 VCC.n9694 VCC.n9693 185
R32450 VCC.n9693 VCC.n9692 185
R32451 VCC.n9710 VCC.n9564 185
R32452 VCC.n9714 VCC.n9564 185
R32453 VCC.n9716 VCC.n9565 185
R32454 VCC.n9716 VCC.n9715 185
R32455 VCC.n9695 VCC.n9567 185
R32456 VCC.n9567 VCC.n9566 185
R32457 VCC.n9634 VCC.n9632 185
R32458 VCC.n9607 VCC.n9606 185
R32459 VCC.n9606 VCC.n9605 185
R32460 VCC.n9649 VCC.n9648 185
R32461 VCC.n9650 VCC.n9649 185
R32462 VCC.n9604 VCC.n9602 185
R32463 VCC.n9652 VCC.n9604 185
R32464 VCC.n9783 VCC.n9782 185
R32465 VCC.n9784 VCC.n9783 185
R32466 VCC.n9516 VCC.n9515 185
R32467 VCC.n9819 VCC.n9516 185
R32468 VCC.n9840 VCC.n9839 185
R32469 VCC.n9841 VCC.n9840 185
R32470 VCC.n9838 VCC.n9504 185
R32471 VCC.n9842 VCC.n9504 185
R32472 VCC.n9822 VCC.n9821 185
R32473 VCC.n9821 VCC.n9820 185
R32474 VCC.n9851 VCC.n9505 185
R32475 VCC.n9545 VCC.n9544 185
R32476 VCC.n9543 VCC.n9542 185
R32477 VCC.n9760 VCC.n9543 185
R32478 VCC.n9763 VCC.n9762 185
R32479 VCC.n9762 VCC.n9761 185
R32480 VCC.n9531 VCC.n9530 185
R32481 VCC.n9785 VCC.n9531 185
R32482 VCC.n9845 VCC.n9480 185
R32483 VCC.n9843 VCC.n9480 185
R32484 VCC.n9479 VCC.n9478 185
R32485 VCC.n9895 VCC.n9479 185
R32486 VCC.n9916 VCC.n9915 185
R32487 VCC.n9916 VCC.n9465 185
R32488 VCC.n9448 VCC.n9447 185
R32489 VCC.n9447 VCC.n9446 185
R32490 VCC.n9953 VCC.n9952 185
R32491 VCC.n9952 VCC.n9951 185
R32492 VCC.n9972 VCC.n9971 185
R32493 VCC.n9973 VCC.n9972 185
R32494 VCC.n9922 VCC.n9921 185
R32495 VCC.n9921 VCC.n9920 185
R32496 VCC.n9899 VCC.n9898 185
R32497 VCC.n9898 VCC.n9897 185
R32498 VCC.n9917 VCC.n9463 185
R32499 VCC.n9918 VCC.n9917 185
R32500 VCC.n9445 VCC.n9444 185
R32501 VCC.n9950 VCC.n9445 185
R32502 VCC.n9430 VCC.n9429 185
R32503 VCC.n9847 VCC.n9846 185
R32504 VCC.n9847 VCC.n9844 185
R32505 VCC.n10402 VCC.n10401 185
R32506 VCC.n10401 VCC.n10400 185
R32507 VCC.n10450 VCC.n10449 185
R32508 VCC.n10451 VCC.n10450 185
R32509 VCC.n10033 VCC.n10031 185
R32510 VCC.n10455 VCC.n10033 185
R32511 VCC.n10013 VCC.n10006 185
R32512 VCC.n10491 VCC.n10013 185
R32513 VCC.n10521 VCC.n10520 185
R32514 VCC.n10522 VCC.n10521 185
R32515 VCC.n10525 VCC.n9983 185
R32516 VCC.n10525 VCC.n10524 185
R32517 VCC.n9987 VCC.n9986 185
R32518 VCC.n9986 VCC.n9985 185
R32519 VCC.n10489 VCC.n10488 185
R32520 VCC.n10490 VCC.n10489 185
R32521 VCC.n10453 VCC.n10016 185
R32522 VCC.n10454 VCC.n10453 185
R32523 VCC.n10032 VCC.n10030 185
R32524 VCC.n10452 VCC.n10032 185
R32525 VCC.n10527 VCC.n10526 185
R32526 VCC.n10404 VCC.n10403 185
R32527 VCC.n10404 VCC.n10399 185
R32528 VCC.n10319 VCC.n10318 185
R32529 VCC.n10318 VCC.n10317 185
R32530 VCC.n10087 VCC.n10086 185
R32531 VCC.n10341 VCC.n10087 185
R32532 VCC.n10072 VCC.n10071 185
R32533 VCC.n10375 VCC.n10072 185
R32534 VCC.n10396 VCC.n10395 185
R32535 VCC.n10397 VCC.n10396 185
R32536 VCC.n10394 VCC.n10060 185
R32537 VCC.n10398 VCC.n10060 185
R32538 VCC.n10339 VCC.n10338 185
R32539 VCC.n10340 VCC.n10339 185
R32540 VCC.n10099 VCC.n10098 185
R32541 VCC.n10316 VCC.n10099 185
R32542 VCC.n10378 VCC.n10377 185
R32543 VCC.n10377 VCC.n10376 185
R32544 VCC.n10408 VCC.n10061 185
R32545 VCC.n10101 VCC.n10100 185
R32546 VCC.n10206 VCC.n10205 185
R32547 VCC.n10207 VCC.n10206 185
R32548 VCC.n10161 VCC.n10159 185
R32549 VCC.n10209 VCC.n10161 185
R32550 VCC.n10251 VCC.n10250 185
R32551 VCC.n10250 VCC.n10249 185
R32552 VCC.n10267 VCC.n10121 185
R32553 VCC.n10271 VCC.n10121 185
R32554 VCC.n10273 VCC.n10122 185
R32555 VCC.n10273 VCC.n10272 185
R32556 VCC.n10212 VCC.n10211 185
R32557 VCC.n10211 VCC.n10210 185
R32558 VCC.n10164 VCC.n10163 185
R32559 VCC.n10163 VCC.n10162 185
R32560 VCC.n10252 VCC.n10124 185
R32561 VCC.n10124 VCC.n10123 185
R32562 VCC.n10191 VCC.n10189 185
R32563 VCC.n10762 VCC.n10761 185
R32564 VCC.n10761 VCC.n10760 185
R32565 VCC.n10801 VCC.n10800 185
R32566 VCC.n10800 VCC.n10799 185
R32567 VCC.n10817 VCC.n10671 185
R32568 VCC.n10821 VCC.n10671 185
R32569 VCC.n10823 VCC.n10672 185
R32570 VCC.n10823 VCC.n10822 185
R32571 VCC.n10802 VCC.n10674 185
R32572 VCC.n10674 VCC.n10673 185
R32573 VCC.n10741 VCC.n10739 185
R32574 VCC.n10714 VCC.n10713 185
R32575 VCC.n10713 VCC.n10712 185
R32576 VCC.n10756 VCC.n10755 185
R32577 VCC.n10757 VCC.n10756 185
R32578 VCC.n10711 VCC.n10709 185
R32579 VCC.n10759 VCC.n10711 185
R32580 VCC.n10890 VCC.n10889 185
R32581 VCC.n10891 VCC.n10890 185
R32582 VCC.n10623 VCC.n10622 185
R32583 VCC.n10926 VCC.n10623 185
R32584 VCC.n10947 VCC.n10946 185
R32585 VCC.n10948 VCC.n10947 185
R32586 VCC.n10945 VCC.n10611 185
R32587 VCC.n10949 VCC.n10611 185
R32588 VCC.n10929 VCC.n10928 185
R32589 VCC.n10928 VCC.n10927 185
R32590 VCC.n10958 VCC.n10612 185
R32591 VCC.n10652 VCC.n10651 185
R32592 VCC.n10650 VCC.n10649 185
R32593 VCC.n10867 VCC.n10650 185
R32594 VCC.n10870 VCC.n10869 185
R32595 VCC.n10869 VCC.n10868 185
R32596 VCC.n10638 VCC.n10637 185
R32597 VCC.n10892 VCC.n10638 185
R32598 VCC.n10952 VCC.n10587 185
R32599 VCC.n10950 VCC.n10587 185
R32600 VCC.n10586 VCC.n10585 185
R32601 VCC.n11002 VCC.n10586 185
R32602 VCC.n11023 VCC.n11022 185
R32603 VCC.n11023 VCC.n10572 185
R32604 VCC.n10555 VCC.n10554 185
R32605 VCC.n10554 VCC.n10553 185
R32606 VCC.n11060 VCC.n11059 185
R32607 VCC.n11059 VCC.n11058 185
R32608 VCC.n11079 VCC.n11078 185
R32609 VCC.n11080 VCC.n11079 185
R32610 VCC.n11029 VCC.n11028 185
R32611 VCC.n11028 VCC.n11027 185
R32612 VCC.n11006 VCC.n11005 185
R32613 VCC.n11005 VCC.n11004 185
R32614 VCC.n11024 VCC.n10570 185
R32615 VCC.n11025 VCC.n11024 185
R32616 VCC.n10552 VCC.n10551 185
R32617 VCC.n11057 VCC.n10552 185
R32618 VCC.n10537 VCC.n10536 185
R32619 VCC.n10954 VCC.n10953 185
R32620 VCC.n10954 VCC.n10951 185
R32621 VCC.n11509 VCC.n11508 185
R32622 VCC.n11508 VCC.n11507 185
R32623 VCC.n11557 VCC.n11556 185
R32624 VCC.n11558 VCC.n11557 185
R32625 VCC.n11140 VCC.n11138 185
R32626 VCC.n11562 VCC.n11140 185
R32627 VCC.n11120 VCC.n11113 185
R32628 VCC.n11598 VCC.n11120 185
R32629 VCC.n11628 VCC.n11627 185
R32630 VCC.n11629 VCC.n11628 185
R32631 VCC.n11632 VCC.n11090 185
R32632 VCC.n11632 VCC.n11631 185
R32633 VCC.n11094 VCC.n11093 185
R32634 VCC.n11093 VCC.n11092 185
R32635 VCC.n11596 VCC.n11595 185
R32636 VCC.n11597 VCC.n11596 185
R32637 VCC.n11560 VCC.n11123 185
R32638 VCC.n11561 VCC.n11560 185
R32639 VCC.n11139 VCC.n11137 185
R32640 VCC.n11559 VCC.n11139 185
R32641 VCC.n11634 VCC.n11633 185
R32642 VCC.n11511 VCC.n11510 185
R32643 VCC.n11511 VCC.n11506 185
R32644 VCC.n11426 VCC.n11425 185
R32645 VCC.n11425 VCC.n11424 185
R32646 VCC.n11194 VCC.n11193 185
R32647 VCC.n11448 VCC.n11194 185
R32648 VCC.n11179 VCC.n11178 185
R32649 VCC.n11482 VCC.n11179 185
R32650 VCC.n11503 VCC.n11502 185
R32651 VCC.n11504 VCC.n11503 185
R32652 VCC.n11501 VCC.n11167 185
R32653 VCC.n11505 VCC.n11167 185
R32654 VCC.n11446 VCC.n11445 185
R32655 VCC.n11447 VCC.n11446 185
R32656 VCC.n11206 VCC.n11205 185
R32657 VCC.n11423 VCC.n11206 185
R32658 VCC.n11485 VCC.n11484 185
R32659 VCC.n11484 VCC.n11483 185
R32660 VCC.n11515 VCC.n11168 185
R32661 VCC.n11208 VCC.n11207 185
R32662 VCC.n11313 VCC.n11312 185
R32663 VCC.n11314 VCC.n11313 185
R32664 VCC.n11268 VCC.n11266 185
R32665 VCC.n11316 VCC.n11268 185
R32666 VCC.n11358 VCC.n11357 185
R32667 VCC.n11357 VCC.n11356 185
R32668 VCC.n11374 VCC.n11228 185
R32669 VCC.n11378 VCC.n11228 185
R32670 VCC.n11380 VCC.n11229 185
R32671 VCC.n11380 VCC.n11379 185
R32672 VCC.n11319 VCC.n11318 185
R32673 VCC.n11318 VCC.n11317 185
R32674 VCC.n11271 VCC.n11270 185
R32675 VCC.n11270 VCC.n11269 185
R32676 VCC.n11359 VCC.n11231 185
R32677 VCC.n11231 VCC.n11230 185
R32678 VCC.n11298 VCC.n11296 185
R32679 VCC.n11869 VCC.n11868 185
R32680 VCC.n11868 VCC.n11867 185
R32681 VCC.n11908 VCC.n11907 185
R32682 VCC.n11907 VCC.n11906 185
R32683 VCC.n11924 VCC.n11778 185
R32684 VCC.n11928 VCC.n11778 185
R32685 VCC.n11930 VCC.n11779 185
R32686 VCC.n11930 VCC.n11929 185
R32687 VCC.n11909 VCC.n11781 185
R32688 VCC.n11781 VCC.n11780 185
R32689 VCC.n11848 VCC.n11846 185
R32690 VCC.n11821 VCC.n11820 185
R32691 VCC.n11820 VCC.n11819 185
R32692 VCC.n11863 VCC.n11862 185
R32693 VCC.n11864 VCC.n11863 185
R32694 VCC.n11818 VCC.n11816 185
R32695 VCC.n11866 VCC.n11818 185
R32696 VCC.n11997 VCC.n11996 185
R32697 VCC.n11998 VCC.n11997 185
R32698 VCC.n11730 VCC.n11729 185
R32699 VCC.n12033 VCC.n11730 185
R32700 VCC.n12054 VCC.n12053 185
R32701 VCC.n12055 VCC.n12054 185
R32702 VCC.n12052 VCC.n11718 185
R32703 VCC.n12056 VCC.n11718 185
R32704 VCC.n12036 VCC.n12035 185
R32705 VCC.n12035 VCC.n12034 185
R32706 VCC.n12065 VCC.n11719 185
R32707 VCC.n11759 VCC.n11758 185
R32708 VCC.n11757 VCC.n11756 185
R32709 VCC.n11974 VCC.n11757 185
R32710 VCC.n11977 VCC.n11976 185
R32711 VCC.n11976 VCC.n11975 185
R32712 VCC.n11745 VCC.n11744 185
R32713 VCC.n11999 VCC.n11745 185
R32714 VCC.n12059 VCC.n11694 185
R32715 VCC.n12057 VCC.n11694 185
R32716 VCC.n11693 VCC.n11692 185
R32717 VCC.n12109 VCC.n11693 185
R32718 VCC.n12130 VCC.n12129 185
R32719 VCC.n12130 VCC.n11679 185
R32720 VCC.n11662 VCC.n11661 185
R32721 VCC.n11661 VCC.n11660 185
R32722 VCC.n12167 VCC.n12166 185
R32723 VCC.n12166 VCC.n12165 185
R32724 VCC.n12186 VCC.n12185 185
R32725 VCC.n12187 VCC.n12186 185
R32726 VCC.n12136 VCC.n12135 185
R32727 VCC.n12135 VCC.n12134 185
R32728 VCC.n12113 VCC.n12112 185
R32729 VCC.n12112 VCC.n12111 185
R32730 VCC.n12131 VCC.n11677 185
R32731 VCC.n12132 VCC.n12131 185
R32732 VCC.n11659 VCC.n11658 185
R32733 VCC.n12164 VCC.n11659 185
R32734 VCC.n11644 VCC.n11643 185
R32735 VCC.n12061 VCC.n12060 185
R32736 VCC.n12061 VCC.n12058 185
R32737 VCC.n12616 VCC.n12615 185
R32738 VCC.n12615 VCC.n12614 185
R32739 VCC.n12664 VCC.n12663 185
R32740 VCC.n12665 VCC.n12664 185
R32741 VCC.n12247 VCC.n12245 185
R32742 VCC.n12669 VCC.n12247 185
R32743 VCC.n12227 VCC.n12220 185
R32744 VCC.n12705 VCC.n12227 185
R32745 VCC.n12735 VCC.n12734 185
R32746 VCC.n12736 VCC.n12735 185
R32747 VCC.n12739 VCC.n12197 185
R32748 VCC.n12739 VCC.n12738 185
R32749 VCC.n12201 VCC.n12200 185
R32750 VCC.n12200 VCC.n12199 185
R32751 VCC.n12703 VCC.n12702 185
R32752 VCC.n12704 VCC.n12703 185
R32753 VCC.n12667 VCC.n12230 185
R32754 VCC.n12668 VCC.n12667 185
R32755 VCC.n12246 VCC.n12244 185
R32756 VCC.n12666 VCC.n12246 185
R32757 VCC.n12741 VCC.n12740 185
R32758 VCC.n12618 VCC.n12617 185
R32759 VCC.n12618 VCC.n12613 185
R32760 VCC.n12533 VCC.n12532 185
R32761 VCC.n12532 VCC.n12531 185
R32762 VCC.n12301 VCC.n12300 185
R32763 VCC.n12555 VCC.n12301 185
R32764 VCC.n12286 VCC.n12285 185
R32765 VCC.n12589 VCC.n12286 185
R32766 VCC.n12610 VCC.n12609 185
R32767 VCC.n12611 VCC.n12610 185
R32768 VCC.n12608 VCC.n12274 185
R32769 VCC.n12612 VCC.n12274 185
R32770 VCC.n12553 VCC.n12552 185
R32771 VCC.n12554 VCC.n12553 185
R32772 VCC.n12313 VCC.n12312 185
R32773 VCC.n12530 VCC.n12313 185
R32774 VCC.n12592 VCC.n12591 185
R32775 VCC.n12591 VCC.n12590 185
R32776 VCC.n12622 VCC.n12275 185
R32777 VCC.n12315 VCC.n12314 185
R32778 VCC.n12420 VCC.n12419 185
R32779 VCC.n12421 VCC.n12420 185
R32780 VCC.n12375 VCC.n12373 185
R32781 VCC.n12423 VCC.n12375 185
R32782 VCC.n12465 VCC.n12464 185
R32783 VCC.n12464 VCC.n12463 185
R32784 VCC.n12481 VCC.n12335 185
R32785 VCC.n12485 VCC.n12335 185
R32786 VCC.n12487 VCC.n12336 185
R32787 VCC.n12487 VCC.n12486 185
R32788 VCC.n12426 VCC.n12425 185
R32789 VCC.n12425 VCC.n12424 185
R32790 VCC.n12378 VCC.n12377 185
R32791 VCC.n12377 VCC.n12376 185
R32792 VCC.n12466 VCC.n12338 185
R32793 VCC.n12338 VCC.n12337 185
R32794 VCC.n12405 VCC.n12403 185
R32795 VCC.n12976 VCC.n12975 185
R32796 VCC.n12975 VCC.n12974 185
R32797 VCC.n13015 VCC.n13014 185
R32798 VCC.n13014 VCC.n13013 185
R32799 VCC.n13031 VCC.n12885 185
R32800 VCC.n13035 VCC.n12885 185
R32801 VCC.n13037 VCC.n12886 185
R32802 VCC.n13037 VCC.n13036 185
R32803 VCC.n13016 VCC.n12888 185
R32804 VCC.n12888 VCC.n12887 185
R32805 VCC.n12955 VCC.n12953 185
R32806 VCC.n12928 VCC.n12927 185
R32807 VCC.n12927 VCC.n12926 185
R32808 VCC.n12970 VCC.n12969 185
R32809 VCC.n12971 VCC.n12970 185
R32810 VCC.n12925 VCC.n12923 185
R32811 VCC.n12973 VCC.n12925 185
R32812 VCC.n13104 VCC.n13103 185
R32813 VCC.n13105 VCC.n13104 185
R32814 VCC.n12837 VCC.n12836 185
R32815 VCC.n13140 VCC.n12837 185
R32816 VCC.n13161 VCC.n13160 185
R32817 VCC.n13162 VCC.n13161 185
R32818 VCC.n13159 VCC.n12825 185
R32819 VCC.n13163 VCC.n12825 185
R32820 VCC.n13143 VCC.n13142 185
R32821 VCC.n13142 VCC.n13141 185
R32822 VCC.n13172 VCC.n12826 185
R32823 VCC.n12866 VCC.n12865 185
R32824 VCC.n12864 VCC.n12863 185
R32825 VCC.n13081 VCC.n12864 185
R32826 VCC.n13084 VCC.n13083 185
R32827 VCC.n13083 VCC.n13082 185
R32828 VCC.n12852 VCC.n12851 185
R32829 VCC.n13106 VCC.n12852 185
R32830 VCC.n13166 VCC.n12801 185
R32831 VCC.n13164 VCC.n12801 185
R32832 VCC.n12800 VCC.n12799 185
R32833 VCC.n13216 VCC.n12800 185
R32834 VCC.n13237 VCC.n13236 185
R32835 VCC.n13237 VCC.n12786 185
R32836 VCC.n12769 VCC.n12768 185
R32837 VCC.n12768 VCC.n12767 185
R32838 VCC.n13274 VCC.n13273 185
R32839 VCC.n13273 VCC.n13272 185
R32840 VCC.n13293 VCC.n13292 185
R32841 VCC.n13294 VCC.n13293 185
R32842 VCC.n13243 VCC.n13242 185
R32843 VCC.n13242 VCC.n13241 185
R32844 VCC.n13220 VCC.n13219 185
R32845 VCC.n13219 VCC.n13218 185
R32846 VCC.n13238 VCC.n12784 185
R32847 VCC.n13239 VCC.n13238 185
R32848 VCC.n12766 VCC.n12765 185
R32849 VCC.n13271 VCC.n12766 185
R32850 VCC.n12751 VCC.n12750 185
R32851 VCC.n13168 VCC.n13167 185
R32852 VCC.n13168 VCC.n13165 185
R32853 VCC.n13723 VCC.n13722 185
R32854 VCC.n13722 VCC.n13721 185
R32855 VCC.n13771 VCC.n13770 185
R32856 VCC.n13772 VCC.n13771 185
R32857 VCC.n13354 VCC.n13352 185
R32858 VCC.n13776 VCC.n13354 185
R32859 VCC.n13334 VCC.n13327 185
R32860 VCC.n13812 VCC.n13334 185
R32861 VCC.n13842 VCC.n13841 185
R32862 VCC.n13843 VCC.n13842 185
R32863 VCC.n13846 VCC.n13304 185
R32864 VCC.n13846 VCC.n13845 185
R32865 VCC.n13308 VCC.n13307 185
R32866 VCC.n13307 VCC.n13306 185
R32867 VCC.n13810 VCC.n13809 185
R32868 VCC.n13811 VCC.n13810 185
R32869 VCC.n13774 VCC.n13337 185
R32870 VCC.n13775 VCC.n13774 185
R32871 VCC.n13353 VCC.n13351 185
R32872 VCC.n13773 VCC.n13353 185
R32873 VCC.n13848 VCC.n13847 185
R32874 VCC.n13725 VCC.n13724 185
R32875 VCC.n13725 VCC.n13720 185
R32876 VCC.n13640 VCC.n13639 185
R32877 VCC.n13639 VCC.n13638 185
R32878 VCC.n13408 VCC.n13407 185
R32879 VCC.n13662 VCC.n13408 185
R32880 VCC.n13393 VCC.n13392 185
R32881 VCC.n13696 VCC.n13393 185
R32882 VCC.n13717 VCC.n13716 185
R32883 VCC.n13718 VCC.n13717 185
R32884 VCC.n13715 VCC.n13381 185
R32885 VCC.n13719 VCC.n13381 185
R32886 VCC.n13660 VCC.n13659 185
R32887 VCC.n13661 VCC.n13660 185
R32888 VCC.n13420 VCC.n13419 185
R32889 VCC.n13637 VCC.n13420 185
R32890 VCC.n13699 VCC.n13698 185
R32891 VCC.n13698 VCC.n13697 185
R32892 VCC.n13729 VCC.n13382 185
R32893 VCC.n13422 VCC.n13421 185
R32894 VCC.n13527 VCC.n13526 185
R32895 VCC.n13528 VCC.n13527 185
R32896 VCC.n13482 VCC.n13480 185
R32897 VCC.n13530 VCC.n13482 185
R32898 VCC.n13572 VCC.n13571 185
R32899 VCC.n13571 VCC.n13570 185
R32900 VCC.n13588 VCC.n13442 185
R32901 VCC.n13592 VCC.n13442 185
R32902 VCC.n13594 VCC.n13443 185
R32903 VCC.n13594 VCC.n13593 185
R32904 VCC.n13533 VCC.n13532 185
R32905 VCC.n13532 VCC.n13531 185
R32906 VCC.n13485 VCC.n13484 185
R32907 VCC.n13484 VCC.n13483 185
R32908 VCC.n13573 VCC.n13445 185
R32909 VCC.n13445 VCC.n13444 185
R32910 VCC.n13512 VCC.n13510 185
R32911 VCC.n14083 VCC.n14082 185
R32912 VCC.n14082 VCC.n14081 185
R32913 VCC.n14122 VCC.n14121 185
R32914 VCC.n14121 VCC.n14120 185
R32915 VCC.n14138 VCC.n13992 185
R32916 VCC.n14142 VCC.n13992 185
R32917 VCC.n14144 VCC.n13993 185
R32918 VCC.n14144 VCC.n14143 185
R32919 VCC.n14123 VCC.n13995 185
R32920 VCC.n13995 VCC.n13994 185
R32921 VCC.n14062 VCC.n14060 185
R32922 VCC.n14035 VCC.n14034 185
R32923 VCC.n14034 VCC.n14033 185
R32924 VCC.n14077 VCC.n14076 185
R32925 VCC.n14078 VCC.n14077 185
R32926 VCC.n14032 VCC.n14030 185
R32927 VCC.n14080 VCC.n14032 185
R32928 VCC.n14211 VCC.n14210 185
R32929 VCC.n14212 VCC.n14211 185
R32930 VCC.n13944 VCC.n13943 185
R32931 VCC.n14247 VCC.n13944 185
R32932 VCC.n14268 VCC.n14267 185
R32933 VCC.n14269 VCC.n14268 185
R32934 VCC.n14266 VCC.n13932 185
R32935 VCC.n14270 VCC.n13932 185
R32936 VCC.n14250 VCC.n14249 185
R32937 VCC.n14249 VCC.n14248 185
R32938 VCC.n14279 VCC.n13933 185
R32939 VCC.n13973 VCC.n13972 185
R32940 VCC.n13971 VCC.n13970 185
R32941 VCC.n14188 VCC.n13971 185
R32942 VCC.n14191 VCC.n14190 185
R32943 VCC.n14190 VCC.n14189 185
R32944 VCC.n13959 VCC.n13958 185
R32945 VCC.n14213 VCC.n13959 185
R32946 VCC.n14273 VCC.n13908 185
R32947 VCC.n14271 VCC.n13908 185
R32948 VCC.n13907 VCC.n13906 185
R32949 VCC.n14323 VCC.n13907 185
R32950 VCC.n14344 VCC.n14343 185
R32951 VCC.n14344 VCC.n13893 185
R32952 VCC.n13876 VCC.n13875 185
R32953 VCC.n13875 VCC.n13874 185
R32954 VCC.n14381 VCC.n14380 185
R32955 VCC.n14380 VCC.n14379 185
R32956 VCC.n14400 VCC.n14399 185
R32957 VCC.n14401 VCC.n14400 185
R32958 VCC.n14350 VCC.n14349 185
R32959 VCC.n14349 VCC.n14348 185
R32960 VCC.n14327 VCC.n14326 185
R32961 VCC.n14326 VCC.n14325 185
R32962 VCC.n14345 VCC.n13891 185
R32963 VCC.n14346 VCC.n14345 185
R32964 VCC.n13873 VCC.n13872 185
R32965 VCC.n14378 VCC.n13873 185
R32966 VCC.n13858 VCC.n13857 185
R32967 VCC.n14275 VCC.n14274 185
R32968 VCC.n14275 VCC.n14272 185
R32969 VCC.n14830 VCC.n14829 185
R32970 VCC.n14829 VCC.n14828 185
R32971 VCC.n14878 VCC.n14877 185
R32972 VCC.n14879 VCC.n14878 185
R32973 VCC.n14461 VCC.n14459 185
R32974 VCC.n14883 VCC.n14461 185
R32975 VCC.n14441 VCC.n14434 185
R32976 VCC.n14919 VCC.n14441 185
R32977 VCC.n14949 VCC.n14948 185
R32978 VCC.n14950 VCC.n14949 185
R32979 VCC.n14953 VCC.n14411 185
R32980 VCC.n14953 VCC.n14952 185
R32981 VCC.n14415 VCC.n14414 185
R32982 VCC.n14414 VCC.n14413 185
R32983 VCC.n14917 VCC.n14916 185
R32984 VCC.n14918 VCC.n14917 185
R32985 VCC.n14881 VCC.n14444 185
R32986 VCC.n14882 VCC.n14881 185
R32987 VCC.n14460 VCC.n14458 185
R32988 VCC.n14880 VCC.n14460 185
R32989 VCC.n14955 VCC.n14954 185
R32990 VCC.n14832 VCC.n14831 185
R32991 VCC.n14832 VCC.n14827 185
R32992 VCC.n14747 VCC.n14746 185
R32993 VCC.n14746 VCC.n14745 185
R32994 VCC.n14515 VCC.n14514 185
R32995 VCC.n14769 VCC.n14515 185
R32996 VCC.n14500 VCC.n14499 185
R32997 VCC.n14803 VCC.n14500 185
R32998 VCC.n14824 VCC.n14823 185
R32999 VCC.n14825 VCC.n14824 185
R33000 VCC.n14822 VCC.n14488 185
R33001 VCC.n14826 VCC.n14488 185
R33002 VCC.n14767 VCC.n14766 185
R33003 VCC.n14768 VCC.n14767 185
R33004 VCC.n14527 VCC.n14526 185
R33005 VCC.n14744 VCC.n14527 185
R33006 VCC.n14806 VCC.n14805 185
R33007 VCC.n14805 VCC.n14804 185
R33008 VCC.n14836 VCC.n14489 185
R33009 VCC.n14529 VCC.n14528 185
R33010 VCC.n14634 VCC.n14633 185
R33011 VCC.n14635 VCC.n14634 185
R33012 VCC.n14589 VCC.n14587 185
R33013 VCC.n14637 VCC.n14589 185
R33014 VCC.n14679 VCC.n14678 185
R33015 VCC.n14678 VCC.n14677 185
R33016 VCC.n14695 VCC.n14549 185
R33017 VCC.n14699 VCC.n14549 185
R33018 VCC.n14701 VCC.n14550 185
R33019 VCC.n14701 VCC.n14700 185
R33020 VCC.n14640 VCC.n14639 185
R33021 VCC.n14639 VCC.n14638 185
R33022 VCC.n14592 VCC.n14591 185
R33023 VCC.n14591 VCC.n14590 185
R33024 VCC.n14680 VCC.n14552 185
R33025 VCC.n14552 VCC.n14551 185
R33026 VCC.n14619 VCC.n14617 185
R33027 VCC.n15190 VCC.n15189 185
R33028 VCC.n15189 VCC.n15188 185
R33029 VCC.n15229 VCC.n15228 185
R33030 VCC.n15228 VCC.n15227 185
R33031 VCC.n15245 VCC.n15099 185
R33032 VCC.n15249 VCC.n15099 185
R33033 VCC.n15251 VCC.n15100 185
R33034 VCC.n15251 VCC.n15250 185
R33035 VCC.n15230 VCC.n15102 185
R33036 VCC.n15102 VCC.n15101 185
R33037 VCC.n15169 VCC.n15167 185
R33038 VCC.n15142 VCC.n15141 185
R33039 VCC.n15141 VCC.n15140 185
R33040 VCC.n15184 VCC.n15183 185
R33041 VCC.n15185 VCC.n15184 185
R33042 VCC.n15139 VCC.n15137 185
R33043 VCC.n15187 VCC.n15139 185
R33044 VCC.n15318 VCC.n15317 185
R33045 VCC.n15319 VCC.n15318 185
R33046 VCC.n15051 VCC.n15050 185
R33047 VCC.n15354 VCC.n15051 185
R33048 VCC.n15375 VCC.n15374 185
R33049 VCC.n15376 VCC.n15375 185
R33050 VCC.n15373 VCC.n15039 185
R33051 VCC.n15377 VCC.n15039 185
R33052 VCC.n15357 VCC.n15356 185
R33053 VCC.n15356 VCC.n15355 185
R33054 VCC.n15386 VCC.n15040 185
R33055 VCC.n15080 VCC.n15079 185
R33056 VCC.n15078 VCC.n15077 185
R33057 VCC.n15295 VCC.n15078 185
R33058 VCC.n15298 VCC.n15297 185
R33059 VCC.n15297 VCC.n15296 185
R33060 VCC.n15066 VCC.n15065 185
R33061 VCC.n15320 VCC.n15066 185
R33062 VCC.n15380 VCC.n15015 185
R33063 VCC.n15378 VCC.n15015 185
R33064 VCC.n15014 VCC.n15013 185
R33065 VCC.n15430 VCC.n15014 185
R33066 VCC.n15451 VCC.n15450 185
R33067 VCC.n15451 VCC.n15000 185
R33068 VCC.n14983 VCC.n14982 185
R33069 VCC.n14982 VCC.n14981 185
R33070 VCC.n15488 VCC.n15487 185
R33071 VCC.n15487 VCC.n15486 185
R33072 VCC.n15507 VCC.n15506 185
R33073 VCC.n15508 VCC.n15507 185
R33074 VCC.n15457 VCC.n15456 185
R33075 VCC.n15456 VCC.n15455 185
R33076 VCC.n15434 VCC.n15433 185
R33077 VCC.n15433 VCC.n15432 185
R33078 VCC.n15452 VCC.n14998 185
R33079 VCC.n15453 VCC.n15452 185
R33080 VCC.n14980 VCC.n14979 185
R33081 VCC.n15485 VCC.n14980 185
R33082 VCC.n14965 VCC.n14964 185
R33083 VCC.n15382 VCC.n15381 185
R33084 VCC.n15382 VCC.n15379 185
R33085 VCC.n15937 VCC.n15936 185
R33086 VCC.n15936 VCC.n15935 185
R33087 VCC.n15985 VCC.n15984 185
R33088 VCC.n15986 VCC.n15985 185
R33089 VCC.n15568 VCC.n15566 185
R33090 VCC.n15990 VCC.n15568 185
R33091 VCC.n15548 VCC.n15541 185
R33092 VCC.n16026 VCC.n15548 185
R33093 VCC.n16056 VCC.n16055 185
R33094 VCC.n16057 VCC.n16056 185
R33095 VCC.n16060 VCC.n15518 185
R33096 VCC.n16060 VCC.n16059 185
R33097 VCC.n15522 VCC.n15521 185
R33098 VCC.n15521 VCC.n15520 185
R33099 VCC.n16024 VCC.n16023 185
R33100 VCC.n16025 VCC.n16024 185
R33101 VCC.n15988 VCC.n15551 185
R33102 VCC.n15989 VCC.n15988 185
R33103 VCC.n15567 VCC.n15565 185
R33104 VCC.n15987 VCC.n15567 185
R33105 VCC.n16062 VCC.n16061 185
R33106 VCC.n15939 VCC.n15938 185
R33107 VCC.n15939 VCC.n15934 185
R33108 VCC.n15854 VCC.n15853 185
R33109 VCC.n15853 VCC.n15852 185
R33110 VCC.n15622 VCC.n15621 185
R33111 VCC.n15876 VCC.n15622 185
R33112 VCC.n15607 VCC.n15606 185
R33113 VCC.n15910 VCC.n15607 185
R33114 VCC.n15931 VCC.n15930 185
R33115 VCC.n15932 VCC.n15931 185
R33116 VCC.n15929 VCC.n15595 185
R33117 VCC.n15933 VCC.n15595 185
R33118 VCC.n15874 VCC.n15873 185
R33119 VCC.n15875 VCC.n15874 185
R33120 VCC.n15634 VCC.n15633 185
R33121 VCC.n15851 VCC.n15634 185
R33122 VCC.n15913 VCC.n15912 185
R33123 VCC.n15912 VCC.n15911 185
R33124 VCC.n15943 VCC.n15596 185
R33125 VCC.n15636 VCC.n15635 185
R33126 VCC.n15741 VCC.n15740 185
R33127 VCC.n15742 VCC.n15741 185
R33128 VCC.n15696 VCC.n15694 185
R33129 VCC.n15744 VCC.n15696 185
R33130 VCC.n15786 VCC.n15785 185
R33131 VCC.n15785 VCC.n15784 185
R33132 VCC.n15802 VCC.n15656 185
R33133 VCC.n15806 VCC.n15656 185
R33134 VCC.n15808 VCC.n15657 185
R33135 VCC.n15808 VCC.n15807 185
R33136 VCC.n15747 VCC.n15746 185
R33137 VCC.n15746 VCC.n15745 185
R33138 VCC.n15699 VCC.n15698 185
R33139 VCC.n15698 VCC.n15697 185
R33140 VCC.n15787 VCC.n15659 185
R33141 VCC.n15659 VCC.n15658 185
R33142 VCC.n15726 VCC.n15724 185
R33143 VCC.n16297 VCC.n16296 185
R33144 VCC.n16296 VCC.n16295 185
R33145 VCC.n16336 VCC.n16335 185
R33146 VCC.n16335 VCC.n16334 185
R33147 VCC.n16352 VCC.n16206 185
R33148 VCC.n16356 VCC.n16206 185
R33149 VCC.n16358 VCC.n16207 185
R33150 VCC.n16358 VCC.n16357 185
R33151 VCC.n16337 VCC.n16209 185
R33152 VCC.n16209 VCC.n16208 185
R33153 VCC.n16276 VCC.n16274 185
R33154 VCC.n16249 VCC.n16248 185
R33155 VCC.n16248 VCC.n16247 185
R33156 VCC.n16291 VCC.n16290 185
R33157 VCC.n16292 VCC.n16291 185
R33158 VCC.n16246 VCC.n16244 185
R33159 VCC.n16294 VCC.n16246 185
R33160 VCC.n16425 VCC.n16424 185
R33161 VCC.n16426 VCC.n16425 185
R33162 VCC.n16158 VCC.n16157 185
R33163 VCC.n16461 VCC.n16158 185
R33164 VCC.n16482 VCC.n16481 185
R33165 VCC.n16483 VCC.n16482 185
R33166 VCC.n16480 VCC.n16146 185
R33167 VCC.n16484 VCC.n16146 185
R33168 VCC.n16464 VCC.n16463 185
R33169 VCC.n16463 VCC.n16462 185
R33170 VCC.n16493 VCC.n16147 185
R33171 VCC.n16187 VCC.n16186 185
R33172 VCC.n16185 VCC.n16184 185
R33173 VCC.n16402 VCC.n16185 185
R33174 VCC.n16405 VCC.n16404 185
R33175 VCC.n16404 VCC.n16403 185
R33176 VCC.n16173 VCC.n16172 185
R33177 VCC.n16427 VCC.n16173 185
R33178 VCC.n16487 VCC.n16122 185
R33179 VCC.n16485 VCC.n16122 185
R33180 VCC.n16121 VCC.n16120 185
R33181 VCC.n16537 VCC.n16121 185
R33182 VCC.n16558 VCC.n16557 185
R33183 VCC.n16558 VCC.n16107 185
R33184 VCC.n16090 VCC.n16089 185
R33185 VCC.n16089 VCC.n16088 185
R33186 VCC.n16595 VCC.n16594 185
R33187 VCC.n16594 VCC.n16593 185
R33188 VCC.n16614 VCC.n16613 185
R33189 VCC.n16615 VCC.n16614 185
R33190 VCC.n16564 VCC.n16563 185
R33191 VCC.n16563 VCC.n16562 185
R33192 VCC.n16541 VCC.n16540 185
R33193 VCC.n16540 VCC.n16539 185
R33194 VCC.n16559 VCC.n16105 185
R33195 VCC.n16560 VCC.n16559 185
R33196 VCC.n16087 VCC.n16086 185
R33197 VCC.n16592 VCC.n16087 185
R33198 VCC.n16072 VCC.n16071 185
R33199 VCC.n16489 VCC.n16488 185
R33200 VCC.n16489 VCC.n16486 185
R33201 VCC.n17044 VCC.n17043 185
R33202 VCC.n17043 VCC.n17042 185
R33203 VCC.n17092 VCC.n17091 185
R33204 VCC.n17093 VCC.n17092 185
R33205 VCC.n16675 VCC.n16673 185
R33206 VCC.n17097 VCC.n16675 185
R33207 VCC.n16655 VCC.n16648 185
R33208 VCC.n17133 VCC.n16655 185
R33209 VCC.n17163 VCC.n17162 185
R33210 VCC.n17164 VCC.n17163 185
R33211 VCC.n17167 VCC.n16625 185
R33212 VCC.n17167 VCC.n17166 185
R33213 VCC.n16629 VCC.n16628 185
R33214 VCC.n16628 VCC.n16627 185
R33215 VCC.n17131 VCC.n17130 185
R33216 VCC.n17132 VCC.n17131 185
R33217 VCC.n17095 VCC.n16658 185
R33218 VCC.n17096 VCC.n17095 185
R33219 VCC.n16674 VCC.n16672 185
R33220 VCC.n17094 VCC.n16674 185
R33221 VCC.n17169 VCC.n17168 185
R33222 VCC.n17046 VCC.n17045 185
R33223 VCC.n17046 VCC.n17041 185
R33224 VCC.n16961 VCC.n16960 185
R33225 VCC.n16960 VCC.n16959 185
R33226 VCC.n16729 VCC.n16728 185
R33227 VCC.n16983 VCC.n16729 185
R33228 VCC.n16714 VCC.n16713 185
R33229 VCC.n17017 VCC.n16714 185
R33230 VCC.n17038 VCC.n17037 185
R33231 VCC.n17039 VCC.n17038 185
R33232 VCC.n17036 VCC.n16702 185
R33233 VCC.n17040 VCC.n16702 185
R33234 VCC.n16981 VCC.n16980 185
R33235 VCC.n16982 VCC.n16981 185
R33236 VCC.n16741 VCC.n16740 185
R33237 VCC.n16958 VCC.n16741 185
R33238 VCC.n17020 VCC.n17019 185
R33239 VCC.n17019 VCC.n17018 185
R33240 VCC.n17050 VCC.n16703 185
R33241 VCC.n16743 VCC.n16742 185
R33242 VCC.n16848 VCC.n16847 185
R33243 VCC.n16849 VCC.n16848 185
R33244 VCC.n16803 VCC.n16801 185
R33245 VCC.n16851 VCC.n16803 185
R33246 VCC.n16893 VCC.n16892 185
R33247 VCC.n16892 VCC.n16891 185
R33248 VCC.n16909 VCC.n16763 185
R33249 VCC.n16913 VCC.n16763 185
R33250 VCC.n16915 VCC.n16764 185
R33251 VCC.n16915 VCC.n16914 185
R33252 VCC.n16854 VCC.n16853 185
R33253 VCC.n16853 VCC.n16852 185
R33254 VCC.n16806 VCC.n16805 185
R33255 VCC.n16805 VCC.n16804 185
R33256 VCC.n16894 VCC.n16766 185
R33257 VCC.n16766 VCC.n16765 185
R33258 VCC.n16833 VCC.n16831 185
R33259 VCC.n17345 VCC.n17344 185
R33260 VCC.n17346 VCC.n17345 185
R33261 VCC.n17265 VCC.n17264 185
R33262 VCC.n17381 VCC.n17265 185
R33263 VCC.n17402 VCC.n17401 185
R33264 VCC.n17403 VCC.n17402 185
R33265 VCC.n17400 VCC.n17253 185
R33266 VCC.n17404 VCC.n17253 185
R33267 VCC.n17384 VCC.n17383 185
R33268 VCC.n17383 VCC.n17382 185
R33269 VCC.n17413 VCC.n17254 185
R33270 VCC.n17294 VCC.n17293 185
R33271 VCC.n17292 VCC.n17291 185
R33272 VCC.n17322 VCC.n17292 185
R33273 VCC.n17325 VCC.n17324 185
R33274 VCC.n17324 VCC.n17323 185
R33275 VCC.n17280 VCC.n17279 185
R33276 VCC.n17347 VCC.n17280 185
R33277 VCC.n17407 VCC.n17229 185
R33278 VCC.n17405 VCC.n17229 185
R33279 VCC.n17228 VCC.n17227 185
R33280 VCC.n17457 VCC.n17228 185
R33281 VCC.n17478 VCC.n17477 185
R33282 VCC.n17478 VCC.n17214 185
R33283 VCC.n17197 VCC.n17196 185
R33284 VCC.n17196 VCC.n17195 185
R33285 VCC.n17515 VCC.n17514 185
R33286 VCC.n17514 VCC.n17513 185
R33287 VCC.n17534 VCC.n17533 185
R33288 VCC.n17535 VCC.n17534 185
R33289 VCC.n17484 VCC.n17483 185
R33290 VCC.n17483 VCC.n17482 185
R33291 VCC.n17461 VCC.n17460 185
R33292 VCC.n17460 VCC.n17459 185
R33293 VCC.n17479 VCC.n17212 185
R33294 VCC.n17480 VCC.n17479 185
R33295 VCC.n17194 VCC.n17193 185
R33296 VCC.n17512 VCC.n17194 185
R33297 VCC.n17179 VCC.n17178 185
R33298 VCC.n17409 VCC.n17408 185
R33299 VCC.n17409 VCC.n17406 185
R33300 VCC.n229 VCC.n227 96.8274
R33301 VCC.n289 VCC.n142 96.8274
R33302 VCC.n360 VCC.n108 96.8274
R33303 VCC.n396 VCC.n82 96.8274
R33304 VCC.n781 VCC.n779 96.8274
R33305 VCC.n841 VCC.n694 96.8274
R33306 VCC.n912 VCC.n660 96.8274
R33307 VCC.n948 VCC.n634 96.8274
R33308 VCC.n1469 VCC.n1217 96.8274
R33309 VCC.n1505 VCC.n1191 96.8274
R33310 VCC.n1339 VCC.n1337 96.8274
R33311 VCC.n1399 VCC.n1252 96.8274
R33312 VCC.n1890 VCC.n1888 96.8274
R33313 VCC.n1950 VCC.n1803 96.8274
R33314 VCC.n2021 VCC.n1769 96.8274
R33315 VCC.n2057 VCC.n1743 96.8274
R33316 VCC.n2578 VCC.n2326 96.8274
R33317 VCC.n2614 VCC.n2300 96.8274
R33318 VCC.n2448 VCC.n2446 96.8274
R33319 VCC.n2508 VCC.n2361 96.8274
R33320 VCC.n2999 VCC.n2997 96.8274
R33321 VCC.n3059 VCC.n2912 96.8274
R33322 VCC.n3130 VCC.n2878 96.8274
R33323 VCC.n3166 VCC.n2852 96.8274
R33324 VCC.n3687 VCC.n3435 96.8274
R33325 VCC.n3723 VCC.n3409 96.8274
R33326 VCC.n3557 VCC.n3555 96.8274
R33327 VCC.n3617 VCC.n3470 96.8274
R33328 VCC.n4108 VCC.n4106 96.8274
R33329 VCC.n4168 VCC.n4021 96.8274
R33330 VCC.n4239 VCC.n3987 96.8274
R33331 VCC.n4275 VCC.n3961 96.8274
R33332 VCC.n4796 VCC.n4544 96.8274
R33333 VCC.n4832 VCC.n4518 96.8274
R33334 VCC.n4666 VCC.n4664 96.8274
R33335 VCC.n4726 VCC.n4579 96.8274
R33336 VCC.n5217 VCC.n5215 96.8274
R33337 VCC.n5277 VCC.n5130 96.8274
R33338 VCC.n5348 VCC.n5096 96.8274
R33339 VCC.n5384 VCC.n5070 96.8274
R33340 VCC.n5905 VCC.n5653 96.8274
R33341 VCC.n5941 VCC.n5627 96.8274
R33342 VCC.n5775 VCC.n5773 96.8274
R33343 VCC.n5835 VCC.n5688 96.8274
R33344 VCC.n6326 VCC.n6324 96.8274
R33345 VCC.n6386 VCC.n6239 96.8274
R33346 VCC.n6457 VCC.n6205 96.8274
R33347 VCC.n6493 VCC.n6179 96.8274
R33348 VCC.n7014 VCC.n6762 96.8274
R33349 VCC.n7050 VCC.n6736 96.8274
R33350 VCC.n6884 VCC.n6882 96.8274
R33351 VCC.n6944 VCC.n6797 96.8274
R33352 VCC.n7435 VCC.n7433 96.8274
R33353 VCC.n7495 VCC.n7348 96.8274
R33354 VCC.n7566 VCC.n7314 96.8274
R33355 VCC.n7602 VCC.n7288 96.8274
R33356 VCC.n8123 VCC.n7871 96.8274
R33357 VCC.n8159 VCC.n7845 96.8274
R33358 VCC.n7993 VCC.n7991 96.8274
R33359 VCC.n8053 VCC.n7906 96.8274
R33360 VCC.n8675 VCC.n8423 96.8274
R33361 VCC.n8711 VCC.n8397 96.8274
R33362 VCC.n8544 VCC.n8542 96.8274
R33363 VCC.n8604 VCC.n8457 96.8274
R33364 VCC.n9232 VCC.n8980 96.8274
R33365 VCC.n9268 VCC.n8954 96.8274
R33366 VCC.n9102 VCC.n9100 96.8274
R33367 VCC.n9162 VCC.n9015 96.8274
R33368 VCC.n9653 VCC.n9651 96.8274
R33369 VCC.n9713 VCC.n9566 96.8274
R33370 VCC.n9784 VCC.n9532 96.8274
R33371 VCC.n9820 VCC.n9506 96.8274
R33372 VCC.n10340 VCC.n10088 96.8274
R33373 VCC.n10376 VCC.n10062 96.8274
R33374 VCC.n10210 VCC.n10208 96.8274
R33375 VCC.n10270 VCC.n10123 96.8274
R33376 VCC.n10760 VCC.n10758 96.8274
R33377 VCC.n10820 VCC.n10673 96.8274
R33378 VCC.n10891 VCC.n10639 96.8274
R33379 VCC.n10927 VCC.n10613 96.8274
R33380 VCC.n11447 VCC.n11195 96.8274
R33381 VCC.n11483 VCC.n11169 96.8274
R33382 VCC.n11317 VCC.n11315 96.8274
R33383 VCC.n11377 VCC.n11230 96.8274
R33384 VCC.n11867 VCC.n11865 96.8274
R33385 VCC.n11927 VCC.n11780 96.8274
R33386 VCC.n11998 VCC.n11746 96.8274
R33387 VCC.n12034 VCC.n11720 96.8274
R33388 VCC.n12554 VCC.n12302 96.8274
R33389 VCC.n12590 VCC.n12276 96.8274
R33390 VCC.n12424 VCC.n12422 96.8274
R33391 VCC.n12484 VCC.n12337 96.8274
R33392 VCC.n12974 VCC.n12972 96.8274
R33393 VCC.n13034 VCC.n12887 96.8274
R33394 VCC.n13105 VCC.n12853 96.8274
R33395 VCC.n13141 VCC.n12827 96.8274
R33396 VCC.n13661 VCC.n13409 96.8274
R33397 VCC.n13697 VCC.n13383 96.8274
R33398 VCC.n13531 VCC.n13529 96.8274
R33399 VCC.n13591 VCC.n13444 96.8274
R33400 VCC.n14081 VCC.n14079 96.8274
R33401 VCC.n14141 VCC.n13994 96.8274
R33402 VCC.n14212 VCC.n13960 96.8274
R33403 VCC.n14248 VCC.n13934 96.8274
R33404 VCC.n14768 VCC.n14516 96.8274
R33405 VCC.n14804 VCC.n14490 96.8274
R33406 VCC.n14638 VCC.n14636 96.8274
R33407 VCC.n14698 VCC.n14551 96.8274
R33408 VCC.n15188 VCC.n15186 96.8274
R33409 VCC.n15248 VCC.n15101 96.8274
R33410 VCC.n15319 VCC.n15067 96.8274
R33411 VCC.n15355 VCC.n15041 96.8274
R33412 VCC.n15875 VCC.n15623 96.8274
R33413 VCC.n15911 VCC.n15597 96.8274
R33414 VCC.n15745 VCC.n15743 96.8274
R33415 VCC.n15805 VCC.n15658 96.8274
R33416 VCC.n16295 VCC.n16293 96.8274
R33417 VCC.n16355 VCC.n16208 96.8274
R33418 VCC.n16426 VCC.n16174 96.8274
R33419 VCC.n16462 VCC.n16148 96.8274
R33420 VCC.n16982 VCC.n16730 96.8274
R33421 VCC.n17018 VCC.n16704 96.8274
R33422 VCC.n16852 VCC.n16850 96.8274
R33423 VCC.n16912 VCC.n16765 96.8274
R33424 VCC.n17346 VCC.n17281 96.8274
R33425 VCC.n17382 VCC.n17255 96.8274
R33426 VCC.n266 VCC.n153 95.0005
R33427 VCC.n267 VCC.n266 95.0005
R33428 VCC.n362 VCC.n93 95.0005
R33429 VCC.n394 VCC.n93 95.0005
R33430 VCC.n818 VCC.n705 95.0005
R33431 VCC.n819 VCC.n818 95.0005
R33432 VCC.n914 VCC.n645 95.0005
R33433 VCC.n946 VCC.n645 95.0005
R33434 VCC.n1471 VCC.n1202 95.0005
R33435 VCC.n1503 VCC.n1202 95.0005
R33436 VCC.n1376 VCC.n1263 95.0005
R33437 VCC.n1377 VCC.n1376 95.0005
R33438 VCC.n1927 VCC.n1814 95.0005
R33439 VCC.n1928 VCC.n1927 95.0005
R33440 VCC.n2023 VCC.n1754 95.0005
R33441 VCC.n2055 VCC.n1754 95.0005
R33442 VCC.n2580 VCC.n2311 95.0005
R33443 VCC.n2612 VCC.n2311 95.0005
R33444 VCC.n2485 VCC.n2372 95.0005
R33445 VCC.n2486 VCC.n2485 95.0005
R33446 VCC.n3036 VCC.n2923 95.0005
R33447 VCC.n3037 VCC.n3036 95.0005
R33448 VCC.n3132 VCC.n2863 95.0005
R33449 VCC.n3164 VCC.n2863 95.0005
R33450 VCC.n3689 VCC.n3420 95.0005
R33451 VCC.n3721 VCC.n3420 95.0005
R33452 VCC.n3594 VCC.n3481 95.0005
R33453 VCC.n3595 VCC.n3594 95.0005
R33454 VCC.n4145 VCC.n4032 95.0005
R33455 VCC.n4146 VCC.n4145 95.0005
R33456 VCC.n4241 VCC.n3972 95.0005
R33457 VCC.n4273 VCC.n3972 95.0005
R33458 VCC.n4798 VCC.n4529 95.0005
R33459 VCC.n4830 VCC.n4529 95.0005
R33460 VCC.n4703 VCC.n4590 95.0005
R33461 VCC.n4704 VCC.n4703 95.0005
R33462 VCC.n5254 VCC.n5141 95.0005
R33463 VCC.n5255 VCC.n5254 95.0005
R33464 VCC.n5350 VCC.n5081 95.0005
R33465 VCC.n5382 VCC.n5081 95.0005
R33466 VCC.n5907 VCC.n5638 95.0005
R33467 VCC.n5939 VCC.n5638 95.0005
R33468 VCC.n5812 VCC.n5699 95.0005
R33469 VCC.n5813 VCC.n5812 95.0005
R33470 VCC.n6363 VCC.n6250 95.0005
R33471 VCC.n6364 VCC.n6363 95.0005
R33472 VCC.n6459 VCC.n6190 95.0005
R33473 VCC.n6491 VCC.n6190 95.0005
R33474 VCC.n7016 VCC.n6747 95.0005
R33475 VCC.n7048 VCC.n6747 95.0005
R33476 VCC.n6921 VCC.n6808 95.0005
R33477 VCC.n6922 VCC.n6921 95.0005
R33478 VCC.n7472 VCC.n7359 95.0005
R33479 VCC.n7473 VCC.n7472 95.0005
R33480 VCC.n7568 VCC.n7299 95.0005
R33481 VCC.n7600 VCC.n7299 95.0005
R33482 VCC.n8125 VCC.n7856 95.0005
R33483 VCC.n8157 VCC.n7856 95.0005
R33484 VCC.n8030 VCC.n7917 95.0005
R33485 VCC.n8031 VCC.n8030 95.0005
R33486 VCC.n8677 VCC.n8408 95.0005
R33487 VCC.n8709 VCC.n8408 95.0005
R33488 VCC.n8581 VCC.n8468 95.0005
R33489 VCC.n8582 VCC.n8581 95.0005
R33490 VCC.n9234 VCC.n8965 95.0005
R33491 VCC.n9266 VCC.n8965 95.0005
R33492 VCC.n9139 VCC.n9026 95.0005
R33493 VCC.n9140 VCC.n9139 95.0005
R33494 VCC.n9690 VCC.n9577 95.0005
R33495 VCC.n9691 VCC.n9690 95.0005
R33496 VCC.n9786 VCC.n9517 95.0005
R33497 VCC.n9818 VCC.n9517 95.0005
R33498 VCC.n10342 VCC.n10073 95.0005
R33499 VCC.n10374 VCC.n10073 95.0005
R33500 VCC.n10247 VCC.n10134 95.0005
R33501 VCC.n10248 VCC.n10247 95.0005
R33502 VCC.n10797 VCC.n10684 95.0005
R33503 VCC.n10798 VCC.n10797 95.0005
R33504 VCC.n10893 VCC.n10624 95.0005
R33505 VCC.n10925 VCC.n10624 95.0005
R33506 VCC.n11449 VCC.n11180 95.0005
R33507 VCC.n11481 VCC.n11180 95.0005
R33508 VCC.n11354 VCC.n11241 95.0005
R33509 VCC.n11355 VCC.n11354 95.0005
R33510 VCC.n11904 VCC.n11791 95.0005
R33511 VCC.n11905 VCC.n11904 95.0005
R33512 VCC.n12000 VCC.n11731 95.0005
R33513 VCC.n12032 VCC.n11731 95.0005
R33514 VCC.n12556 VCC.n12287 95.0005
R33515 VCC.n12588 VCC.n12287 95.0005
R33516 VCC.n12461 VCC.n12348 95.0005
R33517 VCC.n12462 VCC.n12461 95.0005
R33518 VCC.n13011 VCC.n12898 95.0005
R33519 VCC.n13012 VCC.n13011 95.0005
R33520 VCC.n13107 VCC.n12838 95.0005
R33521 VCC.n13139 VCC.n12838 95.0005
R33522 VCC.n13663 VCC.n13394 95.0005
R33523 VCC.n13695 VCC.n13394 95.0005
R33524 VCC.n13568 VCC.n13455 95.0005
R33525 VCC.n13569 VCC.n13568 95.0005
R33526 VCC.n14118 VCC.n14005 95.0005
R33527 VCC.n14119 VCC.n14118 95.0005
R33528 VCC.n14214 VCC.n13945 95.0005
R33529 VCC.n14246 VCC.n13945 95.0005
R33530 VCC.n14770 VCC.n14501 95.0005
R33531 VCC.n14802 VCC.n14501 95.0005
R33532 VCC.n14675 VCC.n14562 95.0005
R33533 VCC.n14676 VCC.n14675 95.0005
R33534 VCC.n15225 VCC.n15112 95.0005
R33535 VCC.n15226 VCC.n15225 95.0005
R33536 VCC.n15321 VCC.n15052 95.0005
R33537 VCC.n15353 VCC.n15052 95.0005
R33538 VCC.n15877 VCC.n15608 95.0005
R33539 VCC.n15909 VCC.n15608 95.0005
R33540 VCC.n15782 VCC.n15669 95.0005
R33541 VCC.n15783 VCC.n15782 95.0005
R33542 VCC.n16332 VCC.n16219 95.0005
R33543 VCC.n16333 VCC.n16332 95.0005
R33544 VCC.n16428 VCC.n16159 95.0005
R33545 VCC.n16460 VCC.n16159 95.0005
R33546 VCC.n16984 VCC.n16715 95.0005
R33547 VCC.n17016 VCC.n16715 95.0005
R33548 VCC.n16889 VCC.n16776 95.0005
R33549 VCC.n16890 VCC.n16889 95.0005
R33550 VCC.n17348 VCC.n17266 95.0005
R33551 VCC.n17380 VCC.n17266 95.0005
R33552 VCC.n473 VCC.n472 93.2412
R33553 VCC.n495 VCC.n494 93.2412
R33554 VCC.n496 VCC.n495 93.2412
R33555 VCC.n547 VCC.n5 93.2412
R33556 VCC.n1025 VCC.n1024 93.2412
R33557 VCC.n1047 VCC.n1046 93.2412
R33558 VCC.n1048 VCC.n1047 93.2412
R33559 VCC.n1101 VCC.n559 93.2412
R33560 VCC.n1585 VCC.n1581 93.2412
R33561 VCC.n1583 VCC.n1143 93.2412
R33562 VCC.n1619 VCC.n1143 93.2412
R33563 VCC.n1653 VCC.n1652 93.2412
R33564 VCC.n2134 VCC.n2133 93.2412
R33565 VCC.n2156 VCC.n2155 93.2412
R33566 VCC.n2157 VCC.n2156 93.2412
R33567 VCC.n2210 VCC.n1668 93.2412
R33568 VCC.n2694 VCC.n2690 93.2412
R33569 VCC.n2692 VCC.n2252 93.2412
R33570 VCC.n2728 VCC.n2252 93.2412
R33571 VCC.n2762 VCC.n2761 93.2412
R33572 VCC.n3243 VCC.n3242 93.2412
R33573 VCC.n3265 VCC.n3264 93.2412
R33574 VCC.n3266 VCC.n3265 93.2412
R33575 VCC.n3319 VCC.n2777 93.2412
R33576 VCC.n3803 VCC.n3799 93.2412
R33577 VCC.n3801 VCC.n3361 93.2412
R33578 VCC.n3837 VCC.n3361 93.2412
R33579 VCC.n3871 VCC.n3870 93.2412
R33580 VCC.n4352 VCC.n4351 93.2412
R33581 VCC.n4374 VCC.n4373 93.2412
R33582 VCC.n4375 VCC.n4374 93.2412
R33583 VCC.n4428 VCC.n3886 93.2412
R33584 VCC.n4912 VCC.n4908 93.2412
R33585 VCC.n4910 VCC.n4470 93.2412
R33586 VCC.n4946 VCC.n4470 93.2412
R33587 VCC.n4980 VCC.n4979 93.2412
R33588 VCC.n5461 VCC.n5460 93.2412
R33589 VCC.n5483 VCC.n5482 93.2412
R33590 VCC.n5484 VCC.n5483 93.2412
R33591 VCC.n5537 VCC.n4995 93.2412
R33592 VCC.n6021 VCC.n6017 93.2412
R33593 VCC.n6019 VCC.n5579 93.2412
R33594 VCC.n6055 VCC.n5579 93.2412
R33595 VCC.n6089 VCC.n6088 93.2412
R33596 VCC.n6570 VCC.n6569 93.2412
R33597 VCC.n6592 VCC.n6591 93.2412
R33598 VCC.n6593 VCC.n6592 93.2412
R33599 VCC.n6646 VCC.n6104 93.2412
R33600 VCC.n7130 VCC.n7126 93.2412
R33601 VCC.n7128 VCC.n6688 93.2412
R33602 VCC.n7164 VCC.n6688 93.2412
R33603 VCC.n7198 VCC.n7197 93.2412
R33604 VCC.n7679 VCC.n7678 93.2412
R33605 VCC.n7701 VCC.n7700 93.2412
R33606 VCC.n7702 VCC.n7701 93.2412
R33607 VCC.n7755 VCC.n7213 93.2412
R33608 VCC.n8239 VCC.n8235 93.2412
R33609 VCC.n8237 VCC.n7797 93.2412
R33610 VCC.n8273 VCC.n7797 93.2412
R33611 VCC.n8307 VCC.n8306 93.2412
R33612 VCC.n8788 VCC.n8787 93.2412
R33613 VCC.n8810 VCC.n8809 93.2412
R33614 VCC.n8811 VCC.n8810 93.2412
R33615 VCC.n8864 VCC.n8322 93.2412
R33616 VCC.n9348 VCC.n9344 93.2412
R33617 VCC.n9346 VCC.n8906 93.2412
R33618 VCC.n9382 VCC.n8906 93.2412
R33619 VCC.n9416 VCC.n9415 93.2412
R33620 VCC.n9897 VCC.n9896 93.2412
R33621 VCC.n9919 VCC.n9918 93.2412
R33622 VCC.n9920 VCC.n9919 93.2412
R33623 VCC.n9973 VCC.n9431 93.2412
R33624 VCC.n10456 VCC.n10452 93.2412
R33625 VCC.n10454 VCC.n10014 93.2412
R33626 VCC.n10490 VCC.n10014 93.2412
R33627 VCC.n10524 VCC.n10523 93.2412
R33628 VCC.n11004 VCC.n11003 93.2412
R33629 VCC.n11026 VCC.n11025 93.2412
R33630 VCC.n11027 VCC.n11026 93.2412
R33631 VCC.n11080 VCC.n10538 93.2412
R33632 VCC.n11563 VCC.n11559 93.2412
R33633 VCC.n11561 VCC.n11121 93.2412
R33634 VCC.n11597 VCC.n11121 93.2412
R33635 VCC.n11631 VCC.n11630 93.2412
R33636 VCC.n12111 VCC.n12110 93.2412
R33637 VCC.n12133 VCC.n12132 93.2412
R33638 VCC.n12134 VCC.n12133 93.2412
R33639 VCC.n12187 VCC.n11645 93.2412
R33640 VCC.n12670 VCC.n12666 93.2412
R33641 VCC.n12668 VCC.n12228 93.2412
R33642 VCC.n12704 VCC.n12228 93.2412
R33643 VCC.n12738 VCC.n12737 93.2412
R33644 VCC.n13218 VCC.n13217 93.2412
R33645 VCC.n13240 VCC.n13239 93.2412
R33646 VCC.n13241 VCC.n13240 93.2412
R33647 VCC.n13294 VCC.n12752 93.2412
R33648 VCC.n13777 VCC.n13773 93.2412
R33649 VCC.n13775 VCC.n13335 93.2412
R33650 VCC.n13811 VCC.n13335 93.2412
R33651 VCC.n13845 VCC.n13844 93.2412
R33652 VCC.n14325 VCC.n14324 93.2412
R33653 VCC.n14347 VCC.n14346 93.2412
R33654 VCC.n14348 VCC.n14347 93.2412
R33655 VCC.n14401 VCC.n13859 93.2412
R33656 VCC.n14884 VCC.n14880 93.2412
R33657 VCC.n14882 VCC.n14442 93.2412
R33658 VCC.n14918 VCC.n14442 93.2412
R33659 VCC.n14952 VCC.n14951 93.2412
R33660 VCC.n15432 VCC.n15431 93.2412
R33661 VCC.n15454 VCC.n15453 93.2412
R33662 VCC.n15455 VCC.n15454 93.2412
R33663 VCC.n15508 VCC.n14966 93.2412
R33664 VCC.n15991 VCC.n15987 93.2412
R33665 VCC.n15989 VCC.n15549 93.2412
R33666 VCC.n16025 VCC.n15549 93.2412
R33667 VCC.n16059 VCC.n16058 93.2412
R33668 VCC.n16539 VCC.n16538 93.2412
R33669 VCC.n16561 VCC.n16560 93.2412
R33670 VCC.n16562 VCC.n16561 93.2412
R33671 VCC.n16615 VCC.n16073 93.2412
R33672 VCC.n17098 VCC.n17094 93.2412
R33673 VCC.n17096 VCC.n16656 93.2412
R33674 VCC.n17132 VCC.n16656 93.2412
R33675 VCC.n17166 VCC.n17165 93.2412
R33676 VCC.n17459 VCC.n17458 93.2412
R33677 VCC.n17481 VCC.n17480 93.2412
R33678 VCC.n17482 VCC.n17481 93.2412
R33679 VCC.n17535 VCC.n17180 93.2412
R33680 VCC.n213 VCC.n194 92.5398
R33681 VCC.n333 VCC.n123 92.5398
R33682 VCC.n430 VCC.n79 92.5398
R33683 VCC.n765 VCC.n746 92.5398
R33684 VCC.n885 VCC.n675 92.5398
R33685 VCC.n982 VCC.n631 92.5398
R33686 VCC.n1442 VCC.n1232 92.5398
R33687 VCC.n1540 VCC.n1188 92.5398
R33688 VCC.n1323 VCC.n1304 92.5398
R33689 VCC.n1874 VCC.n1855 92.5398
R33690 VCC.n1994 VCC.n1784 92.5398
R33691 VCC.n2091 VCC.n1740 92.5398
R33692 VCC.n2551 VCC.n2341 92.5398
R33693 VCC.n2649 VCC.n2297 92.5398
R33694 VCC.n2432 VCC.n2413 92.5398
R33695 VCC.n2983 VCC.n2964 92.5398
R33696 VCC.n3103 VCC.n2893 92.5398
R33697 VCC.n3200 VCC.n2849 92.5398
R33698 VCC.n3660 VCC.n3450 92.5398
R33699 VCC.n3758 VCC.n3406 92.5398
R33700 VCC.n3541 VCC.n3522 92.5398
R33701 VCC.n4092 VCC.n4073 92.5398
R33702 VCC.n4212 VCC.n4002 92.5398
R33703 VCC.n4309 VCC.n3958 92.5398
R33704 VCC.n4769 VCC.n4559 92.5398
R33705 VCC.n4867 VCC.n4515 92.5398
R33706 VCC.n4650 VCC.n4631 92.5398
R33707 VCC.n5201 VCC.n5182 92.5398
R33708 VCC.n5321 VCC.n5111 92.5398
R33709 VCC.n5418 VCC.n5067 92.5398
R33710 VCC.n5878 VCC.n5668 92.5398
R33711 VCC.n5976 VCC.n5624 92.5398
R33712 VCC.n5759 VCC.n5740 92.5398
R33713 VCC.n6310 VCC.n6291 92.5398
R33714 VCC.n6430 VCC.n6220 92.5398
R33715 VCC.n6527 VCC.n6176 92.5398
R33716 VCC.n6987 VCC.n6777 92.5398
R33717 VCC.n7085 VCC.n6733 92.5398
R33718 VCC.n6868 VCC.n6849 92.5398
R33719 VCC.n7419 VCC.n7400 92.5398
R33720 VCC.n7539 VCC.n7329 92.5398
R33721 VCC.n7636 VCC.n7285 92.5398
R33722 VCC.n8096 VCC.n7886 92.5398
R33723 VCC.n8194 VCC.n7842 92.5398
R33724 VCC.n7977 VCC.n7958 92.5398
R33725 VCC.n8648 VCC.n8438 92.5398
R33726 VCC.n8745 VCC.n8394 92.5398
R33727 VCC.n8528 VCC.n8509 92.5398
R33728 VCC.n9205 VCC.n8995 92.5398
R33729 VCC.n9303 VCC.n8951 92.5398
R33730 VCC.n9086 VCC.n9067 92.5398
R33731 VCC.n9637 VCC.n9618 92.5398
R33732 VCC.n9757 VCC.n9547 92.5398
R33733 VCC.n9854 VCC.n9503 92.5398
R33734 VCC.n10313 VCC.n10103 92.5398
R33735 VCC.n10411 VCC.n10059 92.5398
R33736 VCC.n10194 VCC.n10175 92.5398
R33737 VCC.n10744 VCC.n10725 92.5398
R33738 VCC.n10864 VCC.n10654 92.5398
R33739 VCC.n10961 VCC.n10610 92.5398
R33740 VCC.n11420 VCC.n11210 92.5398
R33741 VCC.n11518 VCC.n11166 92.5398
R33742 VCC.n11301 VCC.n11282 92.5398
R33743 VCC.n11851 VCC.n11832 92.5398
R33744 VCC.n11971 VCC.n11761 92.5398
R33745 VCC.n12068 VCC.n11717 92.5398
R33746 VCC.n12527 VCC.n12317 92.5398
R33747 VCC.n12625 VCC.n12273 92.5398
R33748 VCC.n12408 VCC.n12389 92.5398
R33749 VCC.n12958 VCC.n12939 92.5398
R33750 VCC.n13078 VCC.n12868 92.5398
R33751 VCC.n13175 VCC.n12824 92.5398
R33752 VCC.n13634 VCC.n13424 92.5398
R33753 VCC.n13732 VCC.n13380 92.5398
R33754 VCC.n13515 VCC.n13496 92.5398
R33755 VCC.n14065 VCC.n14046 92.5398
R33756 VCC.n14185 VCC.n13975 92.5398
R33757 VCC.n14282 VCC.n13931 92.5398
R33758 VCC.n14741 VCC.n14531 92.5398
R33759 VCC.n14839 VCC.n14487 92.5398
R33760 VCC.n14622 VCC.n14603 92.5398
R33761 VCC.n15172 VCC.n15153 92.5398
R33762 VCC.n15292 VCC.n15082 92.5398
R33763 VCC.n15389 VCC.n15038 92.5398
R33764 VCC.n15848 VCC.n15638 92.5398
R33765 VCC.n15946 VCC.n15594 92.5398
R33766 VCC.n15729 VCC.n15710 92.5398
R33767 VCC.n16279 VCC.n16260 92.5398
R33768 VCC.n16399 VCC.n16189 92.5398
R33769 VCC.n16496 VCC.n16145 92.5398
R33770 VCC.n16955 VCC.n16745 92.5398
R33771 VCC.n17053 VCC.n16701 92.5398
R33772 VCC.n16836 VCC.n16817 92.5398
R33773 VCC.n17319 VCC.n17296 92.5398
R33774 VCC.n17416 VCC.n17252 92.5398
R33775 VCC.n265 VCC.n264 92.5005
R33776 VCC.n266 VCC.n265 92.5005
R33777 VCC.n385 VCC.n94 92.5005
R33778 VCC.n94 VCC.n93 92.5005
R33779 VCC.n817 VCC.n816 92.5005
R33780 VCC.n818 VCC.n817 92.5005
R33781 VCC.n937 VCC.n646 92.5005
R33782 VCC.n646 VCC.n645 92.5005
R33783 VCC.n1494 VCC.n1203 92.5005
R33784 VCC.n1203 VCC.n1202 92.5005
R33785 VCC.n1375 VCC.n1374 92.5005
R33786 VCC.n1376 VCC.n1375 92.5005
R33787 VCC.n1926 VCC.n1925 92.5005
R33788 VCC.n1927 VCC.n1926 92.5005
R33789 VCC.n2046 VCC.n1755 92.5005
R33790 VCC.n1755 VCC.n1754 92.5005
R33791 VCC.n2603 VCC.n2312 92.5005
R33792 VCC.n2312 VCC.n2311 92.5005
R33793 VCC.n2484 VCC.n2483 92.5005
R33794 VCC.n2485 VCC.n2484 92.5005
R33795 VCC.n3035 VCC.n3034 92.5005
R33796 VCC.n3036 VCC.n3035 92.5005
R33797 VCC.n3155 VCC.n2864 92.5005
R33798 VCC.n2864 VCC.n2863 92.5005
R33799 VCC.n3712 VCC.n3421 92.5005
R33800 VCC.n3421 VCC.n3420 92.5005
R33801 VCC.n3593 VCC.n3592 92.5005
R33802 VCC.n3594 VCC.n3593 92.5005
R33803 VCC.n4144 VCC.n4143 92.5005
R33804 VCC.n4145 VCC.n4144 92.5005
R33805 VCC.n4264 VCC.n3973 92.5005
R33806 VCC.n3973 VCC.n3972 92.5005
R33807 VCC.n4821 VCC.n4530 92.5005
R33808 VCC.n4530 VCC.n4529 92.5005
R33809 VCC.n4702 VCC.n4701 92.5005
R33810 VCC.n4703 VCC.n4702 92.5005
R33811 VCC.n5253 VCC.n5252 92.5005
R33812 VCC.n5254 VCC.n5253 92.5005
R33813 VCC.n5373 VCC.n5082 92.5005
R33814 VCC.n5082 VCC.n5081 92.5005
R33815 VCC.n5930 VCC.n5639 92.5005
R33816 VCC.n5639 VCC.n5638 92.5005
R33817 VCC.n5811 VCC.n5810 92.5005
R33818 VCC.n5812 VCC.n5811 92.5005
R33819 VCC.n6362 VCC.n6361 92.5005
R33820 VCC.n6363 VCC.n6362 92.5005
R33821 VCC.n6482 VCC.n6191 92.5005
R33822 VCC.n6191 VCC.n6190 92.5005
R33823 VCC.n7039 VCC.n6748 92.5005
R33824 VCC.n6748 VCC.n6747 92.5005
R33825 VCC.n6920 VCC.n6919 92.5005
R33826 VCC.n6921 VCC.n6920 92.5005
R33827 VCC.n7471 VCC.n7470 92.5005
R33828 VCC.n7472 VCC.n7471 92.5005
R33829 VCC.n7591 VCC.n7300 92.5005
R33830 VCC.n7300 VCC.n7299 92.5005
R33831 VCC.n8148 VCC.n7857 92.5005
R33832 VCC.n7857 VCC.n7856 92.5005
R33833 VCC.n8029 VCC.n8028 92.5005
R33834 VCC.n8030 VCC.n8029 92.5005
R33835 VCC.n8700 VCC.n8409 92.5005
R33836 VCC.n8409 VCC.n8408 92.5005
R33837 VCC.n8580 VCC.n8579 92.5005
R33838 VCC.n8581 VCC.n8580 92.5005
R33839 VCC.n9257 VCC.n8966 92.5005
R33840 VCC.n8966 VCC.n8965 92.5005
R33841 VCC.n9138 VCC.n9137 92.5005
R33842 VCC.n9139 VCC.n9138 92.5005
R33843 VCC.n9689 VCC.n9688 92.5005
R33844 VCC.n9690 VCC.n9689 92.5005
R33845 VCC.n9809 VCC.n9518 92.5005
R33846 VCC.n9518 VCC.n9517 92.5005
R33847 VCC.n10365 VCC.n10074 92.5005
R33848 VCC.n10074 VCC.n10073 92.5005
R33849 VCC.n10246 VCC.n10245 92.5005
R33850 VCC.n10247 VCC.n10246 92.5005
R33851 VCC.n10796 VCC.n10795 92.5005
R33852 VCC.n10797 VCC.n10796 92.5005
R33853 VCC.n10916 VCC.n10625 92.5005
R33854 VCC.n10625 VCC.n10624 92.5005
R33855 VCC.n11472 VCC.n11181 92.5005
R33856 VCC.n11181 VCC.n11180 92.5005
R33857 VCC.n11353 VCC.n11352 92.5005
R33858 VCC.n11354 VCC.n11353 92.5005
R33859 VCC.n11903 VCC.n11902 92.5005
R33860 VCC.n11904 VCC.n11903 92.5005
R33861 VCC.n12023 VCC.n11732 92.5005
R33862 VCC.n11732 VCC.n11731 92.5005
R33863 VCC.n12579 VCC.n12288 92.5005
R33864 VCC.n12288 VCC.n12287 92.5005
R33865 VCC.n12460 VCC.n12459 92.5005
R33866 VCC.n12461 VCC.n12460 92.5005
R33867 VCC.n13010 VCC.n13009 92.5005
R33868 VCC.n13011 VCC.n13010 92.5005
R33869 VCC.n13130 VCC.n12839 92.5005
R33870 VCC.n12839 VCC.n12838 92.5005
R33871 VCC.n13686 VCC.n13395 92.5005
R33872 VCC.n13395 VCC.n13394 92.5005
R33873 VCC.n13567 VCC.n13566 92.5005
R33874 VCC.n13568 VCC.n13567 92.5005
R33875 VCC.n14117 VCC.n14116 92.5005
R33876 VCC.n14118 VCC.n14117 92.5005
R33877 VCC.n14237 VCC.n13946 92.5005
R33878 VCC.n13946 VCC.n13945 92.5005
R33879 VCC.n14793 VCC.n14502 92.5005
R33880 VCC.n14502 VCC.n14501 92.5005
R33881 VCC.n14674 VCC.n14673 92.5005
R33882 VCC.n14675 VCC.n14674 92.5005
R33883 VCC.n15224 VCC.n15223 92.5005
R33884 VCC.n15225 VCC.n15224 92.5005
R33885 VCC.n15344 VCC.n15053 92.5005
R33886 VCC.n15053 VCC.n15052 92.5005
R33887 VCC.n15900 VCC.n15609 92.5005
R33888 VCC.n15609 VCC.n15608 92.5005
R33889 VCC.n15781 VCC.n15780 92.5005
R33890 VCC.n15782 VCC.n15781 92.5005
R33891 VCC.n16331 VCC.n16330 92.5005
R33892 VCC.n16332 VCC.n16331 92.5005
R33893 VCC.n16451 VCC.n16160 92.5005
R33894 VCC.n16160 VCC.n16159 92.5005
R33895 VCC.n17007 VCC.n16716 92.5005
R33896 VCC.n16716 VCC.n16715 92.5005
R33897 VCC.n16888 VCC.n16887 92.5005
R33898 VCC.n16889 VCC.n16888 92.5005
R33899 VCC.n17371 VCC.n17267 92.5005
R33900 VCC.n17267 VCC.n17266 92.5005
R33901 VCC.n211 VCC.t232 74.9043
R33902 VCC.n763 VCC.t387 74.9043
R33903 VCC.n1321 VCC.t485 74.9043
R33904 VCC.n1872 VCC.t18 74.9043
R33905 VCC.n2430 VCC.t141 74.9043
R33906 VCC.n2981 VCC.t599 74.9043
R33907 VCC.n3539 VCC.t4 74.9043
R33908 VCC.n4090 VCC.t551 74.9043
R33909 VCC.n4648 VCC.t412 74.9043
R33910 VCC.n5199 VCC.t350 74.9043
R33911 VCC.n5757 VCC.t621 74.9043
R33912 VCC.n6308 VCC.t332 74.9043
R33913 VCC.n6866 VCC.t235 74.9043
R33914 VCC.n7417 VCC.t601 74.9043
R33915 VCC.n7975 VCC.t105 74.9043
R33916 VCC.n8526 VCC.t83 74.9043
R33917 VCC.n9084 VCC.t422 74.9043
R33918 VCC.n9635 VCC.t321 74.9043
R33919 VCC.n10192 VCC.t47 74.9043
R33920 VCC.n10742 VCC.t22 74.9043
R33921 VCC.n11299 VCC.t228 74.9043
R33922 VCC.n11849 VCC.t505 74.9043
R33923 VCC.n12406 VCC.t261 74.9043
R33924 VCC.n12956 VCC.t560 74.9043
R33925 VCC.n13513 VCC.t628 74.9043
R33926 VCC.n14063 VCC.t208 74.9043
R33927 VCC.n14620 VCC.t353 74.9043
R33928 VCC.n15170 VCC.t50 74.9043
R33929 VCC.n15727 VCC.t527 74.9043
R33930 VCC.n16277 VCC.t419 74.9043
R33931 VCC.n16834 VCC.t608 74.9043
R33932 VCC.t567 VCC.n335 73.0774
R33933 VCC.t390 VCC.n887 73.0774
R33934 VCC.t296 VCC.n1444 73.0774
R33935 VCC.t553 VCC.n1996 73.0774
R33936 VCC.t479 VCC.n2553 73.0774
R33937 VCC.t327 VCC.n3105 73.0774
R33938 VCC.t161 VCC.n3662 73.0774
R33939 VCC.t158 VCC.n4214 73.0774
R33940 VCC.t443 VCC.n4771 73.0774
R33941 VCC.t101 VCC.n5323 73.0774
R33942 VCC.t250 VCC.n5880 73.0774
R33943 VCC.t148 VCC.n6432 73.0774
R33944 VCC.t202 VCC.n6989 73.0774
R33945 VCC.t96 VCC.n7541 73.0774
R33946 VCC.t125 VCC.n8098 73.0774
R33947 VCC.t475 VCC.n8650 73.0774
R33948 VCC.t275 VCC.n9207 73.0774
R33949 VCC.t482 VCC.n9759 73.0774
R33950 VCC.t542 VCC.n10315 73.0774
R33951 VCC.t219 VCC.n10866 73.0774
R33952 VCC.t452 VCC.n11422 73.0774
R33953 VCC.t87 VCC.n11973 73.0774
R33954 VCC.t547 VCC.n12529 73.0774
R33955 VCC.t212 VCC.n13080 73.0774
R33956 VCC.t309 VCC.n13636 73.0774
R33957 VCC.t586 VCC.n14187 73.0774
R33958 VCC.t131 VCC.n14743 73.0774
R33959 VCC.t340 VCC.n15294 73.0774
R33960 VCC.t8 VCC.n15850 73.0774
R33961 VCC.t518 VCC.n16401 73.0774
R33962 VCC.t347 VCC.n16957 73.0774
R33963 VCC.t369 VCC.n17321 73.0774
R33964 VCC.n293 VCC.t10 72.544
R33965 VCC.n845 VCC.t20 72.544
R33966 VCC.n1403 VCC.t466 72.544
R33967 VCC.n1954 VCC.t367 72.544
R33968 VCC.n2512 VCC.t432 72.544
R33969 VCC.n3063 VCC.t468 72.544
R33970 VCC.n3621 VCC.t399 72.544
R33971 VCC.n4172 VCC.t365 72.544
R33972 VCC.n4730 VCC.t362 72.544
R33973 VCC.n5281 VCC.t195 72.544
R33974 VCC.n5839 VCC.t618 72.544
R33975 VCC.n6390 VCC.t596 72.544
R33976 VCC.n6948 VCC.t531 72.544
R33977 VCC.n7499 VCC.t300 72.544
R33978 VCC.n8057 VCC.t632 72.544
R33979 VCC.n8608 VCC.t247 72.544
R33980 VCC.n9166 VCC.t108 72.544
R33981 VCC.n9717 VCC.t272 72.544
R33982 VCC.n10274 VCC.t424 72.544
R33983 VCC.n10824 VCC.t616 72.544
R33984 VCC.n11381 VCC.t380 72.544
R33985 VCC.n11931 VCC.t151 72.544
R33986 VCC.n12488 VCC.t192 72.544
R33987 VCC.n13038 VCC.t318 72.544
R33988 VCC.n13595 VCC.t263 72.544
R33989 VCC.n14145 VCC.t114 72.544
R33990 VCC.n14702 VCC.t206 72.544
R33991 VCC.n15252 VCC.t92 72.544
R33992 VCC.n15809 VCC.t525 72.544
R33993 VCC.n16359 VCC.t253 72.544
R33994 VCC.n16916 VCC.t407 72.544
R33995 VCC.t330 VCC.n525 70.3709
R33996 VCC.t185 VCC.n1077 70.3709
R33997 VCC.n1621 VCC.t343 70.3709
R33998 VCC.t434 VCC.n2186 70.3709
R33999 VCC.n2730 VCC.t111 70.3709
R34000 VCC.t372 VCC.n3295 70.3709
R34001 VCC.n3839 VCC.t155 70.3709
R34002 VCC.t38 VCC.n4404 70.3709
R34003 VCC.n4948 VCC.t459 70.3709
R34004 VCC.t0 VCC.n5513 70.3709
R34005 VCC.n6057 VCC.t440 70.3709
R34006 VCC.t256 VCC.n6622 70.3709
R34007 VCC.n7166 VCC.t53 70.3709
R34008 VCC.t168 VCC.n7731 70.3709
R34009 VCC.n8275 VCC.t376 70.3709
R34010 VCC.t446 VCC.n8840 70.3709
R34011 VCC.n9384 VCC.t402 70.3709
R34012 VCC.t494 VCC.n9949 70.3709
R34013 VCC.n10492 VCC.t356 70.3709
R34014 VCC.t31 VCC.n11056 70.3709
R34015 VCC.n11599 VCC.t14 70.3709
R34016 VCC.t501 VCC.n12163 70.3709
R34017 VCC.n12706 VCC.t397 70.3709
R34018 VCC.t267 VCC.n13270 70.3709
R34019 VCC.n13813 VCC.t134 70.3709
R34020 VCC.t571 VCC.n14377 70.3709
R34021 VCC.n14920 VCC.t472 70.3709
R34022 VCC.t507 VCC.n15484 70.3709
R34023 VCC.n16027 VCC.t58 70.3709
R34024 VCC.t174 VCC.n16591 70.3709
R34025 VCC.n17134 VCC.t565 70.3709
R34026 VCC.t624 VCC.n17511 70.3709
R34027 VCC.n470 VCC.t189 66.8524
R34028 VCC.n1022 VCC.t336 66.8524
R34029 VCC.t286 VCC.n1163 66.8524
R34030 VCC.n2131 VCC.t428 66.8524
R34031 VCC.t290 VCC.n2272 66.8524
R34032 VCC.n3240 VCC.t589 66.8524
R34033 VCC.t574 VCC.n3381 66.8524
R34034 VCC.n4349 VCC.t315 66.8524
R34035 VCC.t533 VCC.n4490 66.8524
R34036 VCC.n5458 VCC.t324 66.8524
R34037 VCC.t25 VCC.n5599 66.8524
R34038 VCC.n6567 VCC.t306 66.8524
R34039 VCC.t225 VCC.n6708 66.8524
R34040 VCC.n7676 VCC.t582 66.8524
R34041 VCC.t279 VCC.n7817 66.8524
R34042 VCC.n8785 VCC.t33 66.8524
R34043 VCC.t538 VCC.n8926 66.8524
R34044 VCC.n9894 VCC.t497 66.8524
R34045 VCC.t237 VCC.n10034 66.8524
R34046 VCC.n11001 VCC.t612 66.8524
R34047 VCC.t117 VCC.n11141 66.8524
R34048 VCC.n12108 VCC.t215 66.8524
R34049 VCC.t178 VCC.n12248 66.8524
R34050 VCC.n13215 VCC.t511 66.8524
R34051 VCC.t606 VCC.n13355 66.8524
R34052 VCC.n14322 VCC.t462 66.8524
R34053 VCC.t74 VCC.n14462 66.8524
R34054 VCC.n15429 VCC.t558 66.8524
R34055 VCC.t488 VCC.n15569 66.8524
R34056 VCC.n16536 VCC.t592 66.8524
R34057 VCC.t122 VCC.n16676 66.8524
R34058 VCC.n17456 VCC.t198 66.8524
R34059 VCC.n428 VCC.t138 65.7697
R34060 VCC.n980 VCC.t128 65.7697
R34061 VCC.n1538 VCC.t64 65.7697
R34062 VCC.n2089 VCC.t384 65.7697
R34063 VCC.n2647 VCC.t409 65.7697
R34064 VCC.n3198 VCC.t182 65.7697
R34065 VCC.n3756 VCC.t521 65.7697
R34066 VCC.n4307 VCC.t163 65.7697
R34067 VCC.n4865 VCC.t42 65.7697
R34068 VCC.n5416 VCC.t170 65.7697
R34069 VCC.n5974 VCC.t221 65.7697
R34070 VCC.n6525 VCC.t241 65.7697
R34071 VCC.n7083 VCC.t392 65.7697
R34072 VCC.n7634 VCC.t515 65.7697
R34073 VCC.n8192 VCC.t98 65.7697
R34074 VCC.n8743 VCC.t61 65.7697
R34075 VCC.n9301 VCC.t80 65.7697
R34076 VCC.n9852 VCC.t90 65.7697
R34077 VCC.n10409 VCC.t67 65.7697
R34078 VCC.n10959 VCC.t78 65.7697
R34079 VCC.n11516 VCC.t415 65.7697
R34080 VCC.n12066 VCC.t545 65.7697
R34081 VCC.n12623 VCC.t359 65.7697
R34082 VCC.n13173 VCC.t70 65.7697
R34083 VCC.n13730 VCC.t294 65.7697
R34084 VCC.n14280 VCC.t311 65.7697
R34085 VCC.n14837 VCC.t283 65.7697
R34086 VCC.n15387 VCC.t455 65.7697
R34087 VCC.n15944 VCC.t144 65.7697
R34088 VCC.n16494 VCC.t245 65.7697
R34089 VCC.n17051 VCC.t45 65.7697
R34090 VCC.n17414 VCC.t578 65.7697
R34091 VCC.n293 VCC.n292 50.4194
R34092 VCC.n845 VCC.n844 50.4194
R34093 VCC.n1403 VCC.n1402 50.4194
R34094 VCC.n1954 VCC.n1953 50.4194
R34095 VCC.n2512 VCC.n2511 50.4194
R34096 VCC.n3063 VCC.n3062 50.4194
R34097 VCC.n3621 VCC.n3620 50.4194
R34098 VCC.n4172 VCC.n4171 50.4194
R34099 VCC.n4730 VCC.n4729 50.4194
R34100 VCC.n5281 VCC.n5280 50.4194
R34101 VCC.n5839 VCC.n5838 50.4194
R34102 VCC.n6390 VCC.n6389 50.4194
R34103 VCC.n6948 VCC.n6947 50.4194
R34104 VCC.n7499 VCC.n7498 50.4194
R34105 VCC.n8057 VCC.n8056 50.4194
R34106 VCC.n8608 VCC.n8607 50.4194
R34107 VCC.n9166 VCC.n9165 50.4194
R34108 VCC.n9717 VCC.n9716 50.4194
R34109 VCC.n10274 VCC.n10273 50.4194
R34110 VCC.n10824 VCC.n10823 50.4194
R34111 VCC.n11381 VCC.n11380 50.4194
R34112 VCC.n11931 VCC.n11930 50.4194
R34113 VCC.n12488 VCC.n12487 50.4194
R34114 VCC.n13038 VCC.n13037 50.4194
R34115 VCC.n13595 VCC.n13594 50.4194
R34116 VCC.n14145 VCC.n14144 50.4194
R34117 VCC.n14702 VCC.n14701 50.4194
R34118 VCC.n15252 VCC.n15251 50.4194
R34119 VCC.n15809 VCC.n15808 50.4194
R34120 VCC.n16359 VCC.n16358 50.4194
R34121 VCC.n16916 VCC.n16915 50.4194
R34122 VCC.n212 VCC.n182 50.3505
R34123 VCC.n230 VCC.n179 50.3505
R34124 VCC.n288 VCC.n143 50.3505
R34125 VCC.n334 VCC.n119 50.3505
R34126 VCC.n359 VCC.n109 50.3505
R34127 VCC.n397 VCC.n83 50.3505
R34128 VCC.n429 VCC.n80 50.3505
R34129 VCC.n764 VCC.n734 50.3505
R34130 VCC.n782 VCC.n731 50.3505
R34131 VCC.n840 VCC.n695 50.3505
R34132 VCC.n886 VCC.n671 50.3505
R34133 VCC.n911 VCC.n661 50.3505
R34134 VCC.n949 VCC.n635 50.3505
R34135 VCC.n981 VCC.n632 50.3505
R34136 VCC.n1443 VCC.n1228 50.3505
R34137 VCC.n1468 VCC.n1218 50.3505
R34138 VCC.n1506 VCC.n1192 50.3505
R34139 VCC.n1539 VCC.n1189 50.3505
R34140 VCC.n1322 VCC.n1292 50.3505
R34141 VCC.n1340 VCC.n1289 50.3505
R34142 VCC.n1398 VCC.n1253 50.3505
R34143 VCC.n1873 VCC.n1843 50.3505
R34144 VCC.n1891 VCC.n1840 50.3505
R34145 VCC.n1949 VCC.n1804 50.3505
R34146 VCC.n1995 VCC.n1780 50.3505
R34147 VCC.n2020 VCC.n1770 50.3505
R34148 VCC.n2058 VCC.n1744 50.3505
R34149 VCC.n2090 VCC.n1741 50.3505
R34150 VCC.n2552 VCC.n2337 50.3505
R34151 VCC.n2577 VCC.n2327 50.3505
R34152 VCC.n2615 VCC.n2301 50.3505
R34153 VCC.n2648 VCC.n2298 50.3505
R34154 VCC.n2431 VCC.n2401 50.3505
R34155 VCC.n2449 VCC.n2398 50.3505
R34156 VCC.n2507 VCC.n2362 50.3505
R34157 VCC.n2982 VCC.n2952 50.3505
R34158 VCC.n3000 VCC.n2949 50.3505
R34159 VCC.n3058 VCC.n2913 50.3505
R34160 VCC.n3104 VCC.n2889 50.3505
R34161 VCC.n3129 VCC.n2879 50.3505
R34162 VCC.n3167 VCC.n2853 50.3505
R34163 VCC.n3199 VCC.n2850 50.3505
R34164 VCC.n3661 VCC.n3446 50.3505
R34165 VCC.n3686 VCC.n3436 50.3505
R34166 VCC.n3724 VCC.n3410 50.3505
R34167 VCC.n3757 VCC.n3407 50.3505
R34168 VCC.n3540 VCC.n3510 50.3505
R34169 VCC.n3558 VCC.n3507 50.3505
R34170 VCC.n3616 VCC.n3471 50.3505
R34171 VCC.n4091 VCC.n4061 50.3505
R34172 VCC.n4109 VCC.n4058 50.3505
R34173 VCC.n4167 VCC.n4022 50.3505
R34174 VCC.n4213 VCC.n3998 50.3505
R34175 VCC.n4238 VCC.n3988 50.3505
R34176 VCC.n4276 VCC.n3962 50.3505
R34177 VCC.n4308 VCC.n3959 50.3505
R34178 VCC.n4770 VCC.n4555 50.3505
R34179 VCC.n4795 VCC.n4545 50.3505
R34180 VCC.n4833 VCC.n4519 50.3505
R34181 VCC.n4866 VCC.n4516 50.3505
R34182 VCC.n4649 VCC.n4619 50.3505
R34183 VCC.n4667 VCC.n4616 50.3505
R34184 VCC.n4725 VCC.n4580 50.3505
R34185 VCC.n5200 VCC.n5170 50.3505
R34186 VCC.n5218 VCC.n5167 50.3505
R34187 VCC.n5276 VCC.n5131 50.3505
R34188 VCC.n5322 VCC.n5107 50.3505
R34189 VCC.n5347 VCC.n5097 50.3505
R34190 VCC.n5385 VCC.n5071 50.3505
R34191 VCC.n5417 VCC.n5068 50.3505
R34192 VCC.n5879 VCC.n5664 50.3505
R34193 VCC.n5904 VCC.n5654 50.3505
R34194 VCC.n5942 VCC.n5628 50.3505
R34195 VCC.n5975 VCC.n5625 50.3505
R34196 VCC.n5758 VCC.n5728 50.3505
R34197 VCC.n5776 VCC.n5725 50.3505
R34198 VCC.n5834 VCC.n5689 50.3505
R34199 VCC.n6309 VCC.n6279 50.3505
R34200 VCC.n6327 VCC.n6276 50.3505
R34201 VCC.n6385 VCC.n6240 50.3505
R34202 VCC.n6431 VCC.n6216 50.3505
R34203 VCC.n6456 VCC.n6206 50.3505
R34204 VCC.n6494 VCC.n6180 50.3505
R34205 VCC.n6526 VCC.n6177 50.3505
R34206 VCC.n6988 VCC.n6773 50.3505
R34207 VCC.n7013 VCC.n6763 50.3505
R34208 VCC.n7051 VCC.n6737 50.3505
R34209 VCC.n7084 VCC.n6734 50.3505
R34210 VCC.n6867 VCC.n6837 50.3505
R34211 VCC.n6885 VCC.n6834 50.3505
R34212 VCC.n6943 VCC.n6798 50.3505
R34213 VCC.n7418 VCC.n7388 50.3505
R34214 VCC.n7436 VCC.n7385 50.3505
R34215 VCC.n7494 VCC.n7349 50.3505
R34216 VCC.n7540 VCC.n7325 50.3505
R34217 VCC.n7565 VCC.n7315 50.3505
R34218 VCC.n7603 VCC.n7289 50.3505
R34219 VCC.n7635 VCC.n7286 50.3505
R34220 VCC.n8097 VCC.n7882 50.3505
R34221 VCC.n8122 VCC.n7872 50.3505
R34222 VCC.n8160 VCC.n7846 50.3505
R34223 VCC.n8193 VCC.n7843 50.3505
R34224 VCC.n7976 VCC.n7946 50.3505
R34225 VCC.n7994 VCC.n7943 50.3505
R34226 VCC.n8052 VCC.n7907 50.3505
R34227 VCC.n8649 VCC.n8434 50.3505
R34228 VCC.n8674 VCC.n8424 50.3505
R34229 VCC.n8712 VCC.n8398 50.3505
R34230 VCC.n8744 VCC.n8395 50.3505
R34231 VCC.n8527 VCC.n8497 50.3505
R34232 VCC.n8545 VCC.n8494 50.3505
R34233 VCC.n8603 VCC.n8458 50.3505
R34234 VCC.n9206 VCC.n8991 50.3505
R34235 VCC.n9231 VCC.n8981 50.3505
R34236 VCC.n9269 VCC.n8955 50.3505
R34237 VCC.n9302 VCC.n8952 50.3505
R34238 VCC.n9085 VCC.n9055 50.3505
R34239 VCC.n9103 VCC.n9052 50.3505
R34240 VCC.n9161 VCC.n9016 50.3505
R34241 VCC.n9636 VCC.n9606 50.3505
R34242 VCC.n9654 VCC.n9603 50.3505
R34243 VCC.n9712 VCC.n9567 50.3505
R34244 VCC.n9758 VCC.n9543 50.3505
R34245 VCC.n9783 VCC.n9533 50.3505
R34246 VCC.n9821 VCC.n9507 50.3505
R34247 VCC.n9853 VCC.n9504 50.3505
R34248 VCC.n10314 VCC.n10099 50.3505
R34249 VCC.n10339 VCC.n10089 50.3505
R34250 VCC.n10377 VCC.n10063 50.3505
R34251 VCC.n10410 VCC.n10060 50.3505
R34252 VCC.n10193 VCC.n10163 50.3505
R34253 VCC.n10211 VCC.n10160 50.3505
R34254 VCC.n10269 VCC.n10124 50.3505
R34255 VCC.n10743 VCC.n10713 50.3505
R34256 VCC.n10761 VCC.n10710 50.3505
R34257 VCC.n10819 VCC.n10674 50.3505
R34258 VCC.n10865 VCC.n10650 50.3505
R34259 VCC.n10890 VCC.n10640 50.3505
R34260 VCC.n10928 VCC.n10614 50.3505
R34261 VCC.n10960 VCC.n10611 50.3505
R34262 VCC.n11421 VCC.n11206 50.3505
R34263 VCC.n11446 VCC.n11196 50.3505
R34264 VCC.n11484 VCC.n11170 50.3505
R34265 VCC.n11517 VCC.n11167 50.3505
R34266 VCC.n11300 VCC.n11270 50.3505
R34267 VCC.n11318 VCC.n11267 50.3505
R34268 VCC.n11376 VCC.n11231 50.3505
R34269 VCC.n11850 VCC.n11820 50.3505
R34270 VCC.n11868 VCC.n11817 50.3505
R34271 VCC.n11926 VCC.n11781 50.3505
R34272 VCC.n11972 VCC.n11757 50.3505
R34273 VCC.n11997 VCC.n11747 50.3505
R34274 VCC.n12035 VCC.n11721 50.3505
R34275 VCC.n12067 VCC.n11718 50.3505
R34276 VCC.n12528 VCC.n12313 50.3505
R34277 VCC.n12553 VCC.n12303 50.3505
R34278 VCC.n12591 VCC.n12277 50.3505
R34279 VCC.n12624 VCC.n12274 50.3505
R34280 VCC.n12407 VCC.n12377 50.3505
R34281 VCC.n12425 VCC.n12374 50.3505
R34282 VCC.n12483 VCC.n12338 50.3505
R34283 VCC.n12957 VCC.n12927 50.3505
R34284 VCC.n12975 VCC.n12924 50.3505
R34285 VCC.n13033 VCC.n12888 50.3505
R34286 VCC.n13079 VCC.n12864 50.3505
R34287 VCC.n13104 VCC.n12854 50.3505
R34288 VCC.n13142 VCC.n12828 50.3505
R34289 VCC.n13174 VCC.n12825 50.3505
R34290 VCC.n13635 VCC.n13420 50.3505
R34291 VCC.n13660 VCC.n13410 50.3505
R34292 VCC.n13698 VCC.n13384 50.3505
R34293 VCC.n13731 VCC.n13381 50.3505
R34294 VCC.n13514 VCC.n13484 50.3505
R34295 VCC.n13532 VCC.n13481 50.3505
R34296 VCC.n13590 VCC.n13445 50.3505
R34297 VCC.n14064 VCC.n14034 50.3505
R34298 VCC.n14082 VCC.n14031 50.3505
R34299 VCC.n14140 VCC.n13995 50.3505
R34300 VCC.n14186 VCC.n13971 50.3505
R34301 VCC.n14211 VCC.n13961 50.3505
R34302 VCC.n14249 VCC.n13935 50.3505
R34303 VCC.n14281 VCC.n13932 50.3505
R34304 VCC.n14742 VCC.n14527 50.3505
R34305 VCC.n14767 VCC.n14517 50.3505
R34306 VCC.n14805 VCC.n14491 50.3505
R34307 VCC.n14838 VCC.n14488 50.3505
R34308 VCC.n14621 VCC.n14591 50.3505
R34309 VCC.n14639 VCC.n14588 50.3505
R34310 VCC.n14697 VCC.n14552 50.3505
R34311 VCC.n15171 VCC.n15141 50.3505
R34312 VCC.n15189 VCC.n15138 50.3505
R34313 VCC.n15247 VCC.n15102 50.3505
R34314 VCC.n15293 VCC.n15078 50.3505
R34315 VCC.n15318 VCC.n15068 50.3505
R34316 VCC.n15356 VCC.n15042 50.3505
R34317 VCC.n15388 VCC.n15039 50.3505
R34318 VCC.n15849 VCC.n15634 50.3505
R34319 VCC.n15874 VCC.n15624 50.3505
R34320 VCC.n15912 VCC.n15598 50.3505
R34321 VCC.n15945 VCC.n15595 50.3505
R34322 VCC.n15728 VCC.n15698 50.3505
R34323 VCC.n15746 VCC.n15695 50.3505
R34324 VCC.n15804 VCC.n15659 50.3505
R34325 VCC.n16278 VCC.n16248 50.3505
R34326 VCC.n16296 VCC.n16245 50.3505
R34327 VCC.n16354 VCC.n16209 50.3505
R34328 VCC.n16400 VCC.n16185 50.3505
R34329 VCC.n16425 VCC.n16175 50.3505
R34330 VCC.n16463 VCC.n16149 50.3505
R34331 VCC.n16495 VCC.n16146 50.3505
R34332 VCC.n16956 VCC.n16741 50.3505
R34333 VCC.n16981 VCC.n16731 50.3505
R34334 VCC.n17019 VCC.n16705 50.3505
R34335 VCC.n17052 VCC.n16702 50.3505
R34336 VCC.n16835 VCC.n16805 50.3505
R34337 VCC.n16853 VCC.n16802 50.3505
R34338 VCC.n16911 VCC.n16766 50.3505
R34339 VCC.n17320 VCC.n17292 50.3505
R34340 VCC.n17345 VCC.n17282 50.3505
R34341 VCC.n17383 VCC.n17256 50.3505
R34342 VCC.n17415 VCC.n17253 50.3505
R34343 VCC.n265 VCC.n154 49.4005
R34344 VCC.n265 VCC.n152 49.4005
R34345 VCC.n363 VCC.n94 49.4005
R34346 VCC.n393 VCC.n94 49.4005
R34347 VCC.n817 VCC.n706 49.4005
R34348 VCC.n817 VCC.n704 49.4005
R34349 VCC.n915 VCC.n646 49.4005
R34350 VCC.n945 VCC.n646 49.4005
R34351 VCC.n1472 VCC.n1203 49.4005
R34352 VCC.n1502 VCC.n1203 49.4005
R34353 VCC.n1375 VCC.n1264 49.4005
R34354 VCC.n1375 VCC.n1262 49.4005
R34355 VCC.n1926 VCC.n1815 49.4005
R34356 VCC.n1926 VCC.n1813 49.4005
R34357 VCC.n2024 VCC.n1755 49.4005
R34358 VCC.n2054 VCC.n1755 49.4005
R34359 VCC.n2581 VCC.n2312 49.4005
R34360 VCC.n2611 VCC.n2312 49.4005
R34361 VCC.n2484 VCC.n2373 49.4005
R34362 VCC.n2484 VCC.n2371 49.4005
R34363 VCC.n3035 VCC.n2924 49.4005
R34364 VCC.n3035 VCC.n2922 49.4005
R34365 VCC.n3133 VCC.n2864 49.4005
R34366 VCC.n3163 VCC.n2864 49.4005
R34367 VCC.n3690 VCC.n3421 49.4005
R34368 VCC.n3720 VCC.n3421 49.4005
R34369 VCC.n3593 VCC.n3482 49.4005
R34370 VCC.n3593 VCC.n3480 49.4005
R34371 VCC.n4144 VCC.n4033 49.4005
R34372 VCC.n4144 VCC.n4031 49.4005
R34373 VCC.n4242 VCC.n3973 49.4005
R34374 VCC.n4272 VCC.n3973 49.4005
R34375 VCC.n4799 VCC.n4530 49.4005
R34376 VCC.n4829 VCC.n4530 49.4005
R34377 VCC.n4702 VCC.n4591 49.4005
R34378 VCC.n4702 VCC.n4589 49.4005
R34379 VCC.n5253 VCC.n5142 49.4005
R34380 VCC.n5253 VCC.n5140 49.4005
R34381 VCC.n5351 VCC.n5082 49.4005
R34382 VCC.n5381 VCC.n5082 49.4005
R34383 VCC.n5908 VCC.n5639 49.4005
R34384 VCC.n5938 VCC.n5639 49.4005
R34385 VCC.n5811 VCC.n5700 49.4005
R34386 VCC.n5811 VCC.n5698 49.4005
R34387 VCC.n6362 VCC.n6251 49.4005
R34388 VCC.n6362 VCC.n6249 49.4005
R34389 VCC.n6460 VCC.n6191 49.4005
R34390 VCC.n6490 VCC.n6191 49.4005
R34391 VCC.n7017 VCC.n6748 49.4005
R34392 VCC.n7047 VCC.n6748 49.4005
R34393 VCC.n6920 VCC.n6809 49.4005
R34394 VCC.n6920 VCC.n6807 49.4005
R34395 VCC.n7471 VCC.n7360 49.4005
R34396 VCC.n7471 VCC.n7358 49.4005
R34397 VCC.n7569 VCC.n7300 49.4005
R34398 VCC.n7599 VCC.n7300 49.4005
R34399 VCC.n8126 VCC.n7857 49.4005
R34400 VCC.n8156 VCC.n7857 49.4005
R34401 VCC.n8029 VCC.n7918 49.4005
R34402 VCC.n8029 VCC.n7916 49.4005
R34403 VCC.n8678 VCC.n8409 49.4005
R34404 VCC.n8708 VCC.n8409 49.4005
R34405 VCC.n8580 VCC.n8469 49.4005
R34406 VCC.n8580 VCC.n8467 49.4005
R34407 VCC.n9235 VCC.n8966 49.4005
R34408 VCC.n9265 VCC.n8966 49.4005
R34409 VCC.n9138 VCC.n9027 49.4005
R34410 VCC.n9138 VCC.n9025 49.4005
R34411 VCC.n9689 VCC.n9578 49.4005
R34412 VCC.n9689 VCC.n9576 49.4005
R34413 VCC.n9787 VCC.n9518 49.4005
R34414 VCC.n9817 VCC.n9518 49.4005
R34415 VCC.n10343 VCC.n10074 49.4005
R34416 VCC.n10373 VCC.n10074 49.4005
R34417 VCC.n10246 VCC.n10135 49.4005
R34418 VCC.n10246 VCC.n10133 49.4005
R34419 VCC.n10796 VCC.n10685 49.4005
R34420 VCC.n10796 VCC.n10683 49.4005
R34421 VCC.n10894 VCC.n10625 49.4005
R34422 VCC.n10924 VCC.n10625 49.4005
R34423 VCC.n11450 VCC.n11181 49.4005
R34424 VCC.n11480 VCC.n11181 49.4005
R34425 VCC.n11353 VCC.n11242 49.4005
R34426 VCC.n11353 VCC.n11240 49.4005
R34427 VCC.n11903 VCC.n11792 49.4005
R34428 VCC.n11903 VCC.n11790 49.4005
R34429 VCC.n12001 VCC.n11732 49.4005
R34430 VCC.n12031 VCC.n11732 49.4005
R34431 VCC.n12557 VCC.n12288 49.4005
R34432 VCC.n12587 VCC.n12288 49.4005
R34433 VCC.n12460 VCC.n12349 49.4005
R34434 VCC.n12460 VCC.n12347 49.4005
R34435 VCC.n13010 VCC.n12899 49.4005
R34436 VCC.n13010 VCC.n12897 49.4005
R34437 VCC.n13108 VCC.n12839 49.4005
R34438 VCC.n13138 VCC.n12839 49.4005
R34439 VCC.n13664 VCC.n13395 49.4005
R34440 VCC.n13694 VCC.n13395 49.4005
R34441 VCC.n13567 VCC.n13456 49.4005
R34442 VCC.n13567 VCC.n13454 49.4005
R34443 VCC.n14117 VCC.n14006 49.4005
R34444 VCC.n14117 VCC.n14004 49.4005
R34445 VCC.n14215 VCC.n13946 49.4005
R34446 VCC.n14245 VCC.n13946 49.4005
R34447 VCC.n14771 VCC.n14502 49.4005
R34448 VCC.n14801 VCC.n14502 49.4005
R34449 VCC.n14674 VCC.n14563 49.4005
R34450 VCC.n14674 VCC.n14561 49.4005
R34451 VCC.n15224 VCC.n15113 49.4005
R34452 VCC.n15224 VCC.n15111 49.4005
R34453 VCC.n15322 VCC.n15053 49.4005
R34454 VCC.n15352 VCC.n15053 49.4005
R34455 VCC.n15878 VCC.n15609 49.4005
R34456 VCC.n15908 VCC.n15609 49.4005
R34457 VCC.n15781 VCC.n15670 49.4005
R34458 VCC.n15781 VCC.n15668 49.4005
R34459 VCC.n16331 VCC.n16220 49.4005
R34460 VCC.n16331 VCC.n16218 49.4005
R34461 VCC.n16429 VCC.n16160 49.4005
R34462 VCC.n16459 VCC.n16160 49.4005
R34463 VCC.n16985 VCC.n16716 49.4005
R34464 VCC.n17015 VCC.n16716 49.4005
R34465 VCC.n16888 VCC.n16777 49.4005
R34466 VCC.n16888 VCC.n16775 49.4005
R34467 VCC.n17349 VCC.n17267 49.4005
R34468 VCC.n17379 VCC.n17267 49.4005
R34469 VCC.n469 VCC.n56 43.1576
R34470 VCC.n474 VCC.n42 43.1576
R34471 VCC.n493 VCC.n40 43.1576
R34472 VCC.n497 VCC.n40 43.1576
R34473 VCC.n524 VCC.n21 43.1576
R34474 VCC.n546 VCC.n6 43.1576
R34475 VCC.n1021 VCC.n608 43.1576
R34476 VCC.n1026 VCC.n594 43.1576
R34477 VCC.n1045 VCC.n592 43.1576
R34478 VCC.n1049 VCC.n592 43.1576
R34479 VCC.n1076 VCC.n573 43.1576
R34480 VCC.n1100 VCC.n560 43.1576
R34481 VCC.n1530 VCC.n1164 43.1576
R34482 VCC.n1586 VCC.n1161 43.1576
R34483 VCC.n1582 VCC.n1144 43.1576
R34484 VCC.n1618 VCC.n1144 43.1576
R34485 VCC.n1622 VCC.n1115 43.1576
R34486 VCC.n1654 VCC.n1113 43.1576
R34487 VCC.n2130 VCC.n1717 43.1576
R34488 VCC.n2135 VCC.n1703 43.1576
R34489 VCC.n2154 VCC.n1701 43.1576
R34490 VCC.n2158 VCC.n1701 43.1576
R34491 VCC.n2185 VCC.n1682 43.1576
R34492 VCC.n2209 VCC.n1669 43.1576
R34493 VCC.n2639 VCC.n2273 43.1576
R34494 VCC.n2695 VCC.n2270 43.1576
R34495 VCC.n2691 VCC.n2253 43.1576
R34496 VCC.n2727 VCC.n2253 43.1576
R34497 VCC.n2731 VCC.n2224 43.1576
R34498 VCC.n2763 VCC.n2222 43.1576
R34499 VCC.n3239 VCC.n2826 43.1576
R34500 VCC.n3244 VCC.n2812 43.1576
R34501 VCC.n3263 VCC.n2810 43.1576
R34502 VCC.n3267 VCC.n2810 43.1576
R34503 VCC.n3294 VCC.n2791 43.1576
R34504 VCC.n3318 VCC.n2778 43.1576
R34505 VCC.n3748 VCC.n3382 43.1576
R34506 VCC.n3804 VCC.n3379 43.1576
R34507 VCC.n3800 VCC.n3362 43.1576
R34508 VCC.n3836 VCC.n3362 43.1576
R34509 VCC.n3840 VCC.n3333 43.1576
R34510 VCC.n3872 VCC.n3331 43.1576
R34511 VCC.n4348 VCC.n3935 43.1576
R34512 VCC.n4353 VCC.n3921 43.1576
R34513 VCC.n4372 VCC.n3919 43.1576
R34514 VCC.n4376 VCC.n3919 43.1576
R34515 VCC.n4403 VCC.n3900 43.1576
R34516 VCC.n4427 VCC.n3887 43.1576
R34517 VCC.n4857 VCC.n4491 43.1576
R34518 VCC.n4913 VCC.n4488 43.1576
R34519 VCC.n4909 VCC.n4471 43.1576
R34520 VCC.n4945 VCC.n4471 43.1576
R34521 VCC.n4949 VCC.n4442 43.1576
R34522 VCC.n4981 VCC.n4440 43.1576
R34523 VCC.n5457 VCC.n5044 43.1576
R34524 VCC.n5462 VCC.n5030 43.1576
R34525 VCC.n5481 VCC.n5028 43.1576
R34526 VCC.n5485 VCC.n5028 43.1576
R34527 VCC.n5512 VCC.n5009 43.1576
R34528 VCC.n5536 VCC.n4996 43.1576
R34529 VCC.n5966 VCC.n5600 43.1576
R34530 VCC.n6022 VCC.n5597 43.1576
R34531 VCC.n6018 VCC.n5580 43.1576
R34532 VCC.n6054 VCC.n5580 43.1576
R34533 VCC.n6058 VCC.n5551 43.1576
R34534 VCC.n6090 VCC.n5549 43.1576
R34535 VCC.n6566 VCC.n6153 43.1576
R34536 VCC.n6571 VCC.n6139 43.1576
R34537 VCC.n6590 VCC.n6137 43.1576
R34538 VCC.n6594 VCC.n6137 43.1576
R34539 VCC.n6621 VCC.n6118 43.1576
R34540 VCC.n6645 VCC.n6105 43.1576
R34541 VCC.n7075 VCC.n6709 43.1576
R34542 VCC.n7131 VCC.n6706 43.1576
R34543 VCC.n7127 VCC.n6689 43.1576
R34544 VCC.n7163 VCC.n6689 43.1576
R34545 VCC.n7167 VCC.n6660 43.1576
R34546 VCC.n7199 VCC.n6658 43.1576
R34547 VCC.n7675 VCC.n7262 43.1576
R34548 VCC.n7680 VCC.n7248 43.1576
R34549 VCC.n7699 VCC.n7246 43.1576
R34550 VCC.n7703 VCC.n7246 43.1576
R34551 VCC.n7730 VCC.n7227 43.1576
R34552 VCC.n7754 VCC.n7214 43.1576
R34553 VCC.n8184 VCC.n7818 43.1576
R34554 VCC.n8240 VCC.n7815 43.1576
R34555 VCC.n8236 VCC.n7798 43.1576
R34556 VCC.n8272 VCC.n7798 43.1576
R34557 VCC.n8276 VCC.n7769 43.1576
R34558 VCC.n8308 VCC.n7767 43.1576
R34559 VCC.n8784 VCC.n8371 43.1576
R34560 VCC.n8789 VCC.n8357 43.1576
R34561 VCC.n8808 VCC.n8355 43.1576
R34562 VCC.n8812 VCC.n8355 43.1576
R34563 VCC.n8839 VCC.n8336 43.1576
R34564 VCC.n8863 VCC.n8323 43.1576
R34565 VCC.n9293 VCC.n8927 43.1576
R34566 VCC.n9349 VCC.n8924 43.1576
R34567 VCC.n9345 VCC.n8907 43.1576
R34568 VCC.n9381 VCC.n8907 43.1576
R34569 VCC.n9385 VCC.n8878 43.1576
R34570 VCC.n9417 VCC.n8876 43.1576
R34571 VCC.n9893 VCC.n9480 43.1576
R34572 VCC.n9898 VCC.n9466 43.1576
R34573 VCC.n9917 VCC.n9464 43.1576
R34574 VCC.n9921 VCC.n9464 43.1576
R34575 VCC.n9948 VCC.n9445 43.1576
R34576 VCC.n9972 VCC.n9432 43.1576
R34577 VCC.n10401 VCC.n10035 43.1576
R34578 VCC.n10457 VCC.n10032 43.1576
R34579 VCC.n10453 VCC.n10015 43.1576
R34580 VCC.n10489 VCC.n10015 43.1576
R34581 VCC.n10493 VCC.n9986 43.1576
R34582 VCC.n10525 VCC.n9984 43.1576
R34583 VCC.n11000 VCC.n10587 43.1576
R34584 VCC.n11005 VCC.n10573 43.1576
R34585 VCC.n11024 VCC.n10571 43.1576
R34586 VCC.n11028 VCC.n10571 43.1576
R34587 VCC.n11055 VCC.n10552 43.1576
R34588 VCC.n11079 VCC.n10539 43.1576
R34589 VCC.n11508 VCC.n11142 43.1576
R34590 VCC.n11564 VCC.n11139 43.1576
R34591 VCC.n11560 VCC.n11122 43.1576
R34592 VCC.n11596 VCC.n11122 43.1576
R34593 VCC.n11600 VCC.n11093 43.1576
R34594 VCC.n11632 VCC.n11091 43.1576
R34595 VCC.n12107 VCC.n11694 43.1576
R34596 VCC.n12112 VCC.n11680 43.1576
R34597 VCC.n12131 VCC.n11678 43.1576
R34598 VCC.n12135 VCC.n11678 43.1576
R34599 VCC.n12162 VCC.n11659 43.1576
R34600 VCC.n12186 VCC.n11646 43.1576
R34601 VCC.n12615 VCC.n12249 43.1576
R34602 VCC.n12671 VCC.n12246 43.1576
R34603 VCC.n12667 VCC.n12229 43.1576
R34604 VCC.n12703 VCC.n12229 43.1576
R34605 VCC.n12707 VCC.n12200 43.1576
R34606 VCC.n12739 VCC.n12198 43.1576
R34607 VCC.n13214 VCC.n12801 43.1576
R34608 VCC.n13219 VCC.n12787 43.1576
R34609 VCC.n13238 VCC.n12785 43.1576
R34610 VCC.n13242 VCC.n12785 43.1576
R34611 VCC.n13269 VCC.n12766 43.1576
R34612 VCC.n13293 VCC.n12753 43.1576
R34613 VCC.n13722 VCC.n13356 43.1576
R34614 VCC.n13778 VCC.n13353 43.1576
R34615 VCC.n13774 VCC.n13336 43.1576
R34616 VCC.n13810 VCC.n13336 43.1576
R34617 VCC.n13814 VCC.n13307 43.1576
R34618 VCC.n13846 VCC.n13305 43.1576
R34619 VCC.n14321 VCC.n13908 43.1576
R34620 VCC.n14326 VCC.n13894 43.1576
R34621 VCC.n14345 VCC.n13892 43.1576
R34622 VCC.n14349 VCC.n13892 43.1576
R34623 VCC.n14376 VCC.n13873 43.1576
R34624 VCC.n14400 VCC.n13860 43.1576
R34625 VCC.n14829 VCC.n14463 43.1576
R34626 VCC.n14885 VCC.n14460 43.1576
R34627 VCC.n14881 VCC.n14443 43.1576
R34628 VCC.n14917 VCC.n14443 43.1576
R34629 VCC.n14921 VCC.n14414 43.1576
R34630 VCC.n14953 VCC.n14412 43.1576
R34631 VCC.n15428 VCC.n15015 43.1576
R34632 VCC.n15433 VCC.n15001 43.1576
R34633 VCC.n15452 VCC.n14999 43.1576
R34634 VCC.n15456 VCC.n14999 43.1576
R34635 VCC.n15483 VCC.n14980 43.1576
R34636 VCC.n15507 VCC.n14967 43.1576
R34637 VCC.n15936 VCC.n15570 43.1576
R34638 VCC.n15992 VCC.n15567 43.1576
R34639 VCC.n15988 VCC.n15550 43.1576
R34640 VCC.n16024 VCC.n15550 43.1576
R34641 VCC.n16028 VCC.n15521 43.1576
R34642 VCC.n16060 VCC.n15519 43.1576
R34643 VCC.n16535 VCC.n16122 43.1576
R34644 VCC.n16540 VCC.n16108 43.1576
R34645 VCC.n16559 VCC.n16106 43.1576
R34646 VCC.n16563 VCC.n16106 43.1576
R34647 VCC.n16590 VCC.n16087 43.1576
R34648 VCC.n16614 VCC.n16074 43.1576
R34649 VCC.n17043 VCC.n16677 43.1576
R34650 VCC.n17099 VCC.n16674 43.1576
R34651 VCC.n17095 VCC.n16657 43.1576
R34652 VCC.n17131 VCC.n16657 43.1576
R34653 VCC.n17135 VCC.n16628 43.1576
R34654 VCC.n17167 VCC.n16626 43.1576
R34655 VCC.n17455 VCC.n17229 43.1576
R34656 VCC.n17460 VCC.n17215 43.1576
R34657 VCC.n17479 VCC.n17213 43.1576
R34658 VCC.n17483 VCC.n17213 43.1576
R34659 VCC.n17510 VCC.n17194 43.1576
R34660 VCC.n17534 VCC.n17181 43.1576
R34661 VCC.n548 VCC.n547 36.8662
R34662 VCC.n1102 VCC.n1101 36.8662
R34663 VCC.n1653 VCC.n1111 36.8662
R34664 VCC.n2211 VCC.n2210 36.8662
R34665 VCC.n2762 VCC.n2220 36.8662
R34666 VCC.n3320 VCC.n3319 36.8662
R34667 VCC.n3871 VCC.n3329 36.8662
R34668 VCC.n4429 VCC.n4428 36.8662
R34669 VCC.n4980 VCC.n4438 36.8662
R34670 VCC.n5538 VCC.n5537 36.8662
R34671 VCC.n6089 VCC.n5547 36.8662
R34672 VCC.n6647 VCC.n6646 36.8662
R34673 VCC.n7198 VCC.n6656 36.8662
R34674 VCC.n7756 VCC.n7755 36.8662
R34675 VCC.n8307 VCC.n7765 36.8662
R34676 VCC.n8865 VCC.n8864 36.8662
R34677 VCC.n9416 VCC.n8874 36.8662
R34678 VCC.n9974 VCC.n9973 36.8662
R34679 VCC.n10524 VCC.n9982 36.8662
R34680 VCC.n11081 VCC.n11080 36.8662
R34681 VCC.n11631 VCC.n11089 36.8662
R34682 VCC.n12188 VCC.n12187 36.8662
R34683 VCC.n12738 VCC.n12196 36.8662
R34684 VCC.n13295 VCC.n13294 36.8662
R34685 VCC.n13845 VCC.n13303 36.8662
R34686 VCC.n14402 VCC.n14401 36.8662
R34687 VCC.n14952 VCC.n14410 36.8662
R34688 VCC.n15509 VCC.n15508 36.8662
R34689 VCC.n16059 VCC.n15517 36.8662
R34690 VCC.n16616 VCC.n16615 36.8662
R34691 VCC.n17166 VCC.n16624 36.8662
R34692 VCC.n17536 VCC.n17535 36.8662
R34693 VCC.n446 VCC.t139 35.5869
R34694 VCC.n998 VCC.t129 35.5869
R34695 VCC.n1556 VCC.t65 35.5869
R34696 VCC.n2107 VCC.t385 35.5869
R34697 VCC.n2665 VCC.t410 35.5869
R34698 VCC.n3216 VCC.t183 35.5869
R34699 VCC.n3774 VCC.t522 35.5869
R34700 VCC.n4325 VCC.t164 35.5869
R34701 VCC.n4883 VCC.t43 35.5869
R34702 VCC.n5434 VCC.t171 35.5869
R34703 VCC.n5992 VCC.t222 35.5869
R34704 VCC.n6543 VCC.t242 35.5869
R34705 VCC.n7101 VCC.t393 35.5869
R34706 VCC.n7652 VCC.t516 35.5869
R34707 VCC.n8210 VCC.t99 35.5869
R34708 VCC.n8761 VCC.t62 35.5869
R34709 VCC.n9319 VCC.t81 35.5869
R34710 VCC.n9870 VCC.t91 35.5869
R34711 VCC.n10427 VCC.t68 35.5869
R34712 VCC.n10977 VCC.t79 35.5869
R34713 VCC.n11534 VCC.t416 35.5869
R34714 VCC.n12084 VCC.t546 35.5869
R34715 VCC.n12641 VCC.t360 35.5869
R34716 VCC.n13191 VCC.t71 35.5869
R34717 VCC.n13748 VCC.t295 35.5869
R34718 VCC.n14298 VCC.t312 35.5869
R34719 VCC.n14855 VCC.t284 35.5869
R34720 VCC.n15405 VCC.t456 35.5869
R34721 VCC.n15962 VCC.t145 35.5869
R34722 VCC.n16512 VCC.t246 35.5869
R34723 VCC.n17069 VCC.t46 35.5869
R34724 VCC.n17432 VCC.t579 35.5869
R34725 VCC.n11 VCC.t331 34.994
R34726 VCC.n1091 VCC.t186 34.994
R34727 VCC.n1640 VCC.t344 34.994
R34728 VCC.n2200 VCC.t435 34.994
R34729 VCC.n2749 VCC.t112 34.994
R34730 VCC.n3309 VCC.t373 34.994
R34731 VCC.n3858 VCC.t156 34.994
R34732 VCC.n4418 VCC.t39 34.994
R34733 VCC.n4967 VCC.t460 34.994
R34734 VCC.n5527 VCC.t1 34.994
R34735 VCC.n6076 VCC.t441 34.994
R34736 VCC.n6636 VCC.t257 34.994
R34737 VCC.n7185 VCC.t54 34.994
R34738 VCC.n7745 VCC.t169 34.994
R34739 VCC.n8294 VCC.t377 34.994
R34740 VCC.n8854 VCC.t447 34.994
R34741 VCC.n9403 VCC.t403 34.994
R34742 VCC.n9963 VCC.t495 34.994
R34743 VCC.n10511 VCC.t357 34.994
R34744 VCC.n11070 VCC.t32 34.994
R34745 VCC.n11618 VCC.t15 34.994
R34746 VCC.n12177 VCC.t502 34.994
R34747 VCC.n12725 VCC.t398 34.994
R34748 VCC.n13284 VCC.t268 34.994
R34749 VCC.n13832 VCC.t135 34.994
R34750 VCC.n14391 VCC.t572 34.994
R34751 VCC.n14939 VCC.t473 34.994
R34752 VCC.n15498 VCC.t508 34.994
R34753 VCC.n16046 VCC.t59 34.994
R34754 VCC.n16605 VCC.t175 34.994
R34755 VCC.n17153 VCC.t566 34.994
R34756 VCC.n17525 VCC.t625 34.994
R34757 VCC.n52 VCC.t190 34.9892
R34758 VCC.n604 VCC.t337 34.9892
R34759 VCC.n1157 VCC.t287 34.9892
R34760 VCC.n1713 VCC.t429 34.9892
R34761 VCC.n2266 VCC.t291 34.9892
R34762 VCC.n2822 VCC.t590 34.9892
R34763 VCC.n3375 VCC.t575 34.9892
R34764 VCC.n3931 VCC.t316 34.9892
R34765 VCC.n4484 VCC.t534 34.9892
R34766 VCC.n5040 VCC.t325 34.9892
R34767 VCC.n5593 VCC.t26 34.9892
R34768 VCC.n6149 VCC.t307 34.9892
R34769 VCC.n6702 VCC.t226 34.9892
R34770 VCC.n7258 VCC.t583 34.9892
R34771 VCC.n7811 VCC.t280 34.9892
R34772 VCC.n8367 VCC.t34 34.9892
R34773 VCC.n8920 VCC.t539 34.9892
R34774 VCC.n9476 VCC.t498 34.9892
R34775 VCC.n10028 VCC.t238 34.9892
R34776 VCC.n10583 VCC.t613 34.9892
R34777 VCC.n11135 VCC.t118 34.9892
R34778 VCC.n11690 VCC.t216 34.9892
R34779 VCC.n12242 VCC.t179 34.9892
R34780 VCC.n12797 VCC.t512 34.9892
R34781 VCC.n13349 VCC.t607 34.9892
R34782 VCC.n13904 VCC.t463 34.9892
R34783 VCC.n14456 VCC.t75 34.9892
R34784 VCC.n15011 VCC.t559 34.9892
R34785 VCC.n15563 VCC.t489 34.9892
R34786 VCC.n16118 VCC.t593 34.9892
R34787 VCC.n16670 VCC.t123 34.9892
R34788 VCC.n17225 VCC.t199 34.9892
R34789 VCC.n311 VCC.t11 34.9619
R34790 VCC.n863 VCC.t21 34.9619
R34791 VCC.n1421 VCC.t467 34.9619
R34792 VCC.n1972 VCC.t368 34.9619
R34793 VCC.n2530 VCC.t433 34.9619
R34794 VCC.n3081 VCC.t469 34.9619
R34795 VCC.n3639 VCC.t400 34.9619
R34796 VCC.n4190 VCC.t366 34.9619
R34797 VCC.n4748 VCC.t363 34.9619
R34798 VCC.n5299 VCC.t196 34.9619
R34799 VCC.n5857 VCC.t619 34.9619
R34800 VCC.n6408 VCC.t597 34.9619
R34801 VCC.n6966 VCC.t532 34.9619
R34802 VCC.n7517 VCC.t301 34.9619
R34803 VCC.n8075 VCC.t633 34.9619
R34804 VCC.n8626 VCC.t248 34.9619
R34805 VCC.n9184 VCC.t109 34.9619
R34806 VCC.n9735 VCC.t273 34.9619
R34807 VCC.n10292 VCC.t425 34.9619
R34808 VCC.n10842 VCC.t617 34.9619
R34809 VCC.n11399 VCC.t381 34.9619
R34810 VCC.n11949 VCC.t152 34.9619
R34811 VCC.n12506 VCC.t193 34.9619
R34812 VCC.n13056 VCC.t319 34.9619
R34813 VCC.n13613 VCC.t264 34.9619
R34814 VCC.n14163 VCC.t115 34.9619
R34815 VCC.n14720 VCC.t207 34.9619
R34816 VCC.n15270 VCC.t93 34.9619
R34817 VCC.n15827 VCC.t526 34.9619
R34818 VCC.n16377 VCC.t254 34.9619
R34819 VCC.n16934 VCC.t408 34.9619
R34820 VCC.n112 VCC.t568 34.945
R34821 VCC.n664 VCC.t391 34.945
R34822 VCC.n1221 VCC.t297 34.945
R34823 VCC.n1773 VCC.t554 34.945
R34824 VCC.n2330 VCC.t480 34.945
R34825 VCC.n2882 VCC.t328 34.945
R34826 VCC.n3439 VCC.t162 34.945
R34827 VCC.n3991 VCC.t159 34.945
R34828 VCC.n4548 VCC.t444 34.945
R34829 VCC.n5100 VCC.t102 34.945
R34830 VCC.n5657 VCC.t251 34.945
R34831 VCC.n6209 VCC.t149 34.945
R34832 VCC.n6766 VCC.t203 34.945
R34833 VCC.n7318 VCC.t97 34.945
R34834 VCC.n7875 VCC.t126 34.945
R34835 VCC.n8427 VCC.t476 34.945
R34836 VCC.n8984 VCC.t276 34.945
R34837 VCC.n9536 VCC.t483 34.945
R34838 VCC.n10092 VCC.t543 34.945
R34839 VCC.n10643 VCC.t220 34.945
R34840 VCC.n11199 VCC.t453 34.945
R34841 VCC.n11750 VCC.t88 34.945
R34842 VCC.n12306 VCC.t548 34.945
R34843 VCC.n12857 VCC.t213 34.945
R34844 VCC.n13413 VCC.t310 34.945
R34845 VCC.n13964 VCC.t587 34.945
R34846 VCC.n14520 VCC.t132 34.945
R34847 VCC.n15071 VCC.t341 34.945
R34848 VCC.n15627 VCC.t9 34.945
R34849 VCC.n16178 VCC.t519 34.945
R34850 VCC.n16734 VCC.t348 34.945
R34851 VCC.n17285 VCC.t370 34.945
R34852 VCC.n237 VCC.t233 34.9423
R34853 VCC.n789 VCC.t388 34.9423
R34854 VCC.n1347 VCC.t486 34.9423
R34855 VCC.n1898 VCC.t19 34.9423
R34856 VCC.n2456 VCC.t142 34.9423
R34857 VCC.n3007 VCC.t600 34.9423
R34858 VCC.n3565 VCC.t5 34.9423
R34859 VCC.n4116 VCC.t552 34.9423
R34860 VCC.n4674 VCC.t413 34.9423
R34861 VCC.n5225 VCC.t351 34.9423
R34862 VCC.n5783 VCC.t622 34.9423
R34863 VCC.n6334 VCC.t333 34.9423
R34864 VCC.n6892 VCC.t236 34.9423
R34865 VCC.n7443 VCC.t602 34.9423
R34866 VCC.n8001 VCC.t106 34.9423
R34867 VCC.n8552 VCC.t84 34.9423
R34868 VCC.n9110 VCC.t423 34.9423
R34869 VCC.n9661 VCC.t322 34.9423
R34870 VCC.n10218 VCC.t48 34.9423
R34871 VCC.n10768 VCC.t23 34.9423
R34872 VCC.n11325 VCC.t229 34.9423
R34873 VCC.n11875 VCC.t506 34.9423
R34874 VCC.n12432 VCC.t262 34.9423
R34875 VCC.n12982 VCC.t561 34.9423
R34876 VCC.n13539 VCC.t629 34.9423
R34877 VCC.n14089 VCC.t209 34.9423
R34878 VCC.n14646 VCC.t354 34.9423
R34879 VCC.n15196 VCC.t51 34.9423
R34880 VCC.n15753 VCC.t528 34.9423
R34881 VCC.n16303 VCC.t420 34.9423
R34882 VCC.n16860 VCC.t609 34.9423
R34883 VCC.n291 VCC.t10 32.8851
R34884 VCC.n843 VCC.t20 32.8851
R34885 VCC.n1401 VCC.t466 32.8851
R34886 VCC.n1952 VCC.t367 32.8851
R34887 VCC.n2510 VCC.t432 32.8851
R34888 VCC.n3061 VCC.t468 32.8851
R34889 VCC.n3619 VCC.t399 32.8851
R34890 VCC.n4170 VCC.t365 32.8851
R34891 VCC.n4728 VCC.t362 32.8851
R34892 VCC.n5279 VCC.t195 32.8851
R34893 VCC.n5837 VCC.t618 32.8851
R34894 VCC.n6388 VCC.t596 32.8851
R34895 VCC.n6946 VCC.t531 32.8851
R34896 VCC.n7497 VCC.t300 32.8851
R34897 VCC.n8055 VCC.t632 32.8851
R34898 VCC.n8606 VCC.t247 32.8851
R34899 VCC.n9164 VCC.t108 32.8851
R34900 VCC.n9715 VCC.t272 32.8851
R34901 VCC.n10272 VCC.t424 32.8851
R34902 VCC.n10822 VCC.t616 32.8851
R34903 VCC.n11379 VCC.t380 32.8851
R34904 VCC.n11929 VCC.t151 32.8851
R34905 VCC.n12486 VCC.t192 32.8851
R34906 VCC.n13036 VCC.t318 32.8851
R34907 VCC.n13593 VCC.t263 32.8851
R34908 VCC.n14143 VCC.t114 32.8851
R34909 VCC.n14700 VCC.t206 32.8851
R34910 VCC.n15250 VCC.t92 32.8851
R34911 VCC.n15807 VCC.t525 32.8851
R34912 VCC.n16357 VCC.t253 32.8851
R34913 VCC.n16914 VCC.t407 32.8851
R34914 VCC.t138 VCC.n418 31.0582
R34915 VCC.t128 VCC.n970 31.0582
R34916 VCC.t64 VCC.n1527 31.0582
R34917 VCC.t384 VCC.n2079 31.0582
R34918 VCC.t409 VCC.n2636 31.0582
R34919 VCC.t182 VCC.n3188 31.0582
R34920 VCC.t521 VCC.n3745 31.0582
R34921 VCC.t163 VCC.n4297 31.0582
R34922 VCC.t42 VCC.n4854 31.0582
R34923 VCC.t170 VCC.n5406 31.0582
R34924 VCC.t221 VCC.n5963 31.0582
R34925 VCC.t241 VCC.n6515 31.0582
R34926 VCC.t392 VCC.n7072 31.0582
R34927 VCC.t515 VCC.n7624 31.0582
R34928 VCC.t98 VCC.n8181 31.0582
R34929 VCC.t61 VCC.n8733 31.0582
R34930 VCC.t80 VCC.n9290 31.0582
R34931 VCC.t90 VCC.n9842 31.0582
R34932 VCC.t67 VCC.n10398 31.0582
R34933 VCC.t78 VCC.n10949 31.0582
R34934 VCC.t415 VCC.n11505 31.0582
R34935 VCC.t545 VCC.n12056 31.0582
R34936 VCC.t359 VCC.n12612 31.0582
R34937 VCC.t70 VCC.n13163 31.0582
R34938 VCC.t294 VCC.n13719 31.0582
R34939 VCC.t311 VCC.n14270 31.0582
R34940 VCC.t283 VCC.n14826 31.0582
R34941 VCC.t455 VCC.n15377 31.0582
R34942 VCC.t144 VCC.n15933 31.0582
R34943 VCC.t245 VCC.n16484 31.0582
R34944 VCC.t45 VCC.n17040 31.0582
R34945 VCC.t578 VCC.n17404 31.0582
R34946 VCC.n228 VCC.n153 29.2313
R34947 VCC.n268 VCC.n267 29.2313
R34948 VCC.n362 VCC.n361 29.2313
R34949 VCC.n395 VCC.n394 29.2313
R34950 VCC.n780 VCC.n705 29.2313
R34951 VCC.n820 VCC.n819 29.2313
R34952 VCC.n914 VCC.n913 29.2313
R34953 VCC.n947 VCC.n946 29.2313
R34954 VCC.n1471 VCC.n1470 29.2313
R34955 VCC.n1504 VCC.n1503 29.2313
R34956 VCC.n1338 VCC.n1263 29.2313
R34957 VCC.n1378 VCC.n1377 29.2313
R34958 VCC.n1889 VCC.n1814 29.2313
R34959 VCC.n1929 VCC.n1928 29.2313
R34960 VCC.n2023 VCC.n2022 29.2313
R34961 VCC.n2056 VCC.n2055 29.2313
R34962 VCC.n2580 VCC.n2579 29.2313
R34963 VCC.n2613 VCC.n2612 29.2313
R34964 VCC.n2447 VCC.n2372 29.2313
R34965 VCC.n2487 VCC.n2486 29.2313
R34966 VCC.n2998 VCC.n2923 29.2313
R34967 VCC.n3038 VCC.n3037 29.2313
R34968 VCC.n3132 VCC.n3131 29.2313
R34969 VCC.n3165 VCC.n3164 29.2313
R34970 VCC.n3689 VCC.n3688 29.2313
R34971 VCC.n3722 VCC.n3721 29.2313
R34972 VCC.n3556 VCC.n3481 29.2313
R34973 VCC.n3596 VCC.n3595 29.2313
R34974 VCC.n4107 VCC.n4032 29.2313
R34975 VCC.n4147 VCC.n4146 29.2313
R34976 VCC.n4241 VCC.n4240 29.2313
R34977 VCC.n4274 VCC.n4273 29.2313
R34978 VCC.n4798 VCC.n4797 29.2313
R34979 VCC.n4831 VCC.n4830 29.2313
R34980 VCC.n4665 VCC.n4590 29.2313
R34981 VCC.n4705 VCC.n4704 29.2313
R34982 VCC.n5216 VCC.n5141 29.2313
R34983 VCC.n5256 VCC.n5255 29.2313
R34984 VCC.n5350 VCC.n5349 29.2313
R34985 VCC.n5383 VCC.n5382 29.2313
R34986 VCC.n5907 VCC.n5906 29.2313
R34987 VCC.n5940 VCC.n5939 29.2313
R34988 VCC.n5774 VCC.n5699 29.2313
R34989 VCC.n5814 VCC.n5813 29.2313
R34990 VCC.n6325 VCC.n6250 29.2313
R34991 VCC.n6365 VCC.n6364 29.2313
R34992 VCC.n6459 VCC.n6458 29.2313
R34993 VCC.n6492 VCC.n6491 29.2313
R34994 VCC.n7016 VCC.n7015 29.2313
R34995 VCC.n7049 VCC.n7048 29.2313
R34996 VCC.n6883 VCC.n6808 29.2313
R34997 VCC.n6923 VCC.n6922 29.2313
R34998 VCC.n7434 VCC.n7359 29.2313
R34999 VCC.n7474 VCC.n7473 29.2313
R35000 VCC.n7568 VCC.n7567 29.2313
R35001 VCC.n7601 VCC.n7600 29.2313
R35002 VCC.n8125 VCC.n8124 29.2313
R35003 VCC.n8158 VCC.n8157 29.2313
R35004 VCC.n7992 VCC.n7917 29.2313
R35005 VCC.n8032 VCC.n8031 29.2313
R35006 VCC.n8677 VCC.n8676 29.2313
R35007 VCC.n8710 VCC.n8709 29.2313
R35008 VCC.n8543 VCC.n8468 29.2313
R35009 VCC.n8583 VCC.n8582 29.2313
R35010 VCC.n9234 VCC.n9233 29.2313
R35011 VCC.n9267 VCC.n9266 29.2313
R35012 VCC.n9101 VCC.n9026 29.2313
R35013 VCC.n9141 VCC.n9140 29.2313
R35014 VCC.n9652 VCC.n9577 29.2313
R35015 VCC.n9692 VCC.n9691 29.2313
R35016 VCC.n9786 VCC.n9785 29.2313
R35017 VCC.n9819 VCC.n9818 29.2313
R35018 VCC.n10342 VCC.n10341 29.2313
R35019 VCC.n10375 VCC.n10374 29.2313
R35020 VCC.n10209 VCC.n10134 29.2313
R35021 VCC.n10249 VCC.n10248 29.2313
R35022 VCC.n10759 VCC.n10684 29.2313
R35023 VCC.n10799 VCC.n10798 29.2313
R35024 VCC.n10893 VCC.n10892 29.2313
R35025 VCC.n10926 VCC.n10925 29.2313
R35026 VCC.n11449 VCC.n11448 29.2313
R35027 VCC.n11482 VCC.n11481 29.2313
R35028 VCC.n11316 VCC.n11241 29.2313
R35029 VCC.n11356 VCC.n11355 29.2313
R35030 VCC.n11866 VCC.n11791 29.2313
R35031 VCC.n11906 VCC.n11905 29.2313
R35032 VCC.n12000 VCC.n11999 29.2313
R35033 VCC.n12033 VCC.n12032 29.2313
R35034 VCC.n12556 VCC.n12555 29.2313
R35035 VCC.n12589 VCC.n12588 29.2313
R35036 VCC.n12423 VCC.n12348 29.2313
R35037 VCC.n12463 VCC.n12462 29.2313
R35038 VCC.n12973 VCC.n12898 29.2313
R35039 VCC.n13013 VCC.n13012 29.2313
R35040 VCC.n13107 VCC.n13106 29.2313
R35041 VCC.n13140 VCC.n13139 29.2313
R35042 VCC.n13663 VCC.n13662 29.2313
R35043 VCC.n13696 VCC.n13695 29.2313
R35044 VCC.n13530 VCC.n13455 29.2313
R35045 VCC.n13570 VCC.n13569 29.2313
R35046 VCC.n14080 VCC.n14005 29.2313
R35047 VCC.n14120 VCC.n14119 29.2313
R35048 VCC.n14214 VCC.n14213 29.2313
R35049 VCC.n14247 VCC.n14246 29.2313
R35050 VCC.n14770 VCC.n14769 29.2313
R35051 VCC.n14803 VCC.n14802 29.2313
R35052 VCC.n14637 VCC.n14562 29.2313
R35053 VCC.n14677 VCC.n14676 29.2313
R35054 VCC.n15187 VCC.n15112 29.2313
R35055 VCC.n15227 VCC.n15226 29.2313
R35056 VCC.n15321 VCC.n15320 29.2313
R35057 VCC.n15354 VCC.n15353 29.2313
R35058 VCC.n15877 VCC.n15876 29.2313
R35059 VCC.n15910 VCC.n15909 29.2313
R35060 VCC.n15744 VCC.n15669 29.2313
R35061 VCC.n15784 VCC.n15783 29.2313
R35062 VCC.n16294 VCC.n16219 29.2313
R35063 VCC.n16334 VCC.n16333 29.2313
R35064 VCC.n16428 VCC.n16427 29.2313
R35065 VCC.n16461 VCC.n16460 29.2313
R35066 VCC.n16984 VCC.n16983 29.2313
R35067 VCC.n17017 VCC.n17016 29.2313
R35068 VCC.n16851 VCC.n16776 29.2313
R35069 VCC.n16891 VCC.n16890 29.2313
R35070 VCC.n17348 VCC.n17347 29.2313
R35071 VCC.n17381 VCC.n17380 29.2313
R35072 VCC.n419 VCC.t189 26.3894
R35073 VCC.n494 VCC.n41 26.3894
R35074 VCC.n496 VCC.n22 26.3894
R35075 VCC.n971 VCC.t336 26.3894
R35076 VCC.n1046 VCC.n593 26.3894
R35077 VCC.n1048 VCC.n574 26.3894
R35078 VCC.n1529 VCC.t286 26.3894
R35079 VCC.n1584 VCC.n1583 26.3894
R35080 VCC.n1620 VCC.n1619 26.3894
R35081 VCC.n2080 VCC.t428 26.3894
R35082 VCC.n2155 VCC.n1702 26.3894
R35083 VCC.n2157 VCC.n1683 26.3894
R35084 VCC.n2638 VCC.t290 26.3894
R35085 VCC.n2693 VCC.n2692 26.3894
R35086 VCC.n2729 VCC.n2728 26.3894
R35087 VCC.n3189 VCC.t589 26.3894
R35088 VCC.n3264 VCC.n2811 26.3894
R35089 VCC.n3266 VCC.n2792 26.3894
R35090 VCC.n3747 VCC.t574 26.3894
R35091 VCC.n3802 VCC.n3801 26.3894
R35092 VCC.n3838 VCC.n3837 26.3894
R35093 VCC.n4298 VCC.t315 26.3894
R35094 VCC.n4373 VCC.n3920 26.3894
R35095 VCC.n4375 VCC.n3901 26.3894
R35096 VCC.n4856 VCC.t533 26.3894
R35097 VCC.n4911 VCC.n4910 26.3894
R35098 VCC.n4947 VCC.n4946 26.3894
R35099 VCC.n5407 VCC.t324 26.3894
R35100 VCC.n5482 VCC.n5029 26.3894
R35101 VCC.n5484 VCC.n5010 26.3894
R35102 VCC.n5965 VCC.t25 26.3894
R35103 VCC.n6020 VCC.n6019 26.3894
R35104 VCC.n6056 VCC.n6055 26.3894
R35105 VCC.n6516 VCC.t306 26.3894
R35106 VCC.n6591 VCC.n6138 26.3894
R35107 VCC.n6593 VCC.n6119 26.3894
R35108 VCC.n7074 VCC.t225 26.3894
R35109 VCC.n7129 VCC.n7128 26.3894
R35110 VCC.n7165 VCC.n7164 26.3894
R35111 VCC.n7625 VCC.t582 26.3894
R35112 VCC.n7700 VCC.n7247 26.3894
R35113 VCC.n7702 VCC.n7228 26.3894
R35114 VCC.n8183 VCC.t279 26.3894
R35115 VCC.n8238 VCC.n8237 26.3894
R35116 VCC.n8274 VCC.n8273 26.3894
R35117 VCC.n8734 VCC.t33 26.3894
R35118 VCC.n8809 VCC.n8356 26.3894
R35119 VCC.n8811 VCC.n8337 26.3894
R35120 VCC.n9292 VCC.t538 26.3894
R35121 VCC.n9347 VCC.n9346 26.3894
R35122 VCC.n9383 VCC.n9382 26.3894
R35123 VCC.n9843 VCC.t497 26.3894
R35124 VCC.n9918 VCC.n9465 26.3894
R35125 VCC.n9920 VCC.n9446 26.3894
R35126 VCC.n10400 VCC.t237 26.3894
R35127 VCC.n10455 VCC.n10454 26.3894
R35128 VCC.n10491 VCC.n10490 26.3894
R35129 VCC.n10950 VCC.t612 26.3894
R35130 VCC.n11025 VCC.n10572 26.3894
R35131 VCC.n11027 VCC.n10553 26.3894
R35132 VCC.n11507 VCC.t117 26.3894
R35133 VCC.n11562 VCC.n11561 26.3894
R35134 VCC.n11598 VCC.n11597 26.3894
R35135 VCC.n12057 VCC.t215 26.3894
R35136 VCC.n12132 VCC.n11679 26.3894
R35137 VCC.n12134 VCC.n11660 26.3894
R35138 VCC.n12614 VCC.t178 26.3894
R35139 VCC.n12669 VCC.n12668 26.3894
R35140 VCC.n12705 VCC.n12704 26.3894
R35141 VCC.n13164 VCC.t511 26.3894
R35142 VCC.n13239 VCC.n12786 26.3894
R35143 VCC.n13241 VCC.n12767 26.3894
R35144 VCC.n13721 VCC.t606 26.3894
R35145 VCC.n13776 VCC.n13775 26.3894
R35146 VCC.n13812 VCC.n13811 26.3894
R35147 VCC.n14271 VCC.t462 26.3894
R35148 VCC.n14346 VCC.n13893 26.3894
R35149 VCC.n14348 VCC.n13874 26.3894
R35150 VCC.n14828 VCC.t74 26.3894
R35151 VCC.n14883 VCC.n14882 26.3894
R35152 VCC.n14919 VCC.n14918 26.3894
R35153 VCC.n15378 VCC.t558 26.3894
R35154 VCC.n15453 VCC.n15000 26.3894
R35155 VCC.n15455 VCC.n14981 26.3894
R35156 VCC.n15935 VCC.t488 26.3894
R35157 VCC.n15990 VCC.n15989 26.3894
R35158 VCC.n16026 VCC.n16025 26.3894
R35159 VCC.n16485 VCC.t592 26.3894
R35160 VCC.n16560 VCC.n16107 26.3894
R35161 VCC.n16562 VCC.n16088 26.3894
R35162 VCC.n17042 VCC.t122 26.3894
R35163 VCC.n17097 VCC.n17096 26.3894
R35164 VCC.n17133 VCC.n17132 26.3894
R35165 VCC.n17405 VCC.t198 26.3894
R35166 VCC.n17480 VCC.n17214 26.3894
R35167 VCC.n17482 VCC.n17195 26.3894
R35168 VCC.n227 VCC.n226 25.5774
R35169 VCC.n290 VCC.n289 25.5774
R35170 VCC.n337 VCC.n108 25.5774
R35171 VCC.n417 VCC.n82 25.5774
R35172 VCC.n779 VCC.n778 25.5774
R35173 VCC.n842 VCC.n841 25.5774
R35174 VCC.n889 VCC.n660 25.5774
R35175 VCC.n969 VCC.n634 25.5774
R35176 VCC.n1446 VCC.n1217 25.5774
R35177 VCC.n1526 VCC.n1191 25.5774
R35178 VCC.n1337 VCC.n1336 25.5774
R35179 VCC.n1400 VCC.n1399 25.5774
R35180 VCC.n1888 VCC.n1887 25.5774
R35181 VCC.n1951 VCC.n1950 25.5774
R35182 VCC.n1998 VCC.n1769 25.5774
R35183 VCC.n2078 VCC.n1743 25.5774
R35184 VCC.n2555 VCC.n2326 25.5774
R35185 VCC.n2635 VCC.n2300 25.5774
R35186 VCC.n2446 VCC.n2445 25.5774
R35187 VCC.n2509 VCC.n2508 25.5774
R35188 VCC.n2997 VCC.n2996 25.5774
R35189 VCC.n3060 VCC.n3059 25.5774
R35190 VCC.n3107 VCC.n2878 25.5774
R35191 VCC.n3187 VCC.n2852 25.5774
R35192 VCC.n3664 VCC.n3435 25.5774
R35193 VCC.n3744 VCC.n3409 25.5774
R35194 VCC.n3555 VCC.n3554 25.5774
R35195 VCC.n3618 VCC.n3617 25.5774
R35196 VCC.n4106 VCC.n4105 25.5774
R35197 VCC.n4169 VCC.n4168 25.5774
R35198 VCC.n4216 VCC.n3987 25.5774
R35199 VCC.n4296 VCC.n3961 25.5774
R35200 VCC.n4773 VCC.n4544 25.5774
R35201 VCC.n4853 VCC.n4518 25.5774
R35202 VCC.n4664 VCC.n4663 25.5774
R35203 VCC.n4727 VCC.n4726 25.5774
R35204 VCC.n5215 VCC.n5214 25.5774
R35205 VCC.n5278 VCC.n5277 25.5774
R35206 VCC.n5325 VCC.n5096 25.5774
R35207 VCC.n5405 VCC.n5070 25.5774
R35208 VCC.n5882 VCC.n5653 25.5774
R35209 VCC.n5962 VCC.n5627 25.5774
R35210 VCC.n5773 VCC.n5772 25.5774
R35211 VCC.n5836 VCC.n5835 25.5774
R35212 VCC.n6324 VCC.n6323 25.5774
R35213 VCC.n6387 VCC.n6386 25.5774
R35214 VCC.n6434 VCC.n6205 25.5774
R35215 VCC.n6514 VCC.n6179 25.5774
R35216 VCC.n6991 VCC.n6762 25.5774
R35217 VCC.n7071 VCC.n6736 25.5774
R35218 VCC.n6882 VCC.n6881 25.5774
R35219 VCC.n6945 VCC.n6944 25.5774
R35220 VCC.n7433 VCC.n7432 25.5774
R35221 VCC.n7496 VCC.n7495 25.5774
R35222 VCC.n7543 VCC.n7314 25.5774
R35223 VCC.n7623 VCC.n7288 25.5774
R35224 VCC.n8100 VCC.n7871 25.5774
R35225 VCC.n8180 VCC.n7845 25.5774
R35226 VCC.n7991 VCC.n7990 25.5774
R35227 VCC.n8054 VCC.n8053 25.5774
R35228 VCC.n8652 VCC.n8423 25.5774
R35229 VCC.n8732 VCC.n8397 25.5774
R35230 VCC.n8542 VCC.n8541 25.5774
R35231 VCC.n8605 VCC.n8604 25.5774
R35232 VCC.n9209 VCC.n8980 25.5774
R35233 VCC.n9289 VCC.n8954 25.5774
R35234 VCC.n9100 VCC.n9099 25.5774
R35235 VCC.n9163 VCC.n9162 25.5774
R35236 VCC.n9651 VCC.n9650 25.5774
R35237 VCC.n9714 VCC.n9713 25.5774
R35238 VCC.n9761 VCC.n9532 25.5774
R35239 VCC.n9841 VCC.n9506 25.5774
R35240 VCC.n10317 VCC.n10088 25.5774
R35241 VCC.n10397 VCC.n10062 25.5774
R35242 VCC.n10208 VCC.n10207 25.5774
R35243 VCC.n10271 VCC.n10270 25.5774
R35244 VCC.n10758 VCC.n10757 25.5774
R35245 VCC.n10821 VCC.n10820 25.5774
R35246 VCC.n10868 VCC.n10639 25.5774
R35247 VCC.n10948 VCC.n10613 25.5774
R35248 VCC.n11424 VCC.n11195 25.5774
R35249 VCC.n11504 VCC.n11169 25.5774
R35250 VCC.n11315 VCC.n11314 25.5774
R35251 VCC.n11378 VCC.n11377 25.5774
R35252 VCC.n11865 VCC.n11864 25.5774
R35253 VCC.n11928 VCC.n11927 25.5774
R35254 VCC.n11975 VCC.n11746 25.5774
R35255 VCC.n12055 VCC.n11720 25.5774
R35256 VCC.n12531 VCC.n12302 25.5774
R35257 VCC.n12611 VCC.n12276 25.5774
R35258 VCC.n12422 VCC.n12421 25.5774
R35259 VCC.n12485 VCC.n12484 25.5774
R35260 VCC.n12972 VCC.n12971 25.5774
R35261 VCC.n13035 VCC.n13034 25.5774
R35262 VCC.n13082 VCC.n12853 25.5774
R35263 VCC.n13162 VCC.n12827 25.5774
R35264 VCC.n13638 VCC.n13409 25.5774
R35265 VCC.n13718 VCC.n13383 25.5774
R35266 VCC.n13529 VCC.n13528 25.5774
R35267 VCC.n13592 VCC.n13591 25.5774
R35268 VCC.n14079 VCC.n14078 25.5774
R35269 VCC.n14142 VCC.n14141 25.5774
R35270 VCC.n14189 VCC.n13960 25.5774
R35271 VCC.n14269 VCC.n13934 25.5774
R35272 VCC.n14745 VCC.n14516 25.5774
R35273 VCC.n14825 VCC.n14490 25.5774
R35274 VCC.n14636 VCC.n14635 25.5774
R35275 VCC.n14699 VCC.n14698 25.5774
R35276 VCC.n15186 VCC.n15185 25.5774
R35277 VCC.n15249 VCC.n15248 25.5774
R35278 VCC.n15296 VCC.n15067 25.5774
R35279 VCC.n15376 VCC.n15041 25.5774
R35280 VCC.n15852 VCC.n15623 25.5774
R35281 VCC.n15932 VCC.n15597 25.5774
R35282 VCC.n15743 VCC.n15742 25.5774
R35283 VCC.n15806 VCC.n15805 25.5774
R35284 VCC.n16293 VCC.n16292 25.5774
R35285 VCC.n16356 VCC.n16355 25.5774
R35286 VCC.n16403 VCC.n16174 25.5774
R35287 VCC.n16483 VCC.n16148 25.5774
R35288 VCC.n16959 VCC.n16730 25.5774
R35289 VCC.n17039 VCC.n16704 25.5774
R35290 VCC.n16850 VCC.n16849 25.5774
R35291 VCC.n16913 VCC.n16912 25.5774
R35292 VCC.n17323 VCC.n17281 25.5774
R35293 VCC.n17403 VCC.n17255 25.5774
R35294 VCC.n336 VCC.t567 23.7505
R35295 VCC.n888 VCC.t390 23.7505
R35296 VCC.n1445 VCC.t296 23.7505
R35297 VCC.n1997 VCC.t553 23.7505
R35298 VCC.n2554 VCC.t479 23.7505
R35299 VCC.n3106 VCC.t327 23.7505
R35300 VCC.n3663 VCC.t161 23.7505
R35301 VCC.n4215 VCC.t158 23.7505
R35302 VCC.n4772 VCC.t443 23.7505
R35303 VCC.n5324 VCC.t101 23.7505
R35304 VCC.n5881 VCC.t250 23.7505
R35305 VCC.n6433 VCC.t148 23.7505
R35306 VCC.n6990 VCC.t202 23.7505
R35307 VCC.n7542 VCC.t96 23.7505
R35308 VCC.n8099 VCC.t125 23.7505
R35309 VCC.n8651 VCC.t475 23.7505
R35310 VCC.n9208 VCC.t275 23.7505
R35311 VCC.n9760 VCC.t482 23.7505
R35312 VCC.n10316 VCC.t542 23.7505
R35313 VCC.n10867 VCC.t219 23.7505
R35314 VCC.n11423 VCC.t452 23.7505
R35315 VCC.n11974 VCC.t87 23.7505
R35316 VCC.n12530 VCC.t547 23.7505
R35317 VCC.n13081 VCC.t212 23.7505
R35318 VCC.n13637 VCC.t309 23.7505
R35319 VCC.n14188 VCC.t586 23.7505
R35320 VCC.n14744 VCC.t131 23.7505
R35321 VCC.n15295 VCC.t340 23.7505
R35322 VCC.n15851 VCC.t8 23.7505
R35323 VCC.n16402 VCC.t518 23.7505
R35324 VCC.n16958 VCC.t347 23.7505
R35325 VCC.n17322 VCC.t369 23.7505
R35326 VCC.n473 VCC.n471 22.8709
R35327 VCC.n526 VCC.t330 22.8709
R35328 VCC.n527 VCC.n526 22.8709
R35329 VCC.n1025 VCC.n1023 22.8709
R35330 VCC.n1078 VCC.t185 22.8709
R35331 VCC.n1079 VCC.n1078 22.8709
R35332 VCC.n1581 VCC.n1580 22.8709
R35333 VCC.t343 VCC.n1114 22.8709
R35334 VCC.n1651 VCC.n1114 22.8709
R35335 VCC.n2134 VCC.n2132 22.8709
R35336 VCC.n2187 VCC.t434 22.8709
R35337 VCC.n2188 VCC.n2187 22.8709
R35338 VCC.n2690 VCC.n2689 22.8709
R35339 VCC.t111 VCC.n2223 22.8709
R35340 VCC.n2760 VCC.n2223 22.8709
R35341 VCC.n3243 VCC.n3241 22.8709
R35342 VCC.n3296 VCC.t372 22.8709
R35343 VCC.n3297 VCC.n3296 22.8709
R35344 VCC.n3799 VCC.n3798 22.8709
R35345 VCC.t155 VCC.n3332 22.8709
R35346 VCC.n3869 VCC.n3332 22.8709
R35347 VCC.n4352 VCC.n4350 22.8709
R35348 VCC.n4405 VCC.t38 22.8709
R35349 VCC.n4406 VCC.n4405 22.8709
R35350 VCC.n4908 VCC.n4907 22.8709
R35351 VCC.t459 VCC.n4441 22.8709
R35352 VCC.n4978 VCC.n4441 22.8709
R35353 VCC.n5461 VCC.n5459 22.8709
R35354 VCC.n5514 VCC.t0 22.8709
R35355 VCC.n5515 VCC.n5514 22.8709
R35356 VCC.n6017 VCC.n6016 22.8709
R35357 VCC.t440 VCC.n5550 22.8709
R35358 VCC.n6087 VCC.n5550 22.8709
R35359 VCC.n6570 VCC.n6568 22.8709
R35360 VCC.n6623 VCC.t256 22.8709
R35361 VCC.n6624 VCC.n6623 22.8709
R35362 VCC.n7126 VCC.n7125 22.8709
R35363 VCC.t53 VCC.n6659 22.8709
R35364 VCC.n7196 VCC.n6659 22.8709
R35365 VCC.n7679 VCC.n7677 22.8709
R35366 VCC.n7732 VCC.t168 22.8709
R35367 VCC.n7733 VCC.n7732 22.8709
R35368 VCC.n8235 VCC.n8234 22.8709
R35369 VCC.t376 VCC.n7768 22.8709
R35370 VCC.n8305 VCC.n7768 22.8709
R35371 VCC.n8788 VCC.n8786 22.8709
R35372 VCC.n8841 VCC.t446 22.8709
R35373 VCC.n8842 VCC.n8841 22.8709
R35374 VCC.n9344 VCC.n9343 22.8709
R35375 VCC.t402 VCC.n8877 22.8709
R35376 VCC.n9414 VCC.n8877 22.8709
R35377 VCC.n9897 VCC.n9895 22.8709
R35378 VCC.n9950 VCC.t494 22.8709
R35379 VCC.n9951 VCC.n9950 22.8709
R35380 VCC.n10452 VCC.n10451 22.8709
R35381 VCC.t356 VCC.n9985 22.8709
R35382 VCC.n10522 VCC.n9985 22.8709
R35383 VCC.n11004 VCC.n11002 22.8709
R35384 VCC.n11057 VCC.t31 22.8709
R35385 VCC.n11058 VCC.n11057 22.8709
R35386 VCC.n11559 VCC.n11558 22.8709
R35387 VCC.t14 VCC.n11092 22.8709
R35388 VCC.n11629 VCC.n11092 22.8709
R35389 VCC.n12111 VCC.n12109 22.8709
R35390 VCC.n12164 VCC.t501 22.8709
R35391 VCC.n12165 VCC.n12164 22.8709
R35392 VCC.n12666 VCC.n12665 22.8709
R35393 VCC.t397 VCC.n12199 22.8709
R35394 VCC.n12736 VCC.n12199 22.8709
R35395 VCC.n13218 VCC.n13216 22.8709
R35396 VCC.n13271 VCC.t267 22.8709
R35397 VCC.n13272 VCC.n13271 22.8709
R35398 VCC.n13773 VCC.n13772 22.8709
R35399 VCC.t134 VCC.n13306 22.8709
R35400 VCC.n13843 VCC.n13306 22.8709
R35401 VCC.n14325 VCC.n14323 22.8709
R35402 VCC.n14378 VCC.t571 22.8709
R35403 VCC.n14379 VCC.n14378 22.8709
R35404 VCC.n14880 VCC.n14879 22.8709
R35405 VCC.t472 VCC.n14413 22.8709
R35406 VCC.n14950 VCC.n14413 22.8709
R35407 VCC.n15432 VCC.n15430 22.8709
R35408 VCC.n15485 VCC.t507 22.8709
R35409 VCC.n15486 VCC.n15485 22.8709
R35410 VCC.n15987 VCC.n15986 22.8709
R35411 VCC.t58 VCC.n15520 22.8709
R35412 VCC.n16057 VCC.n15520 22.8709
R35413 VCC.n16539 VCC.n16537 22.8709
R35414 VCC.n16592 VCC.t174 22.8709
R35415 VCC.n16593 VCC.n16592 22.8709
R35416 VCC.n17094 VCC.n17093 22.8709
R35417 VCC.t565 VCC.n16627 22.8709
R35418 VCC.n17164 VCC.n16627 22.8709
R35419 VCC.n17459 VCC.n17457 22.8709
R35420 VCC.n17512 VCC.t624 22.8709
R35421 VCC.n17513 VCC.n17512 22.8709
R35422 VCC.n211 VCC.n210 21.9236
R35423 VCC.t232 VCC.n181 21.9236
R35424 VCC.n335 VCC.n120 21.9236
R35425 VCC.n428 VCC.n427 21.9236
R35426 VCC.n763 VCC.n762 21.9236
R35427 VCC.t387 VCC.n733 21.9236
R35428 VCC.n887 VCC.n672 21.9236
R35429 VCC.n980 VCC.n979 21.9236
R35430 VCC.n1444 VCC.n1229 21.9236
R35431 VCC.n1538 VCC.n1537 21.9236
R35432 VCC.n1321 VCC.n1320 21.9236
R35433 VCC.t485 VCC.n1291 21.9236
R35434 VCC.n1872 VCC.n1871 21.9236
R35435 VCC.t18 VCC.n1842 21.9236
R35436 VCC.n1996 VCC.n1781 21.9236
R35437 VCC.n2089 VCC.n2088 21.9236
R35438 VCC.n2553 VCC.n2338 21.9236
R35439 VCC.n2647 VCC.n2646 21.9236
R35440 VCC.n2430 VCC.n2429 21.9236
R35441 VCC.t141 VCC.n2400 21.9236
R35442 VCC.n2981 VCC.n2980 21.9236
R35443 VCC.t599 VCC.n2951 21.9236
R35444 VCC.n3105 VCC.n2890 21.9236
R35445 VCC.n3198 VCC.n3197 21.9236
R35446 VCC.n3662 VCC.n3447 21.9236
R35447 VCC.n3756 VCC.n3755 21.9236
R35448 VCC.n3539 VCC.n3538 21.9236
R35449 VCC.t4 VCC.n3509 21.9236
R35450 VCC.n4090 VCC.n4089 21.9236
R35451 VCC.t551 VCC.n4060 21.9236
R35452 VCC.n4214 VCC.n3999 21.9236
R35453 VCC.n4307 VCC.n4306 21.9236
R35454 VCC.n4771 VCC.n4556 21.9236
R35455 VCC.n4865 VCC.n4864 21.9236
R35456 VCC.n4648 VCC.n4647 21.9236
R35457 VCC.t412 VCC.n4618 21.9236
R35458 VCC.n5199 VCC.n5198 21.9236
R35459 VCC.t350 VCC.n5169 21.9236
R35460 VCC.n5323 VCC.n5108 21.9236
R35461 VCC.n5416 VCC.n5415 21.9236
R35462 VCC.n5880 VCC.n5665 21.9236
R35463 VCC.n5974 VCC.n5973 21.9236
R35464 VCC.n5757 VCC.n5756 21.9236
R35465 VCC.t621 VCC.n5727 21.9236
R35466 VCC.n6308 VCC.n6307 21.9236
R35467 VCC.t332 VCC.n6278 21.9236
R35468 VCC.n6432 VCC.n6217 21.9236
R35469 VCC.n6525 VCC.n6524 21.9236
R35470 VCC.n6989 VCC.n6774 21.9236
R35471 VCC.n7083 VCC.n7082 21.9236
R35472 VCC.n6866 VCC.n6865 21.9236
R35473 VCC.t235 VCC.n6836 21.9236
R35474 VCC.n7417 VCC.n7416 21.9236
R35475 VCC.t601 VCC.n7387 21.9236
R35476 VCC.n7541 VCC.n7326 21.9236
R35477 VCC.n7634 VCC.n7633 21.9236
R35478 VCC.n8098 VCC.n7883 21.9236
R35479 VCC.n8192 VCC.n8191 21.9236
R35480 VCC.n7975 VCC.n7974 21.9236
R35481 VCC.t105 VCC.n7945 21.9236
R35482 VCC.n8650 VCC.n8435 21.9236
R35483 VCC.n8743 VCC.n8742 21.9236
R35484 VCC.n8526 VCC.n8525 21.9236
R35485 VCC.t83 VCC.n8496 21.9236
R35486 VCC.n9207 VCC.n8992 21.9236
R35487 VCC.n9301 VCC.n9300 21.9236
R35488 VCC.n9084 VCC.n9083 21.9236
R35489 VCC.t422 VCC.n9054 21.9236
R35490 VCC.n9635 VCC.n9634 21.9236
R35491 VCC.t321 VCC.n9605 21.9236
R35492 VCC.n9759 VCC.n9544 21.9236
R35493 VCC.n9852 VCC.n9851 21.9236
R35494 VCC.n10315 VCC.n10100 21.9236
R35495 VCC.n10409 VCC.n10408 21.9236
R35496 VCC.n10192 VCC.n10191 21.9236
R35497 VCC.t47 VCC.n10162 21.9236
R35498 VCC.n10742 VCC.n10741 21.9236
R35499 VCC.t22 VCC.n10712 21.9236
R35500 VCC.n10866 VCC.n10651 21.9236
R35501 VCC.n10959 VCC.n10958 21.9236
R35502 VCC.n11422 VCC.n11207 21.9236
R35503 VCC.n11516 VCC.n11515 21.9236
R35504 VCC.n11299 VCC.n11298 21.9236
R35505 VCC.t228 VCC.n11269 21.9236
R35506 VCC.n11849 VCC.n11848 21.9236
R35507 VCC.t505 VCC.n11819 21.9236
R35508 VCC.n11973 VCC.n11758 21.9236
R35509 VCC.n12066 VCC.n12065 21.9236
R35510 VCC.n12529 VCC.n12314 21.9236
R35511 VCC.n12623 VCC.n12622 21.9236
R35512 VCC.n12406 VCC.n12405 21.9236
R35513 VCC.t261 VCC.n12376 21.9236
R35514 VCC.n12956 VCC.n12955 21.9236
R35515 VCC.t560 VCC.n12926 21.9236
R35516 VCC.n13080 VCC.n12865 21.9236
R35517 VCC.n13173 VCC.n13172 21.9236
R35518 VCC.n13636 VCC.n13421 21.9236
R35519 VCC.n13730 VCC.n13729 21.9236
R35520 VCC.n13513 VCC.n13512 21.9236
R35521 VCC.t628 VCC.n13483 21.9236
R35522 VCC.n14063 VCC.n14062 21.9236
R35523 VCC.t208 VCC.n14033 21.9236
R35524 VCC.n14187 VCC.n13972 21.9236
R35525 VCC.n14280 VCC.n14279 21.9236
R35526 VCC.n14743 VCC.n14528 21.9236
R35527 VCC.n14837 VCC.n14836 21.9236
R35528 VCC.n14620 VCC.n14619 21.9236
R35529 VCC.t353 VCC.n14590 21.9236
R35530 VCC.n15170 VCC.n15169 21.9236
R35531 VCC.t50 VCC.n15140 21.9236
R35532 VCC.n15294 VCC.n15079 21.9236
R35533 VCC.n15387 VCC.n15386 21.9236
R35534 VCC.n15850 VCC.n15635 21.9236
R35535 VCC.n15944 VCC.n15943 21.9236
R35536 VCC.n15727 VCC.n15726 21.9236
R35537 VCC.t527 VCC.n15697 21.9236
R35538 VCC.n16277 VCC.n16276 21.9236
R35539 VCC.t419 VCC.n16247 21.9236
R35540 VCC.n16401 VCC.n16186 21.9236
R35541 VCC.n16494 VCC.n16493 21.9236
R35542 VCC.n16957 VCC.n16742 21.9236
R35543 VCC.n17051 VCC.n17050 21.9236
R35544 VCC.n16834 VCC.n16833 21.9236
R35545 VCC.t608 VCC.n16804 21.9236
R35546 VCC.n17321 VCC.n17293 21.9236
R35547 VCC.n17414 VCC.n17413 21.9236
R35548 VCC.n420 VCC.n419 19.3524
R35549 VCC.n972 VCC.n971 19.3524
R35550 VCC.n1529 VCC.n1528 19.3524
R35551 VCC.n2081 VCC.n2080 19.3524
R35552 VCC.n2638 VCC.n2637 19.3524
R35553 VCC.n3190 VCC.n3189 19.3524
R35554 VCC.n3747 VCC.n3746 19.3524
R35555 VCC.n4299 VCC.n4298 19.3524
R35556 VCC.n4856 VCC.n4855 19.3524
R35557 VCC.n5408 VCC.n5407 19.3524
R35558 VCC.n5965 VCC.n5964 19.3524
R35559 VCC.n6517 VCC.n6516 19.3524
R35560 VCC.n7074 VCC.n7073 19.3524
R35561 VCC.n7626 VCC.n7625 19.3524
R35562 VCC.n8183 VCC.n8182 19.3524
R35563 VCC.n8735 VCC.n8734 19.3524
R35564 VCC.n9292 VCC.n9291 19.3524
R35565 VCC.n9844 VCC.n9843 19.3524
R35566 VCC.n10400 VCC.n10399 19.3524
R35567 VCC.n10951 VCC.n10950 19.3524
R35568 VCC.n11507 VCC.n11506 19.3524
R35569 VCC.n12058 VCC.n12057 19.3524
R35570 VCC.n12614 VCC.n12613 19.3524
R35571 VCC.n13165 VCC.n13164 19.3524
R35572 VCC.n13721 VCC.n13720 19.3524
R35573 VCC.n14272 VCC.n14271 19.3524
R35574 VCC.n14828 VCC.n14827 19.3524
R35575 VCC.n15379 VCC.n15378 19.3524
R35576 VCC.n15935 VCC.n15934 19.3524
R35577 VCC.n16486 VCC.n16485 19.3524
R35578 VCC.n17042 VCC.n17041 19.3524
R35579 VCC.n17406 VCC.n17405 19.3524
R35580 VCC.n180 VCC.n154 15.2005
R35581 VCC.n269 VCC.n152 15.2005
R35582 VCC.n363 VCC.n107 15.2005
R35583 VCC.n393 VCC.n92 15.2005
R35584 VCC.n732 VCC.n706 15.2005
R35585 VCC.n821 VCC.n704 15.2005
R35586 VCC.n915 VCC.n659 15.2005
R35587 VCC.n945 VCC.n644 15.2005
R35588 VCC.n1472 VCC.n1216 15.2005
R35589 VCC.n1502 VCC.n1201 15.2005
R35590 VCC.n1290 VCC.n1264 15.2005
R35591 VCC.n1379 VCC.n1262 15.2005
R35592 VCC.n1841 VCC.n1815 15.2005
R35593 VCC.n1930 VCC.n1813 15.2005
R35594 VCC.n2024 VCC.n1768 15.2005
R35595 VCC.n2054 VCC.n1753 15.2005
R35596 VCC.n2581 VCC.n2325 15.2005
R35597 VCC.n2611 VCC.n2310 15.2005
R35598 VCC.n2399 VCC.n2373 15.2005
R35599 VCC.n2488 VCC.n2371 15.2005
R35600 VCC.n2950 VCC.n2924 15.2005
R35601 VCC.n3039 VCC.n2922 15.2005
R35602 VCC.n3133 VCC.n2877 15.2005
R35603 VCC.n3163 VCC.n2862 15.2005
R35604 VCC.n3690 VCC.n3434 15.2005
R35605 VCC.n3720 VCC.n3419 15.2005
R35606 VCC.n3508 VCC.n3482 15.2005
R35607 VCC.n3597 VCC.n3480 15.2005
R35608 VCC.n4059 VCC.n4033 15.2005
R35609 VCC.n4148 VCC.n4031 15.2005
R35610 VCC.n4242 VCC.n3986 15.2005
R35611 VCC.n4272 VCC.n3971 15.2005
R35612 VCC.n4799 VCC.n4543 15.2005
R35613 VCC.n4829 VCC.n4528 15.2005
R35614 VCC.n4617 VCC.n4591 15.2005
R35615 VCC.n4706 VCC.n4589 15.2005
R35616 VCC.n5168 VCC.n5142 15.2005
R35617 VCC.n5257 VCC.n5140 15.2005
R35618 VCC.n5351 VCC.n5095 15.2005
R35619 VCC.n5381 VCC.n5080 15.2005
R35620 VCC.n5908 VCC.n5652 15.2005
R35621 VCC.n5938 VCC.n5637 15.2005
R35622 VCC.n5726 VCC.n5700 15.2005
R35623 VCC.n5815 VCC.n5698 15.2005
R35624 VCC.n6277 VCC.n6251 15.2005
R35625 VCC.n6366 VCC.n6249 15.2005
R35626 VCC.n6460 VCC.n6204 15.2005
R35627 VCC.n6490 VCC.n6189 15.2005
R35628 VCC.n7017 VCC.n6761 15.2005
R35629 VCC.n7047 VCC.n6746 15.2005
R35630 VCC.n6835 VCC.n6809 15.2005
R35631 VCC.n6924 VCC.n6807 15.2005
R35632 VCC.n7386 VCC.n7360 15.2005
R35633 VCC.n7475 VCC.n7358 15.2005
R35634 VCC.n7569 VCC.n7313 15.2005
R35635 VCC.n7599 VCC.n7298 15.2005
R35636 VCC.n8126 VCC.n7870 15.2005
R35637 VCC.n8156 VCC.n7855 15.2005
R35638 VCC.n7944 VCC.n7918 15.2005
R35639 VCC.n8033 VCC.n7916 15.2005
R35640 VCC.n8678 VCC.n8422 15.2005
R35641 VCC.n8708 VCC.n8407 15.2005
R35642 VCC.n8495 VCC.n8469 15.2005
R35643 VCC.n8584 VCC.n8467 15.2005
R35644 VCC.n9235 VCC.n8979 15.2005
R35645 VCC.n9265 VCC.n8964 15.2005
R35646 VCC.n9053 VCC.n9027 15.2005
R35647 VCC.n9142 VCC.n9025 15.2005
R35648 VCC.n9604 VCC.n9578 15.2005
R35649 VCC.n9693 VCC.n9576 15.2005
R35650 VCC.n9787 VCC.n9531 15.2005
R35651 VCC.n9817 VCC.n9516 15.2005
R35652 VCC.n10343 VCC.n10087 15.2005
R35653 VCC.n10373 VCC.n10072 15.2005
R35654 VCC.n10161 VCC.n10135 15.2005
R35655 VCC.n10250 VCC.n10133 15.2005
R35656 VCC.n10711 VCC.n10685 15.2005
R35657 VCC.n10800 VCC.n10683 15.2005
R35658 VCC.n10894 VCC.n10638 15.2005
R35659 VCC.n10924 VCC.n10623 15.2005
R35660 VCC.n11450 VCC.n11194 15.2005
R35661 VCC.n11480 VCC.n11179 15.2005
R35662 VCC.n11268 VCC.n11242 15.2005
R35663 VCC.n11357 VCC.n11240 15.2005
R35664 VCC.n11818 VCC.n11792 15.2005
R35665 VCC.n11907 VCC.n11790 15.2005
R35666 VCC.n12001 VCC.n11745 15.2005
R35667 VCC.n12031 VCC.n11730 15.2005
R35668 VCC.n12557 VCC.n12301 15.2005
R35669 VCC.n12587 VCC.n12286 15.2005
R35670 VCC.n12375 VCC.n12349 15.2005
R35671 VCC.n12464 VCC.n12347 15.2005
R35672 VCC.n12925 VCC.n12899 15.2005
R35673 VCC.n13014 VCC.n12897 15.2005
R35674 VCC.n13108 VCC.n12852 15.2005
R35675 VCC.n13138 VCC.n12837 15.2005
R35676 VCC.n13664 VCC.n13408 15.2005
R35677 VCC.n13694 VCC.n13393 15.2005
R35678 VCC.n13482 VCC.n13456 15.2005
R35679 VCC.n13571 VCC.n13454 15.2005
R35680 VCC.n14032 VCC.n14006 15.2005
R35681 VCC.n14121 VCC.n14004 15.2005
R35682 VCC.n14215 VCC.n13959 15.2005
R35683 VCC.n14245 VCC.n13944 15.2005
R35684 VCC.n14771 VCC.n14515 15.2005
R35685 VCC.n14801 VCC.n14500 15.2005
R35686 VCC.n14589 VCC.n14563 15.2005
R35687 VCC.n14678 VCC.n14561 15.2005
R35688 VCC.n15139 VCC.n15113 15.2005
R35689 VCC.n15228 VCC.n15111 15.2005
R35690 VCC.n15322 VCC.n15066 15.2005
R35691 VCC.n15352 VCC.n15051 15.2005
R35692 VCC.n15878 VCC.n15622 15.2005
R35693 VCC.n15908 VCC.n15607 15.2005
R35694 VCC.n15696 VCC.n15670 15.2005
R35695 VCC.n15785 VCC.n15668 15.2005
R35696 VCC.n16246 VCC.n16220 15.2005
R35697 VCC.n16335 VCC.n16218 15.2005
R35698 VCC.n16429 VCC.n16173 15.2005
R35699 VCC.n16459 VCC.n16158 15.2005
R35700 VCC.n16985 VCC.n16729 15.2005
R35701 VCC.n17015 VCC.n16714 15.2005
R35702 VCC.n16803 VCC.n16777 15.2005
R35703 VCC.n16892 VCC.n16775 15.2005
R35704 VCC.n17349 VCC.n17280 15.2005
R35705 VCC.n17379 VCC.n17265 15.2005
R35706 VCC.n225 VCC.n179 13.3005
R35707 VCC.n288 VCC.n140 13.3005
R35708 VCC.n338 VCC.n109 13.3005
R35709 VCC.n416 VCC.n83 13.3005
R35710 VCC.n777 VCC.n731 13.3005
R35711 VCC.n840 VCC.n692 13.3005
R35712 VCC.n890 VCC.n661 13.3005
R35713 VCC.n968 VCC.n635 13.3005
R35714 VCC.n1447 VCC.n1218 13.3005
R35715 VCC.n1525 VCC.n1192 13.3005
R35716 VCC.n1335 VCC.n1289 13.3005
R35717 VCC.n1398 VCC.n1250 13.3005
R35718 VCC.n1886 VCC.n1840 13.3005
R35719 VCC.n1949 VCC.n1801 13.3005
R35720 VCC.n1999 VCC.n1770 13.3005
R35721 VCC.n2077 VCC.n1744 13.3005
R35722 VCC.n2556 VCC.n2327 13.3005
R35723 VCC.n2634 VCC.n2301 13.3005
R35724 VCC.n2444 VCC.n2398 13.3005
R35725 VCC.n2507 VCC.n2359 13.3005
R35726 VCC.n2995 VCC.n2949 13.3005
R35727 VCC.n3058 VCC.n2910 13.3005
R35728 VCC.n3108 VCC.n2879 13.3005
R35729 VCC.n3186 VCC.n2853 13.3005
R35730 VCC.n3665 VCC.n3436 13.3005
R35731 VCC.n3743 VCC.n3410 13.3005
R35732 VCC.n3553 VCC.n3507 13.3005
R35733 VCC.n3616 VCC.n3468 13.3005
R35734 VCC.n4104 VCC.n4058 13.3005
R35735 VCC.n4167 VCC.n4019 13.3005
R35736 VCC.n4217 VCC.n3988 13.3005
R35737 VCC.n4295 VCC.n3962 13.3005
R35738 VCC.n4774 VCC.n4545 13.3005
R35739 VCC.n4852 VCC.n4519 13.3005
R35740 VCC.n4662 VCC.n4616 13.3005
R35741 VCC.n4725 VCC.n4577 13.3005
R35742 VCC.n5213 VCC.n5167 13.3005
R35743 VCC.n5276 VCC.n5128 13.3005
R35744 VCC.n5326 VCC.n5097 13.3005
R35745 VCC.n5404 VCC.n5071 13.3005
R35746 VCC.n5883 VCC.n5654 13.3005
R35747 VCC.n5961 VCC.n5628 13.3005
R35748 VCC.n5771 VCC.n5725 13.3005
R35749 VCC.n5834 VCC.n5686 13.3005
R35750 VCC.n6322 VCC.n6276 13.3005
R35751 VCC.n6385 VCC.n6237 13.3005
R35752 VCC.n6435 VCC.n6206 13.3005
R35753 VCC.n6513 VCC.n6180 13.3005
R35754 VCC.n6992 VCC.n6763 13.3005
R35755 VCC.n7070 VCC.n6737 13.3005
R35756 VCC.n6880 VCC.n6834 13.3005
R35757 VCC.n6943 VCC.n6795 13.3005
R35758 VCC.n7431 VCC.n7385 13.3005
R35759 VCC.n7494 VCC.n7346 13.3005
R35760 VCC.n7544 VCC.n7315 13.3005
R35761 VCC.n7622 VCC.n7289 13.3005
R35762 VCC.n8101 VCC.n7872 13.3005
R35763 VCC.n8179 VCC.n7846 13.3005
R35764 VCC.n7989 VCC.n7943 13.3005
R35765 VCC.n8052 VCC.n7904 13.3005
R35766 VCC.n8653 VCC.n8424 13.3005
R35767 VCC.n8731 VCC.n8398 13.3005
R35768 VCC.n8540 VCC.n8494 13.3005
R35769 VCC.n8603 VCC.n8455 13.3005
R35770 VCC.n9210 VCC.n8981 13.3005
R35771 VCC.n9288 VCC.n8955 13.3005
R35772 VCC.n9098 VCC.n9052 13.3005
R35773 VCC.n9161 VCC.n9013 13.3005
R35774 VCC.n9649 VCC.n9603 13.3005
R35775 VCC.n9712 VCC.n9564 13.3005
R35776 VCC.n9762 VCC.n9533 13.3005
R35777 VCC.n9840 VCC.n9507 13.3005
R35778 VCC.n10318 VCC.n10089 13.3005
R35779 VCC.n10396 VCC.n10063 13.3005
R35780 VCC.n10206 VCC.n10160 13.3005
R35781 VCC.n10269 VCC.n10121 13.3005
R35782 VCC.n10756 VCC.n10710 13.3005
R35783 VCC.n10819 VCC.n10671 13.3005
R35784 VCC.n10869 VCC.n10640 13.3005
R35785 VCC.n10947 VCC.n10614 13.3005
R35786 VCC.n11425 VCC.n11196 13.3005
R35787 VCC.n11503 VCC.n11170 13.3005
R35788 VCC.n11313 VCC.n11267 13.3005
R35789 VCC.n11376 VCC.n11228 13.3005
R35790 VCC.n11863 VCC.n11817 13.3005
R35791 VCC.n11926 VCC.n11778 13.3005
R35792 VCC.n11976 VCC.n11747 13.3005
R35793 VCC.n12054 VCC.n11721 13.3005
R35794 VCC.n12532 VCC.n12303 13.3005
R35795 VCC.n12610 VCC.n12277 13.3005
R35796 VCC.n12420 VCC.n12374 13.3005
R35797 VCC.n12483 VCC.n12335 13.3005
R35798 VCC.n12970 VCC.n12924 13.3005
R35799 VCC.n13033 VCC.n12885 13.3005
R35800 VCC.n13083 VCC.n12854 13.3005
R35801 VCC.n13161 VCC.n12828 13.3005
R35802 VCC.n13639 VCC.n13410 13.3005
R35803 VCC.n13717 VCC.n13384 13.3005
R35804 VCC.n13527 VCC.n13481 13.3005
R35805 VCC.n13590 VCC.n13442 13.3005
R35806 VCC.n14077 VCC.n14031 13.3005
R35807 VCC.n14140 VCC.n13992 13.3005
R35808 VCC.n14190 VCC.n13961 13.3005
R35809 VCC.n14268 VCC.n13935 13.3005
R35810 VCC.n14746 VCC.n14517 13.3005
R35811 VCC.n14824 VCC.n14491 13.3005
R35812 VCC.n14634 VCC.n14588 13.3005
R35813 VCC.n14697 VCC.n14549 13.3005
R35814 VCC.n15184 VCC.n15138 13.3005
R35815 VCC.n15247 VCC.n15099 13.3005
R35816 VCC.n15297 VCC.n15068 13.3005
R35817 VCC.n15375 VCC.n15042 13.3005
R35818 VCC.n15853 VCC.n15624 13.3005
R35819 VCC.n15931 VCC.n15598 13.3005
R35820 VCC.n15741 VCC.n15695 13.3005
R35821 VCC.n15804 VCC.n15656 13.3005
R35822 VCC.n16291 VCC.n16245 13.3005
R35823 VCC.n16354 VCC.n16206 13.3005
R35824 VCC.n16404 VCC.n16175 13.3005
R35825 VCC.n16482 VCC.n16149 13.3005
R35826 VCC.n16960 VCC.n16731 13.3005
R35827 VCC.n17038 VCC.n16705 13.3005
R35828 VCC.n16848 VCC.n16802 13.3005
R35829 VCC.n16911 VCC.n16763 13.3005
R35830 VCC.n17324 VCC.n17282 13.3005
R35831 VCC.n17402 VCC.n17256 13.3005
R35832 VCC.n493 VCC.n492 12.2148
R35833 VCC.n497 VCC.n23 12.2148
R35834 VCC.n1045 VCC.n1044 12.2148
R35835 VCC.n1049 VCC.n575 12.2148
R35836 VCC.n1582 VCC.n1162 12.2148
R35837 VCC.n1618 VCC.n1142 12.2148
R35838 VCC.n2154 VCC.n2153 12.2148
R35839 VCC.n2158 VCC.n1684 12.2148
R35840 VCC.n2691 VCC.n2271 12.2148
R35841 VCC.n2727 VCC.n2251 12.2148
R35842 VCC.n3263 VCC.n3262 12.2148
R35843 VCC.n3267 VCC.n2793 12.2148
R35844 VCC.n3800 VCC.n3380 12.2148
R35845 VCC.n3836 VCC.n3360 12.2148
R35846 VCC.n4372 VCC.n4371 12.2148
R35847 VCC.n4376 VCC.n3902 12.2148
R35848 VCC.n4909 VCC.n4489 12.2148
R35849 VCC.n4945 VCC.n4469 12.2148
R35850 VCC.n5481 VCC.n5480 12.2148
R35851 VCC.n5485 VCC.n5011 12.2148
R35852 VCC.n6018 VCC.n5598 12.2148
R35853 VCC.n6054 VCC.n5578 12.2148
R35854 VCC.n6590 VCC.n6589 12.2148
R35855 VCC.n6594 VCC.n6120 12.2148
R35856 VCC.n7127 VCC.n6707 12.2148
R35857 VCC.n7163 VCC.n6687 12.2148
R35858 VCC.n7699 VCC.n7698 12.2148
R35859 VCC.n7703 VCC.n7229 12.2148
R35860 VCC.n8236 VCC.n7816 12.2148
R35861 VCC.n8272 VCC.n7796 12.2148
R35862 VCC.n8808 VCC.n8807 12.2148
R35863 VCC.n8812 VCC.n8338 12.2148
R35864 VCC.n9345 VCC.n8925 12.2148
R35865 VCC.n9381 VCC.n8905 12.2148
R35866 VCC.n9917 VCC.n9916 12.2148
R35867 VCC.n9921 VCC.n9447 12.2148
R35868 VCC.n10453 VCC.n10033 12.2148
R35869 VCC.n10489 VCC.n10013 12.2148
R35870 VCC.n11024 VCC.n11023 12.2148
R35871 VCC.n11028 VCC.n10554 12.2148
R35872 VCC.n11560 VCC.n11140 12.2148
R35873 VCC.n11596 VCC.n11120 12.2148
R35874 VCC.n12131 VCC.n12130 12.2148
R35875 VCC.n12135 VCC.n11661 12.2148
R35876 VCC.n12667 VCC.n12247 12.2148
R35877 VCC.n12703 VCC.n12227 12.2148
R35878 VCC.n13238 VCC.n13237 12.2148
R35879 VCC.n13242 VCC.n12768 12.2148
R35880 VCC.n13774 VCC.n13354 12.2148
R35881 VCC.n13810 VCC.n13334 12.2148
R35882 VCC.n14345 VCC.n14344 12.2148
R35883 VCC.n14349 VCC.n13875 12.2148
R35884 VCC.n14881 VCC.n14461 12.2148
R35885 VCC.n14917 VCC.n14441 12.2148
R35886 VCC.n15452 VCC.n15451 12.2148
R35887 VCC.n15456 VCC.n14982 12.2148
R35888 VCC.n15988 VCC.n15568 12.2148
R35889 VCC.n16024 VCC.n15548 12.2148
R35890 VCC.n16559 VCC.n16558 12.2148
R35891 VCC.n16563 VCC.n16089 12.2148
R35892 VCC.n17095 VCC.n16675 12.2148
R35893 VCC.n17131 VCC.n16655 12.2148
R35894 VCC.n17479 VCC.n17478 12.2148
R35895 VCC.n17483 VCC.n17196 12.2148
R35896 VCC.n212 VCC.n208 11.4005
R35897 VCC.n334 VCC.n121 11.4005
R35898 VCC.n429 VCC.n81 11.4005
R35899 VCC.n764 VCC.n760 11.4005
R35900 VCC.n886 VCC.n673 11.4005
R35901 VCC.n981 VCC.n633 11.4005
R35902 VCC.n1443 VCC.n1230 11.4005
R35903 VCC.n1539 VCC.n1190 11.4005
R35904 VCC.n1322 VCC.n1318 11.4005
R35905 VCC.n1873 VCC.n1869 11.4005
R35906 VCC.n1995 VCC.n1782 11.4005
R35907 VCC.n2090 VCC.n1742 11.4005
R35908 VCC.n2552 VCC.n2339 11.4005
R35909 VCC.n2648 VCC.n2299 11.4005
R35910 VCC.n2431 VCC.n2427 11.4005
R35911 VCC.n2982 VCC.n2978 11.4005
R35912 VCC.n3104 VCC.n2891 11.4005
R35913 VCC.n3199 VCC.n2851 11.4005
R35914 VCC.n3661 VCC.n3448 11.4005
R35915 VCC.n3757 VCC.n3408 11.4005
R35916 VCC.n3540 VCC.n3536 11.4005
R35917 VCC.n4091 VCC.n4087 11.4005
R35918 VCC.n4213 VCC.n4000 11.4005
R35919 VCC.n4308 VCC.n3960 11.4005
R35920 VCC.n4770 VCC.n4557 11.4005
R35921 VCC.n4866 VCC.n4517 11.4005
R35922 VCC.n4649 VCC.n4645 11.4005
R35923 VCC.n5200 VCC.n5196 11.4005
R35924 VCC.n5322 VCC.n5109 11.4005
R35925 VCC.n5417 VCC.n5069 11.4005
R35926 VCC.n5879 VCC.n5666 11.4005
R35927 VCC.n5975 VCC.n5626 11.4005
R35928 VCC.n5758 VCC.n5754 11.4005
R35929 VCC.n6309 VCC.n6305 11.4005
R35930 VCC.n6431 VCC.n6218 11.4005
R35931 VCC.n6526 VCC.n6178 11.4005
R35932 VCC.n6988 VCC.n6775 11.4005
R35933 VCC.n7084 VCC.n6735 11.4005
R35934 VCC.n6867 VCC.n6863 11.4005
R35935 VCC.n7418 VCC.n7414 11.4005
R35936 VCC.n7540 VCC.n7327 11.4005
R35937 VCC.n7635 VCC.n7287 11.4005
R35938 VCC.n8097 VCC.n7884 11.4005
R35939 VCC.n8193 VCC.n7844 11.4005
R35940 VCC.n7976 VCC.n7972 11.4005
R35941 VCC.n8649 VCC.n8436 11.4005
R35942 VCC.n8744 VCC.n8396 11.4005
R35943 VCC.n8527 VCC.n8523 11.4005
R35944 VCC.n9206 VCC.n8993 11.4005
R35945 VCC.n9302 VCC.n8953 11.4005
R35946 VCC.n9085 VCC.n9081 11.4005
R35947 VCC.n9636 VCC.n9632 11.4005
R35948 VCC.n9758 VCC.n9545 11.4005
R35949 VCC.n9853 VCC.n9505 11.4005
R35950 VCC.n10314 VCC.n10101 11.4005
R35951 VCC.n10410 VCC.n10061 11.4005
R35952 VCC.n10193 VCC.n10189 11.4005
R35953 VCC.n10743 VCC.n10739 11.4005
R35954 VCC.n10865 VCC.n10652 11.4005
R35955 VCC.n10960 VCC.n10612 11.4005
R35956 VCC.n11421 VCC.n11208 11.4005
R35957 VCC.n11517 VCC.n11168 11.4005
R35958 VCC.n11300 VCC.n11296 11.4005
R35959 VCC.n11850 VCC.n11846 11.4005
R35960 VCC.n11972 VCC.n11759 11.4005
R35961 VCC.n12067 VCC.n11719 11.4005
R35962 VCC.n12528 VCC.n12315 11.4005
R35963 VCC.n12624 VCC.n12275 11.4005
R35964 VCC.n12407 VCC.n12403 11.4005
R35965 VCC.n12957 VCC.n12953 11.4005
R35966 VCC.n13079 VCC.n12866 11.4005
R35967 VCC.n13174 VCC.n12826 11.4005
R35968 VCC.n13635 VCC.n13422 11.4005
R35969 VCC.n13731 VCC.n13382 11.4005
R35970 VCC.n13514 VCC.n13510 11.4005
R35971 VCC.n14064 VCC.n14060 11.4005
R35972 VCC.n14186 VCC.n13973 11.4005
R35973 VCC.n14281 VCC.n13933 11.4005
R35974 VCC.n14742 VCC.n14529 11.4005
R35975 VCC.n14838 VCC.n14489 11.4005
R35976 VCC.n14621 VCC.n14617 11.4005
R35977 VCC.n15171 VCC.n15167 11.4005
R35978 VCC.n15293 VCC.n15080 11.4005
R35979 VCC.n15388 VCC.n15040 11.4005
R35980 VCC.n15849 VCC.n15636 11.4005
R35981 VCC.n15945 VCC.n15596 11.4005
R35982 VCC.n15728 VCC.n15724 11.4005
R35983 VCC.n16278 VCC.n16274 11.4005
R35984 VCC.n16400 VCC.n16187 11.4005
R35985 VCC.n16495 VCC.n16147 11.4005
R35986 VCC.n16956 VCC.n16743 11.4005
R35987 VCC.n17052 VCC.n16703 11.4005
R35988 VCC.n16835 VCC.n16831 11.4005
R35989 VCC.n17320 VCC.n17294 11.4005
R35990 VCC.n17415 VCC.n17254 11.4005
R35991 VCC.n474 VCC.n55 10.5862
R35992 VCC.n528 VCC.n21 10.5862
R35993 VCC.n1026 VCC.n607 10.5862
R35994 VCC.n1080 VCC.n573 10.5862
R35995 VCC.n1579 VCC.n1161 10.5862
R35996 VCC.n1650 VCC.n1115 10.5862
R35997 VCC.n2135 VCC.n1716 10.5862
R35998 VCC.n2189 VCC.n1682 10.5862
R35999 VCC.n2688 VCC.n2270 10.5862
R36000 VCC.n2759 VCC.n2224 10.5862
R36001 VCC.n3244 VCC.n2825 10.5862
R36002 VCC.n3298 VCC.n2791 10.5862
R36003 VCC.n3797 VCC.n3379 10.5862
R36004 VCC.n3868 VCC.n3333 10.5862
R36005 VCC.n4353 VCC.n3934 10.5862
R36006 VCC.n4407 VCC.n3900 10.5862
R36007 VCC.n4906 VCC.n4488 10.5862
R36008 VCC.n4977 VCC.n4442 10.5862
R36009 VCC.n5462 VCC.n5043 10.5862
R36010 VCC.n5516 VCC.n5009 10.5862
R36011 VCC.n6015 VCC.n5597 10.5862
R36012 VCC.n6086 VCC.n5551 10.5862
R36013 VCC.n6571 VCC.n6152 10.5862
R36014 VCC.n6625 VCC.n6118 10.5862
R36015 VCC.n7124 VCC.n6706 10.5862
R36016 VCC.n7195 VCC.n6660 10.5862
R36017 VCC.n7680 VCC.n7261 10.5862
R36018 VCC.n7734 VCC.n7227 10.5862
R36019 VCC.n8233 VCC.n7815 10.5862
R36020 VCC.n8304 VCC.n7769 10.5862
R36021 VCC.n8789 VCC.n8370 10.5862
R36022 VCC.n8843 VCC.n8336 10.5862
R36023 VCC.n9342 VCC.n8924 10.5862
R36024 VCC.n9413 VCC.n8878 10.5862
R36025 VCC.n9898 VCC.n9479 10.5862
R36026 VCC.n9952 VCC.n9445 10.5862
R36027 VCC.n10450 VCC.n10032 10.5862
R36028 VCC.n10521 VCC.n9986 10.5862
R36029 VCC.n11005 VCC.n10586 10.5862
R36030 VCC.n11059 VCC.n10552 10.5862
R36031 VCC.n11557 VCC.n11139 10.5862
R36032 VCC.n11628 VCC.n11093 10.5862
R36033 VCC.n12112 VCC.n11693 10.5862
R36034 VCC.n12166 VCC.n11659 10.5862
R36035 VCC.n12664 VCC.n12246 10.5862
R36036 VCC.n12735 VCC.n12200 10.5862
R36037 VCC.n13219 VCC.n12800 10.5862
R36038 VCC.n13273 VCC.n12766 10.5862
R36039 VCC.n13771 VCC.n13353 10.5862
R36040 VCC.n13842 VCC.n13307 10.5862
R36041 VCC.n14326 VCC.n13907 10.5862
R36042 VCC.n14380 VCC.n13873 10.5862
R36043 VCC.n14878 VCC.n14460 10.5862
R36044 VCC.n14949 VCC.n14414 10.5862
R36045 VCC.n15433 VCC.n15014 10.5862
R36046 VCC.n15487 VCC.n14980 10.5862
R36047 VCC.n15985 VCC.n15567 10.5862
R36048 VCC.n16056 VCC.n15521 10.5862
R36049 VCC.n16540 VCC.n16121 10.5862
R36050 VCC.n16594 VCC.n16087 10.5862
R36051 VCC.n17092 VCC.n16674 10.5862
R36052 VCC.n17163 VCC.n16628 10.5862
R36053 VCC.n17460 VCC.n17228 10.5862
R36054 VCC.n17514 VCC.n17194 10.5862
R36055 VCC.n425 VCC.n420 10.5561
R36056 VCC.n977 VCC.n972 10.5561
R36057 VCC.n1535 VCC.n1528 10.5561
R36058 VCC.n2086 VCC.n2081 10.5561
R36059 VCC.n2644 VCC.n2637 10.5561
R36060 VCC.n3195 VCC.n3190 10.5561
R36061 VCC.n3753 VCC.n3746 10.5561
R36062 VCC.n4304 VCC.n4299 10.5561
R36063 VCC.n4862 VCC.n4855 10.5561
R36064 VCC.n5413 VCC.n5408 10.5561
R36065 VCC.n5971 VCC.n5964 10.5561
R36066 VCC.n6522 VCC.n6517 10.5561
R36067 VCC.n7080 VCC.n7073 10.5561
R36068 VCC.n7631 VCC.n7626 10.5561
R36069 VCC.n8189 VCC.n8182 10.5561
R36070 VCC.n8740 VCC.n8735 10.5561
R36071 VCC.n9298 VCC.n9291 10.5561
R36072 VCC.n9849 VCC.n9844 10.5561
R36073 VCC.n10406 VCC.n10399 10.5561
R36074 VCC.n10956 VCC.n10951 10.5561
R36075 VCC.n11513 VCC.n11506 10.5561
R36076 VCC.n12063 VCC.n12058 10.5561
R36077 VCC.n12620 VCC.n12613 10.5561
R36078 VCC.n13170 VCC.n13165 10.5561
R36079 VCC.n13727 VCC.n13720 10.5561
R36080 VCC.n14277 VCC.n14272 10.5561
R36081 VCC.n14834 VCC.n14827 10.5561
R36082 VCC.n15384 VCC.n15379 10.5561
R36083 VCC.n15941 VCC.n15934 10.5561
R36084 VCC.n16491 VCC.n16486 10.5561
R36085 VCC.n17048 VCC.n17041 10.5561
R36086 VCC.n17411 VCC.n17406 10.5561
R36087 VCC.n549 VCC.n548 9.80483
R36088 VCC.n1103 VCC.n1102 9.80483
R36089 VCC.n1657 VCC.n1111 9.80483
R36090 VCC.n2212 VCC.n2211 9.80483
R36091 VCC.n2766 VCC.n2220 9.80483
R36092 VCC.n3321 VCC.n3320 9.80483
R36093 VCC.n3875 VCC.n3329 9.80483
R36094 VCC.n4430 VCC.n4429 9.80483
R36095 VCC.n4984 VCC.n4438 9.80483
R36096 VCC.n5539 VCC.n5538 9.80483
R36097 VCC.n6093 VCC.n5547 9.80483
R36098 VCC.n6648 VCC.n6647 9.80483
R36099 VCC.n7202 VCC.n6656 9.80483
R36100 VCC.n7757 VCC.n7756 9.80483
R36101 VCC.n8311 VCC.n7765 9.80483
R36102 VCC.n8866 VCC.n8865 9.80483
R36103 VCC.n9420 VCC.n8874 9.80483
R36104 VCC.n9975 VCC.n9974 9.80483
R36105 VCC.n10528 VCC.n9982 9.80483
R36106 VCC.n11082 VCC.n11081 9.80483
R36107 VCC.n11635 VCC.n11089 9.80483
R36108 VCC.n12189 VCC.n12188 9.80483
R36109 VCC.n12742 VCC.n12196 9.80483
R36110 VCC.n13296 VCC.n13295 9.80483
R36111 VCC.n13849 VCC.n13303 9.80483
R36112 VCC.n14403 VCC.n14402 9.80483
R36113 VCC.n14956 VCC.n14410 9.80483
R36114 VCC.n15510 VCC.n15509 9.80483
R36115 VCC.n16063 VCC.n15517 9.80483
R36116 VCC.n16617 VCC.n16616 9.80483
R36117 VCC.n17170 VCC.n16624 9.80483
R36118 VCC.n17537 VCC.n17536 9.80483
R36119 VCC.n424 VCC.n65 9.38146
R36120 VCC.n976 VCC.n617 9.38146
R36121 VCC.n2085 VCC.n1726 9.38146
R36122 VCC.n3194 VCC.n2835 9.38146
R36123 VCC.n4303 VCC.n3944 9.38146
R36124 VCC.n5412 VCC.n5053 9.38146
R36125 VCC.n6521 VCC.n6162 9.38146
R36126 VCC.n7630 VCC.n7271 9.38146
R36127 VCC.n8739 VCC.n8380 9.38146
R36128 VCC.n9848 VCC.n9489 9.38146
R36129 VCC.n10955 VCC.n10596 9.38146
R36130 VCC.n12062 VCC.n11703 9.38146
R36131 VCC.n13169 VCC.n12810 9.38146
R36132 VCC.n14276 VCC.n13917 9.38146
R36133 VCC.n15383 VCC.n15024 9.38146
R36134 VCC.n16490 VCC.n16131 9.38146
R36135 VCC.n17410 VCC.n17238 9.38146
R36136 VCC.n1534 VCC.n1174 9.38145
R36137 VCC.n2643 VCC.n2283 9.38145
R36138 VCC.n3752 VCC.n3392 9.38145
R36139 VCC.n4861 VCC.n4501 9.38145
R36140 VCC.n5970 VCC.n5610 9.38145
R36141 VCC.n7079 VCC.n6719 9.38145
R36142 VCC.n8188 VCC.n7828 9.38145
R36143 VCC.n9297 VCC.n8937 9.38145
R36144 VCC.n10405 VCC.n10045 9.38145
R36145 VCC.n11512 VCC.n11152 9.38145
R36146 VCC.n12619 VCC.n12259 9.38145
R36147 VCC.n13726 VCC.n13366 9.38145
R36148 VCC.n14833 VCC.n14473 9.38145
R36149 VCC.n15940 VCC.n15580 9.38145
R36150 VCC.n17047 VCC.n16687 9.38145
R36151 VCC.n233 VCC.n232 9.3005
R36152 VCC.n202 VCC.n201 9.3005
R36153 VCC.n298 VCC.n297 9.3005
R36154 VCC.n273 VCC.n272 9.3005
R36155 VCC.n161 VCC.n160 9.3005
R36156 VCC.n162 VCC.n156 9.3005
R36157 VCC.n151 VCC.n150 9.3005
R36158 VCC.n152 VCC.n151 9.3005
R36159 VCC.n267 VCC.n152 9.3005
R36160 VCC.n145 VCC.n144 9.3005
R36161 VCC.n287 VCC.n134 9.3005
R36162 VCC.n288 VCC.n287 9.3005
R36163 VCC.n289 VCC.n288 9.3005
R36164 VCC.n139 VCC.n137 9.3005
R36165 VCC.n295 VCC.n294 9.3005
R36166 VCC.n177 VCC.n176 9.3005
R36167 VCC.n214 VCC.n213 9.3005
R36168 VCC.n213 VCC.n212 9.3005
R36169 VCC.n212 VCC.n211 9.3005
R36170 VCC.n196 VCC.n195 9.3005
R36171 VCC.n223 VCC.n222 9.3005
R36172 VCC.n223 VCC.n179 9.3005
R36173 VCC.n227 VCC.n179 9.3005
R36174 VCC.n170 VCC.n169 9.3005
R36175 VCC.n169 VCC.n154 9.3005
R36176 VCC.n154 VCC.n153 9.3005
R36177 VCC.n248 VCC.n168 9.3005
R36178 VCC.n250 VCC.n249 9.3005
R36179 VCC.n357 VCC.n356 9.3005
R36180 VCC.n327 VCC.n326 9.3005
R36181 VCC.n433 VCC.n432 9.3005
R36182 VCC.n400 VCC.n399 9.3005
R36183 VCC.n389 VCC.n95 9.3005
R36184 VCC.n388 VCC.n387 9.3005
R36185 VCC.n85 VCC.n84 9.3005
R36186 VCC.n78 VCC.n76 9.3005
R36187 VCC.n111 VCC.n110 9.3005
R36188 VCC.n325 VCC.n320 9.3005
R36189 VCC.n365 VCC.n105 9.3005
R36190 VCC.n98 VCC.n97 9.3005
R36191 VCC.n392 VCC.n90 9.3005
R36192 VCC.n393 VCC.n392 9.3005
R36193 VCC.n394 VCC.n393 9.3005
R36194 VCC.n413 VCC.n73 9.3005
R36195 VCC.n413 VCC.n83 9.3005
R36196 VCC.n83 VCC.n82 9.3005
R36197 VCC.n430 VCC.n68 9.3005
R36198 VCC.n430 VCC.n429 9.3005
R36199 VCC.n429 VCC.n428 9.3005
R36200 VCC.n333 VCC.n332 9.3005
R36201 VCC.n334 VCC.n333 9.3005
R36202 VCC.n335 VCC.n334 9.3005
R36203 VCC.n342 VCC.n341 9.3005
R36204 VCC.n341 VCC.n109 9.3005
R36205 VCC.n109 VCC.n108 9.3005
R36206 VCC.n364 VCC.n104 9.3005
R36207 VCC.n364 VCC.n363 9.3005
R36208 VCC.n363 VCC.n362 9.3005
R36209 VCC.n477 VCC.n476 9.3005
R36210 VCC.n523 VCC.n522 9.3005
R36211 VCC.n524 VCC.n523 9.3005
R36212 VCC.n525 VCC.n524 9.3005
R36213 VCC.n8 VCC.n7 9.3005
R36214 VCC.n516 VCC.n515 9.3005
R36215 VCC.n544 VCC.n543 9.3005
R36216 VCC.n532 VCC.n531 9.3005
R36217 VCC.n531 VCC.n6 9.3005
R36218 VCC.n6 VCC.n5 9.3005
R36219 VCC.n490 VCC.n489 9.3005
R36220 VCC.n490 VCC.n42 9.3005
R36221 VCC.n472 VCC.n42 9.3005
R36222 VCC.n469 VCC.n468 9.3005
R36223 VCC.n470 VCC.n469 9.3005
R36224 VCC.n425 VCC.n424 9.3005
R36225 VCC.n785 VCC.n784 9.3005
R36226 VCC.n754 VCC.n753 9.3005
R36227 VCC.n850 VCC.n849 9.3005
R36228 VCC.n825 VCC.n824 9.3005
R36229 VCC.n713 VCC.n712 9.3005
R36230 VCC.n714 VCC.n708 9.3005
R36231 VCC.n703 VCC.n702 9.3005
R36232 VCC.n704 VCC.n703 9.3005
R36233 VCC.n819 VCC.n704 9.3005
R36234 VCC.n697 VCC.n696 9.3005
R36235 VCC.n839 VCC.n686 9.3005
R36236 VCC.n840 VCC.n839 9.3005
R36237 VCC.n841 VCC.n840 9.3005
R36238 VCC.n691 VCC.n689 9.3005
R36239 VCC.n847 VCC.n846 9.3005
R36240 VCC.n729 VCC.n728 9.3005
R36241 VCC.n766 VCC.n765 9.3005
R36242 VCC.n765 VCC.n764 9.3005
R36243 VCC.n764 VCC.n763 9.3005
R36244 VCC.n748 VCC.n747 9.3005
R36245 VCC.n775 VCC.n774 9.3005
R36246 VCC.n775 VCC.n731 9.3005
R36247 VCC.n779 VCC.n731 9.3005
R36248 VCC.n722 VCC.n721 9.3005
R36249 VCC.n721 VCC.n706 9.3005
R36250 VCC.n706 VCC.n705 9.3005
R36251 VCC.n800 VCC.n720 9.3005
R36252 VCC.n802 VCC.n801 9.3005
R36253 VCC.n909 VCC.n908 9.3005
R36254 VCC.n879 VCC.n878 9.3005
R36255 VCC.n985 VCC.n984 9.3005
R36256 VCC.n952 VCC.n951 9.3005
R36257 VCC.n941 VCC.n647 9.3005
R36258 VCC.n940 VCC.n939 9.3005
R36259 VCC.n637 VCC.n636 9.3005
R36260 VCC.n630 VCC.n628 9.3005
R36261 VCC.n663 VCC.n662 9.3005
R36262 VCC.n877 VCC.n872 9.3005
R36263 VCC.n917 VCC.n657 9.3005
R36264 VCC.n650 VCC.n649 9.3005
R36265 VCC.n944 VCC.n642 9.3005
R36266 VCC.n945 VCC.n944 9.3005
R36267 VCC.n946 VCC.n945 9.3005
R36268 VCC.n965 VCC.n625 9.3005
R36269 VCC.n965 VCC.n635 9.3005
R36270 VCC.n635 VCC.n634 9.3005
R36271 VCC.n982 VCC.n620 9.3005
R36272 VCC.n982 VCC.n981 9.3005
R36273 VCC.n981 VCC.n980 9.3005
R36274 VCC.n885 VCC.n884 9.3005
R36275 VCC.n886 VCC.n885 9.3005
R36276 VCC.n887 VCC.n886 9.3005
R36277 VCC.n894 VCC.n893 9.3005
R36278 VCC.n893 VCC.n661 9.3005
R36279 VCC.n661 VCC.n660 9.3005
R36280 VCC.n916 VCC.n656 9.3005
R36281 VCC.n916 VCC.n915 9.3005
R36282 VCC.n915 VCC.n914 9.3005
R36283 VCC.n1075 VCC.n1074 9.3005
R36284 VCC.n1076 VCC.n1075 9.3005
R36285 VCC.n1077 VCC.n1076 9.3005
R36286 VCC.n1021 VCC.n1020 9.3005
R36287 VCC.n1022 VCC.n1021 9.3005
R36288 VCC.n1029 VCC.n1028 9.3005
R36289 VCC.n1042 VCC.n1041 9.3005
R36290 VCC.n1042 VCC.n594 9.3005
R36291 VCC.n1024 VCC.n594 9.3005
R36292 VCC.n1068 VCC.n1067 9.3005
R36293 VCC.n1084 VCC.n1083 9.3005
R36294 VCC.n1083 VCC.n560 9.3005
R36295 VCC.n560 VCC.n559 9.3005
R36296 VCC.n562 VCC.n561 9.3005
R36297 VCC.n1098 VCC.n1097 9.3005
R36298 VCC.n977 VCC.n976 9.3005
R36299 VCC.n1140 VCC.n1139 9.3005
R36300 VCC.n1125 VCC.n1124 9.3005
R36301 VCC.n1123 VCC.n1122 9.3005
R36302 VCC.n1595 VCC.n1594 9.3005
R36303 VCC.n1588 VCC.n1587 9.3005
R36304 VCC.n1587 VCC.n1586 9.3005
R36305 VCC.n1586 VCC.n1585 9.3005
R36306 VCC.n1648 VCC.n1647 9.3005
R36307 VCC.n1648 VCC.n1113 9.3005
R36308 VCC.n1652 VCC.n1113 9.3005
R36309 VCC.n1624 VCC.n1623 9.3005
R36310 VCC.n1623 VCC.n1622 9.3005
R36311 VCC.n1622 VCC.n1621 9.3005
R36312 VCC.n1577 VCC.n1164 9.3005
R36313 VCC.n1164 VCC.n1163 9.3005
R36314 VCC.n1535 VCC.n1534 9.3005
R36315 VCC.n1543 VCC.n1542 9.3005
R36316 VCC.n1509 VCC.n1508 9.3005
R36317 VCC.n1498 VCC.n1204 9.3005
R36318 VCC.n1207 VCC.n1206 9.3005
R36319 VCC.n1451 VCC.n1450 9.3005
R36320 VCC.n1450 VCC.n1218 9.3005
R36321 VCC.n1218 VCC.n1217 9.3005
R36322 VCC.n1220 VCC.n1219 9.3005
R36323 VCC.n1466 VCC.n1465 9.3005
R36324 VCC.n1473 VCC.n1213 9.3005
R36325 VCC.n1473 VCC.n1472 9.3005
R36326 VCC.n1472 VCC.n1471 9.3005
R36327 VCC.n1474 VCC.n1214 9.3005
R36328 VCC.n1497 VCC.n1496 9.3005
R36329 VCC.n1501 VCC.n1199 9.3005
R36330 VCC.n1502 VCC.n1501 9.3005
R36331 VCC.n1503 VCC.n1502 9.3005
R36332 VCC.n1194 VCC.n1193 9.3005
R36333 VCC.n1522 VCC.n1182 9.3005
R36334 VCC.n1522 VCC.n1192 9.3005
R36335 VCC.n1192 VCC.n1191 9.3005
R36336 VCC.n1187 VCC.n1185 9.3005
R36337 VCC.n1540 VCC.n1177 9.3005
R36338 VCC.n1540 VCC.n1539 9.3005
R36339 VCC.n1539 VCC.n1538 9.3005
R36340 VCC.n1442 VCC.n1441 9.3005
R36341 VCC.n1443 VCC.n1442 9.3005
R36342 VCC.n1444 VCC.n1443 9.3005
R36343 VCC.n1434 VCC.n1430 9.3005
R36344 VCC.n1436 VCC.n1435 9.3005
R36345 VCC.n1408 VCC.n1407 9.3005
R36346 VCC.n1383 VCC.n1382 9.3005
R36347 VCC.n1271 VCC.n1270 9.3005
R36348 VCC.n1360 VCC.n1359 9.3005
R36349 VCC.n1333 VCC.n1332 9.3005
R36350 VCC.n1333 VCC.n1289 9.3005
R36351 VCC.n1337 VCC.n1289 9.3005
R36352 VCC.n1287 VCC.n1286 9.3005
R36353 VCC.n1343 VCC.n1342 9.3005
R36354 VCC.n1280 VCC.n1279 9.3005
R36355 VCC.n1279 VCC.n1264 9.3005
R36356 VCC.n1264 VCC.n1263 9.3005
R36357 VCC.n1358 VCC.n1278 9.3005
R36358 VCC.n1272 VCC.n1266 9.3005
R36359 VCC.n1261 VCC.n1260 9.3005
R36360 VCC.n1262 VCC.n1261 9.3005
R36361 VCC.n1377 VCC.n1262 9.3005
R36362 VCC.n1255 VCC.n1254 9.3005
R36363 VCC.n1397 VCC.n1244 9.3005
R36364 VCC.n1398 VCC.n1397 9.3005
R36365 VCC.n1399 VCC.n1398 9.3005
R36366 VCC.n1249 VCC.n1247 9.3005
R36367 VCC.n1405 VCC.n1404 9.3005
R36368 VCC.n1324 VCC.n1323 9.3005
R36369 VCC.n1323 VCC.n1322 9.3005
R36370 VCC.n1322 VCC.n1321 9.3005
R36371 VCC.n1306 VCC.n1305 9.3005
R36372 VCC.n1312 VCC.n1311 9.3005
R36373 VCC.n1894 VCC.n1893 9.3005
R36374 VCC.n1863 VCC.n1862 9.3005
R36375 VCC.n1959 VCC.n1958 9.3005
R36376 VCC.n1934 VCC.n1933 9.3005
R36377 VCC.n1822 VCC.n1821 9.3005
R36378 VCC.n1823 VCC.n1817 9.3005
R36379 VCC.n1812 VCC.n1811 9.3005
R36380 VCC.n1813 VCC.n1812 9.3005
R36381 VCC.n1928 VCC.n1813 9.3005
R36382 VCC.n1806 VCC.n1805 9.3005
R36383 VCC.n1948 VCC.n1795 9.3005
R36384 VCC.n1949 VCC.n1948 9.3005
R36385 VCC.n1950 VCC.n1949 9.3005
R36386 VCC.n1800 VCC.n1798 9.3005
R36387 VCC.n1956 VCC.n1955 9.3005
R36388 VCC.n1838 VCC.n1837 9.3005
R36389 VCC.n1875 VCC.n1874 9.3005
R36390 VCC.n1874 VCC.n1873 9.3005
R36391 VCC.n1873 VCC.n1872 9.3005
R36392 VCC.n1857 VCC.n1856 9.3005
R36393 VCC.n1884 VCC.n1883 9.3005
R36394 VCC.n1884 VCC.n1840 9.3005
R36395 VCC.n1888 VCC.n1840 9.3005
R36396 VCC.n1831 VCC.n1830 9.3005
R36397 VCC.n1830 VCC.n1815 9.3005
R36398 VCC.n1815 VCC.n1814 9.3005
R36399 VCC.n1909 VCC.n1829 9.3005
R36400 VCC.n1911 VCC.n1910 9.3005
R36401 VCC.n2018 VCC.n2017 9.3005
R36402 VCC.n1988 VCC.n1987 9.3005
R36403 VCC.n2094 VCC.n2093 9.3005
R36404 VCC.n2061 VCC.n2060 9.3005
R36405 VCC.n2050 VCC.n1756 9.3005
R36406 VCC.n2049 VCC.n2048 9.3005
R36407 VCC.n1746 VCC.n1745 9.3005
R36408 VCC.n1739 VCC.n1737 9.3005
R36409 VCC.n1772 VCC.n1771 9.3005
R36410 VCC.n1986 VCC.n1981 9.3005
R36411 VCC.n2026 VCC.n1766 9.3005
R36412 VCC.n1759 VCC.n1758 9.3005
R36413 VCC.n2053 VCC.n1751 9.3005
R36414 VCC.n2054 VCC.n2053 9.3005
R36415 VCC.n2055 VCC.n2054 9.3005
R36416 VCC.n2074 VCC.n1734 9.3005
R36417 VCC.n2074 VCC.n1744 9.3005
R36418 VCC.n1744 VCC.n1743 9.3005
R36419 VCC.n2091 VCC.n1729 9.3005
R36420 VCC.n2091 VCC.n2090 9.3005
R36421 VCC.n2090 VCC.n2089 9.3005
R36422 VCC.n1994 VCC.n1993 9.3005
R36423 VCC.n1995 VCC.n1994 9.3005
R36424 VCC.n1996 VCC.n1995 9.3005
R36425 VCC.n2003 VCC.n2002 9.3005
R36426 VCC.n2002 VCC.n1770 9.3005
R36427 VCC.n1770 VCC.n1769 9.3005
R36428 VCC.n2025 VCC.n1765 9.3005
R36429 VCC.n2025 VCC.n2024 9.3005
R36430 VCC.n2024 VCC.n2023 9.3005
R36431 VCC.n2184 VCC.n2183 9.3005
R36432 VCC.n2185 VCC.n2184 9.3005
R36433 VCC.n2186 VCC.n2185 9.3005
R36434 VCC.n2130 VCC.n2129 9.3005
R36435 VCC.n2131 VCC.n2130 9.3005
R36436 VCC.n2138 VCC.n2137 9.3005
R36437 VCC.n2151 VCC.n2150 9.3005
R36438 VCC.n2151 VCC.n1703 9.3005
R36439 VCC.n2133 VCC.n1703 9.3005
R36440 VCC.n2177 VCC.n2176 9.3005
R36441 VCC.n2193 VCC.n2192 9.3005
R36442 VCC.n2192 VCC.n1669 9.3005
R36443 VCC.n1669 VCC.n1668 9.3005
R36444 VCC.n1671 VCC.n1670 9.3005
R36445 VCC.n2207 VCC.n2206 9.3005
R36446 VCC.n2086 VCC.n2085 9.3005
R36447 VCC.n2249 VCC.n2248 9.3005
R36448 VCC.n2234 VCC.n2233 9.3005
R36449 VCC.n2232 VCC.n2231 9.3005
R36450 VCC.n2704 VCC.n2703 9.3005
R36451 VCC.n2697 VCC.n2696 9.3005
R36452 VCC.n2696 VCC.n2695 9.3005
R36453 VCC.n2695 VCC.n2694 9.3005
R36454 VCC.n2757 VCC.n2756 9.3005
R36455 VCC.n2757 VCC.n2222 9.3005
R36456 VCC.n2761 VCC.n2222 9.3005
R36457 VCC.n2733 VCC.n2732 9.3005
R36458 VCC.n2732 VCC.n2731 9.3005
R36459 VCC.n2731 VCC.n2730 9.3005
R36460 VCC.n2686 VCC.n2273 9.3005
R36461 VCC.n2273 VCC.n2272 9.3005
R36462 VCC.n2644 VCC.n2643 9.3005
R36463 VCC.n2652 VCC.n2651 9.3005
R36464 VCC.n2618 VCC.n2617 9.3005
R36465 VCC.n2607 VCC.n2313 9.3005
R36466 VCC.n2316 VCC.n2315 9.3005
R36467 VCC.n2560 VCC.n2559 9.3005
R36468 VCC.n2559 VCC.n2327 9.3005
R36469 VCC.n2327 VCC.n2326 9.3005
R36470 VCC.n2329 VCC.n2328 9.3005
R36471 VCC.n2575 VCC.n2574 9.3005
R36472 VCC.n2582 VCC.n2322 9.3005
R36473 VCC.n2582 VCC.n2581 9.3005
R36474 VCC.n2581 VCC.n2580 9.3005
R36475 VCC.n2583 VCC.n2323 9.3005
R36476 VCC.n2606 VCC.n2605 9.3005
R36477 VCC.n2610 VCC.n2308 9.3005
R36478 VCC.n2611 VCC.n2610 9.3005
R36479 VCC.n2612 VCC.n2611 9.3005
R36480 VCC.n2303 VCC.n2302 9.3005
R36481 VCC.n2631 VCC.n2291 9.3005
R36482 VCC.n2631 VCC.n2301 9.3005
R36483 VCC.n2301 VCC.n2300 9.3005
R36484 VCC.n2296 VCC.n2294 9.3005
R36485 VCC.n2649 VCC.n2286 9.3005
R36486 VCC.n2649 VCC.n2648 9.3005
R36487 VCC.n2648 VCC.n2647 9.3005
R36488 VCC.n2551 VCC.n2550 9.3005
R36489 VCC.n2552 VCC.n2551 9.3005
R36490 VCC.n2553 VCC.n2552 9.3005
R36491 VCC.n2543 VCC.n2539 9.3005
R36492 VCC.n2545 VCC.n2544 9.3005
R36493 VCC.n2517 VCC.n2516 9.3005
R36494 VCC.n2492 VCC.n2491 9.3005
R36495 VCC.n2380 VCC.n2379 9.3005
R36496 VCC.n2469 VCC.n2468 9.3005
R36497 VCC.n2442 VCC.n2441 9.3005
R36498 VCC.n2442 VCC.n2398 9.3005
R36499 VCC.n2446 VCC.n2398 9.3005
R36500 VCC.n2396 VCC.n2395 9.3005
R36501 VCC.n2452 VCC.n2451 9.3005
R36502 VCC.n2389 VCC.n2388 9.3005
R36503 VCC.n2388 VCC.n2373 9.3005
R36504 VCC.n2373 VCC.n2372 9.3005
R36505 VCC.n2467 VCC.n2387 9.3005
R36506 VCC.n2381 VCC.n2375 9.3005
R36507 VCC.n2370 VCC.n2369 9.3005
R36508 VCC.n2371 VCC.n2370 9.3005
R36509 VCC.n2486 VCC.n2371 9.3005
R36510 VCC.n2364 VCC.n2363 9.3005
R36511 VCC.n2506 VCC.n2353 9.3005
R36512 VCC.n2507 VCC.n2506 9.3005
R36513 VCC.n2508 VCC.n2507 9.3005
R36514 VCC.n2358 VCC.n2356 9.3005
R36515 VCC.n2514 VCC.n2513 9.3005
R36516 VCC.n2433 VCC.n2432 9.3005
R36517 VCC.n2432 VCC.n2431 9.3005
R36518 VCC.n2431 VCC.n2430 9.3005
R36519 VCC.n2415 VCC.n2414 9.3005
R36520 VCC.n2421 VCC.n2420 9.3005
R36521 VCC.n3003 VCC.n3002 9.3005
R36522 VCC.n2972 VCC.n2971 9.3005
R36523 VCC.n3068 VCC.n3067 9.3005
R36524 VCC.n3043 VCC.n3042 9.3005
R36525 VCC.n2931 VCC.n2930 9.3005
R36526 VCC.n2932 VCC.n2926 9.3005
R36527 VCC.n2921 VCC.n2920 9.3005
R36528 VCC.n2922 VCC.n2921 9.3005
R36529 VCC.n3037 VCC.n2922 9.3005
R36530 VCC.n2915 VCC.n2914 9.3005
R36531 VCC.n3057 VCC.n2904 9.3005
R36532 VCC.n3058 VCC.n3057 9.3005
R36533 VCC.n3059 VCC.n3058 9.3005
R36534 VCC.n2909 VCC.n2907 9.3005
R36535 VCC.n3065 VCC.n3064 9.3005
R36536 VCC.n2947 VCC.n2946 9.3005
R36537 VCC.n2984 VCC.n2983 9.3005
R36538 VCC.n2983 VCC.n2982 9.3005
R36539 VCC.n2982 VCC.n2981 9.3005
R36540 VCC.n2966 VCC.n2965 9.3005
R36541 VCC.n2993 VCC.n2992 9.3005
R36542 VCC.n2993 VCC.n2949 9.3005
R36543 VCC.n2997 VCC.n2949 9.3005
R36544 VCC.n2940 VCC.n2939 9.3005
R36545 VCC.n2939 VCC.n2924 9.3005
R36546 VCC.n2924 VCC.n2923 9.3005
R36547 VCC.n3018 VCC.n2938 9.3005
R36548 VCC.n3020 VCC.n3019 9.3005
R36549 VCC.n3127 VCC.n3126 9.3005
R36550 VCC.n3097 VCC.n3096 9.3005
R36551 VCC.n3203 VCC.n3202 9.3005
R36552 VCC.n3170 VCC.n3169 9.3005
R36553 VCC.n3159 VCC.n2865 9.3005
R36554 VCC.n3158 VCC.n3157 9.3005
R36555 VCC.n2855 VCC.n2854 9.3005
R36556 VCC.n2848 VCC.n2846 9.3005
R36557 VCC.n2881 VCC.n2880 9.3005
R36558 VCC.n3095 VCC.n3090 9.3005
R36559 VCC.n3135 VCC.n2875 9.3005
R36560 VCC.n2868 VCC.n2867 9.3005
R36561 VCC.n3162 VCC.n2860 9.3005
R36562 VCC.n3163 VCC.n3162 9.3005
R36563 VCC.n3164 VCC.n3163 9.3005
R36564 VCC.n3183 VCC.n2843 9.3005
R36565 VCC.n3183 VCC.n2853 9.3005
R36566 VCC.n2853 VCC.n2852 9.3005
R36567 VCC.n3200 VCC.n2838 9.3005
R36568 VCC.n3200 VCC.n3199 9.3005
R36569 VCC.n3199 VCC.n3198 9.3005
R36570 VCC.n3103 VCC.n3102 9.3005
R36571 VCC.n3104 VCC.n3103 9.3005
R36572 VCC.n3105 VCC.n3104 9.3005
R36573 VCC.n3112 VCC.n3111 9.3005
R36574 VCC.n3111 VCC.n2879 9.3005
R36575 VCC.n2879 VCC.n2878 9.3005
R36576 VCC.n3134 VCC.n2874 9.3005
R36577 VCC.n3134 VCC.n3133 9.3005
R36578 VCC.n3133 VCC.n3132 9.3005
R36579 VCC.n3293 VCC.n3292 9.3005
R36580 VCC.n3294 VCC.n3293 9.3005
R36581 VCC.n3295 VCC.n3294 9.3005
R36582 VCC.n3239 VCC.n3238 9.3005
R36583 VCC.n3240 VCC.n3239 9.3005
R36584 VCC.n3247 VCC.n3246 9.3005
R36585 VCC.n3260 VCC.n3259 9.3005
R36586 VCC.n3260 VCC.n2812 9.3005
R36587 VCC.n3242 VCC.n2812 9.3005
R36588 VCC.n3286 VCC.n3285 9.3005
R36589 VCC.n3302 VCC.n3301 9.3005
R36590 VCC.n3301 VCC.n2778 9.3005
R36591 VCC.n2778 VCC.n2777 9.3005
R36592 VCC.n2780 VCC.n2779 9.3005
R36593 VCC.n3316 VCC.n3315 9.3005
R36594 VCC.n3195 VCC.n3194 9.3005
R36595 VCC.n3358 VCC.n3357 9.3005
R36596 VCC.n3343 VCC.n3342 9.3005
R36597 VCC.n3341 VCC.n3340 9.3005
R36598 VCC.n3813 VCC.n3812 9.3005
R36599 VCC.n3806 VCC.n3805 9.3005
R36600 VCC.n3805 VCC.n3804 9.3005
R36601 VCC.n3804 VCC.n3803 9.3005
R36602 VCC.n3866 VCC.n3865 9.3005
R36603 VCC.n3866 VCC.n3331 9.3005
R36604 VCC.n3870 VCC.n3331 9.3005
R36605 VCC.n3842 VCC.n3841 9.3005
R36606 VCC.n3841 VCC.n3840 9.3005
R36607 VCC.n3840 VCC.n3839 9.3005
R36608 VCC.n3795 VCC.n3382 9.3005
R36609 VCC.n3382 VCC.n3381 9.3005
R36610 VCC.n3753 VCC.n3752 9.3005
R36611 VCC.n3761 VCC.n3760 9.3005
R36612 VCC.n3727 VCC.n3726 9.3005
R36613 VCC.n3716 VCC.n3422 9.3005
R36614 VCC.n3425 VCC.n3424 9.3005
R36615 VCC.n3669 VCC.n3668 9.3005
R36616 VCC.n3668 VCC.n3436 9.3005
R36617 VCC.n3436 VCC.n3435 9.3005
R36618 VCC.n3438 VCC.n3437 9.3005
R36619 VCC.n3684 VCC.n3683 9.3005
R36620 VCC.n3691 VCC.n3431 9.3005
R36621 VCC.n3691 VCC.n3690 9.3005
R36622 VCC.n3690 VCC.n3689 9.3005
R36623 VCC.n3692 VCC.n3432 9.3005
R36624 VCC.n3715 VCC.n3714 9.3005
R36625 VCC.n3719 VCC.n3417 9.3005
R36626 VCC.n3720 VCC.n3719 9.3005
R36627 VCC.n3721 VCC.n3720 9.3005
R36628 VCC.n3412 VCC.n3411 9.3005
R36629 VCC.n3740 VCC.n3400 9.3005
R36630 VCC.n3740 VCC.n3410 9.3005
R36631 VCC.n3410 VCC.n3409 9.3005
R36632 VCC.n3405 VCC.n3403 9.3005
R36633 VCC.n3758 VCC.n3395 9.3005
R36634 VCC.n3758 VCC.n3757 9.3005
R36635 VCC.n3757 VCC.n3756 9.3005
R36636 VCC.n3660 VCC.n3659 9.3005
R36637 VCC.n3661 VCC.n3660 9.3005
R36638 VCC.n3662 VCC.n3661 9.3005
R36639 VCC.n3652 VCC.n3648 9.3005
R36640 VCC.n3654 VCC.n3653 9.3005
R36641 VCC.n3626 VCC.n3625 9.3005
R36642 VCC.n3601 VCC.n3600 9.3005
R36643 VCC.n3489 VCC.n3488 9.3005
R36644 VCC.n3578 VCC.n3577 9.3005
R36645 VCC.n3551 VCC.n3550 9.3005
R36646 VCC.n3551 VCC.n3507 9.3005
R36647 VCC.n3555 VCC.n3507 9.3005
R36648 VCC.n3505 VCC.n3504 9.3005
R36649 VCC.n3561 VCC.n3560 9.3005
R36650 VCC.n3498 VCC.n3497 9.3005
R36651 VCC.n3497 VCC.n3482 9.3005
R36652 VCC.n3482 VCC.n3481 9.3005
R36653 VCC.n3576 VCC.n3496 9.3005
R36654 VCC.n3490 VCC.n3484 9.3005
R36655 VCC.n3479 VCC.n3478 9.3005
R36656 VCC.n3480 VCC.n3479 9.3005
R36657 VCC.n3595 VCC.n3480 9.3005
R36658 VCC.n3473 VCC.n3472 9.3005
R36659 VCC.n3615 VCC.n3462 9.3005
R36660 VCC.n3616 VCC.n3615 9.3005
R36661 VCC.n3617 VCC.n3616 9.3005
R36662 VCC.n3467 VCC.n3465 9.3005
R36663 VCC.n3623 VCC.n3622 9.3005
R36664 VCC.n3542 VCC.n3541 9.3005
R36665 VCC.n3541 VCC.n3540 9.3005
R36666 VCC.n3540 VCC.n3539 9.3005
R36667 VCC.n3524 VCC.n3523 9.3005
R36668 VCC.n3530 VCC.n3529 9.3005
R36669 VCC.n4112 VCC.n4111 9.3005
R36670 VCC.n4081 VCC.n4080 9.3005
R36671 VCC.n4177 VCC.n4176 9.3005
R36672 VCC.n4152 VCC.n4151 9.3005
R36673 VCC.n4040 VCC.n4039 9.3005
R36674 VCC.n4041 VCC.n4035 9.3005
R36675 VCC.n4030 VCC.n4029 9.3005
R36676 VCC.n4031 VCC.n4030 9.3005
R36677 VCC.n4146 VCC.n4031 9.3005
R36678 VCC.n4024 VCC.n4023 9.3005
R36679 VCC.n4166 VCC.n4013 9.3005
R36680 VCC.n4167 VCC.n4166 9.3005
R36681 VCC.n4168 VCC.n4167 9.3005
R36682 VCC.n4018 VCC.n4016 9.3005
R36683 VCC.n4174 VCC.n4173 9.3005
R36684 VCC.n4056 VCC.n4055 9.3005
R36685 VCC.n4093 VCC.n4092 9.3005
R36686 VCC.n4092 VCC.n4091 9.3005
R36687 VCC.n4091 VCC.n4090 9.3005
R36688 VCC.n4075 VCC.n4074 9.3005
R36689 VCC.n4102 VCC.n4101 9.3005
R36690 VCC.n4102 VCC.n4058 9.3005
R36691 VCC.n4106 VCC.n4058 9.3005
R36692 VCC.n4049 VCC.n4048 9.3005
R36693 VCC.n4048 VCC.n4033 9.3005
R36694 VCC.n4033 VCC.n4032 9.3005
R36695 VCC.n4127 VCC.n4047 9.3005
R36696 VCC.n4129 VCC.n4128 9.3005
R36697 VCC.n4236 VCC.n4235 9.3005
R36698 VCC.n4206 VCC.n4205 9.3005
R36699 VCC.n4312 VCC.n4311 9.3005
R36700 VCC.n4279 VCC.n4278 9.3005
R36701 VCC.n4268 VCC.n3974 9.3005
R36702 VCC.n4267 VCC.n4266 9.3005
R36703 VCC.n3964 VCC.n3963 9.3005
R36704 VCC.n3957 VCC.n3955 9.3005
R36705 VCC.n3990 VCC.n3989 9.3005
R36706 VCC.n4204 VCC.n4199 9.3005
R36707 VCC.n4244 VCC.n3984 9.3005
R36708 VCC.n3977 VCC.n3976 9.3005
R36709 VCC.n4271 VCC.n3969 9.3005
R36710 VCC.n4272 VCC.n4271 9.3005
R36711 VCC.n4273 VCC.n4272 9.3005
R36712 VCC.n4292 VCC.n3952 9.3005
R36713 VCC.n4292 VCC.n3962 9.3005
R36714 VCC.n3962 VCC.n3961 9.3005
R36715 VCC.n4309 VCC.n3947 9.3005
R36716 VCC.n4309 VCC.n4308 9.3005
R36717 VCC.n4308 VCC.n4307 9.3005
R36718 VCC.n4212 VCC.n4211 9.3005
R36719 VCC.n4213 VCC.n4212 9.3005
R36720 VCC.n4214 VCC.n4213 9.3005
R36721 VCC.n4221 VCC.n4220 9.3005
R36722 VCC.n4220 VCC.n3988 9.3005
R36723 VCC.n3988 VCC.n3987 9.3005
R36724 VCC.n4243 VCC.n3983 9.3005
R36725 VCC.n4243 VCC.n4242 9.3005
R36726 VCC.n4242 VCC.n4241 9.3005
R36727 VCC.n4402 VCC.n4401 9.3005
R36728 VCC.n4403 VCC.n4402 9.3005
R36729 VCC.n4404 VCC.n4403 9.3005
R36730 VCC.n4348 VCC.n4347 9.3005
R36731 VCC.n4349 VCC.n4348 9.3005
R36732 VCC.n4356 VCC.n4355 9.3005
R36733 VCC.n4369 VCC.n4368 9.3005
R36734 VCC.n4369 VCC.n3921 9.3005
R36735 VCC.n4351 VCC.n3921 9.3005
R36736 VCC.n4395 VCC.n4394 9.3005
R36737 VCC.n4411 VCC.n4410 9.3005
R36738 VCC.n4410 VCC.n3887 9.3005
R36739 VCC.n3887 VCC.n3886 9.3005
R36740 VCC.n3889 VCC.n3888 9.3005
R36741 VCC.n4425 VCC.n4424 9.3005
R36742 VCC.n4304 VCC.n4303 9.3005
R36743 VCC.n4467 VCC.n4466 9.3005
R36744 VCC.n4452 VCC.n4451 9.3005
R36745 VCC.n4450 VCC.n4449 9.3005
R36746 VCC.n4922 VCC.n4921 9.3005
R36747 VCC.n4915 VCC.n4914 9.3005
R36748 VCC.n4914 VCC.n4913 9.3005
R36749 VCC.n4913 VCC.n4912 9.3005
R36750 VCC.n4975 VCC.n4974 9.3005
R36751 VCC.n4975 VCC.n4440 9.3005
R36752 VCC.n4979 VCC.n4440 9.3005
R36753 VCC.n4951 VCC.n4950 9.3005
R36754 VCC.n4950 VCC.n4949 9.3005
R36755 VCC.n4949 VCC.n4948 9.3005
R36756 VCC.n4904 VCC.n4491 9.3005
R36757 VCC.n4491 VCC.n4490 9.3005
R36758 VCC.n4862 VCC.n4861 9.3005
R36759 VCC.n4870 VCC.n4869 9.3005
R36760 VCC.n4836 VCC.n4835 9.3005
R36761 VCC.n4825 VCC.n4531 9.3005
R36762 VCC.n4534 VCC.n4533 9.3005
R36763 VCC.n4778 VCC.n4777 9.3005
R36764 VCC.n4777 VCC.n4545 9.3005
R36765 VCC.n4545 VCC.n4544 9.3005
R36766 VCC.n4547 VCC.n4546 9.3005
R36767 VCC.n4793 VCC.n4792 9.3005
R36768 VCC.n4800 VCC.n4540 9.3005
R36769 VCC.n4800 VCC.n4799 9.3005
R36770 VCC.n4799 VCC.n4798 9.3005
R36771 VCC.n4801 VCC.n4541 9.3005
R36772 VCC.n4824 VCC.n4823 9.3005
R36773 VCC.n4828 VCC.n4526 9.3005
R36774 VCC.n4829 VCC.n4828 9.3005
R36775 VCC.n4830 VCC.n4829 9.3005
R36776 VCC.n4521 VCC.n4520 9.3005
R36777 VCC.n4849 VCC.n4509 9.3005
R36778 VCC.n4849 VCC.n4519 9.3005
R36779 VCC.n4519 VCC.n4518 9.3005
R36780 VCC.n4514 VCC.n4512 9.3005
R36781 VCC.n4867 VCC.n4504 9.3005
R36782 VCC.n4867 VCC.n4866 9.3005
R36783 VCC.n4866 VCC.n4865 9.3005
R36784 VCC.n4769 VCC.n4768 9.3005
R36785 VCC.n4770 VCC.n4769 9.3005
R36786 VCC.n4771 VCC.n4770 9.3005
R36787 VCC.n4761 VCC.n4757 9.3005
R36788 VCC.n4763 VCC.n4762 9.3005
R36789 VCC.n4735 VCC.n4734 9.3005
R36790 VCC.n4710 VCC.n4709 9.3005
R36791 VCC.n4598 VCC.n4597 9.3005
R36792 VCC.n4687 VCC.n4686 9.3005
R36793 VCC.n4660 VCC.n4659 9.3005
R36794 VCC.n4660 VCC.n4616 9.3005
R36795 VCC.n4664 VCC.n4616 9.3005
R36796 VCC.n4614 VCC.n4613 9.3005
R36797 VCC.n4670 VCC.n4669 9.3005
R36798 VCC.n4607 VCC.n4606 9.3005
R36799 VCC.n4606 VCC.n4591 9.3005
R36800 VCC.n4591 VCC.n4590 9.3005
R36801 VCC.n4685 VCC.n4605 9.3005
R36802 VCC.n4599 VCC.n4593 9.3005
R36803 VCC.n4588 VCC.n4587 9.3005
R36804 VCC.n4589 VCC.n4588 9.3005
R36805 VCC.n4704 VCC.n4589 9.3005
R36806 VCC.n4582 VCC.n4581 9.3005
R36807 VCC.n4724 VCC.n4571 9.3005
R36808 VCC.n4725 VCC.n4724 9.3005
R36809 VCC.n4726 VCC.n4725 9.3005
R36810 VCC.n4576 VCC.n4574 9.3005
R36811 VCC.n4732 VCC.n4731 9.3005
R36812 VCC.n4651 VCC.n4650 9.3005
R36813 VCC.n4650 VCC.n4649 9.3005
R36814 VCC.n4649 VCC.n4648 9.3005
R36815 VCC.n4633 VCC.n4632 9.3005
R36816 VCC.n4639 VCC.n4638 9.3005
R36817 VCC.n5221 VCC.n5220 9.3005
R36818 VCC.n5190 VCC.n5189 9.3005
R36819 VCC.n5286 VCC.n5285 9.3005
R36820 VCC.n5261 VCC.n5260 9.3005
R36821 VCC.n5149 VCC.n5148 9.3005
R36822 VCC.n5150 VCC.n5144 9.3005
R36823 VCC.n5139 VCC.n5138 9.3005
R36824 VCC.n5140 VCC.n5139 9.3005
R36825 VCC.n5255 VCC.n5140 9.3005
R36826 VCC.n5133 VCC.n5132 9.3005
R36827 VCC.n5275 VCC.n5122 9.3005
R36828 VCC.n5276 VCC.n5275 9.3005
R36829 VCC.n5277 VCC.n5276 9.3005
R36830 VCC.n5127 VCC.n5125 9.3005
R36831 VCC.n5283 VCC.n5282 9.3005
R36832 VCC.n5165 VCC.n5164 9.3005
R36833 VCC.n5202 VCC.n5201 9.3005
R36834 VCC.n5201 VCC.n5200 9.3005
R36835 VCC.n5200 VCC.n5199 9.3005
R36836 VCC.n5184 VCC.n5183 9.3005
R36837 VCC.n5211 VCC.n5210 9.3005
R36838 VCC.n5211 VCC.n5167 9.3005
R36839 VCC.n5215 VCC.n5167 9.3005
R36840 VCC.n5158 VCC.n5157 9.3005
R36841 VCC.n5157 VCC.n5142 9.3005
R36842 VCC.n5142 VCC.n5141 9.3005
R36843 VCC.n5236 VCC.n5156 9.3005
R36844 VCC.n5238 VCC.n5237 9.3005
R36845 VCC.n5345 VCC.n5344 9.3005
R36846 VCC.n5315 VCC.n5314 9.3005
R36847 VCC.n5421 VCC.n5420 9.3005
R36848 VCC.n5388 VCC.n5387 9.3005
R36849 VCC.n5377 VCC.n5083 9.3005
R36850 VCC.n5376 VCC.n5375 9.3005
R36851 VCC.n5073 VCC.n5072 9.3005
R36852 VCC.n5066 VCC.n5064 9.3005
R36853 VCC.n5099 VCC.n5098 9.3005
R36854 VCC.n5313 VCC.n5308 9.3005
R36855 VCC.n5353 VCC.n5093 9.3005
R36856 VCC.n5086 VCC.n5085 9.3005
R36857 VCC.n5380 VCC.n5078 9.3005
R36858 VCC.n5381 VCC.n5380 9.3005
R36859 VCC.n5382 VCC.n5381 9.3005
R36860 VCC.n5401 VCC.n5061 9.3005
R36861 VCC.n5401 VCC.n5071 9.3005
R36862 VCC.n5071 VCC.n5070 9.3005
R36863 VCC.n5418 VCC.n5056 9.3005
R36864 VCC.n5418 VCC.n5417 9.3005
R36865 VCC.n5417 VCC.n5416 9.3005
R36866 VCC.n5321 VCC.n5320 9.3005
R36867 VCC.n5322 VCC.n5321 9.3005
R36868 VCC.n5323 VCC.n5322 9.3005
R36869 VCC.n5330 VCC.n5329 9.3005
R36870 VCC.n5329 VCC.n5097 9.3005
R36871 VCC.n5097 VCC.n5096 9.3005
R36872 VCC.n5352 VCC.n5092 9.3005
R36873 VCC.n5352 VCC.n5351 9.3005
R36874 VCC.n5351 VCC.n5350 9.3005
R36875 VCC.n5511 VCC.n5510 9.3005
R36876 VCC.n5512 VCC.n5511 9.3005
R36877 VCC.n5513 VCC.n5512 9.3005
R36878 VCC.n5457 VCC.n5456 9.3005
R36879 VCC.n5458 VCC.n5457 9.3005
R36880 VCC.n5465 VCC.n5464 9.3005
R36881 VCC.n5478 VCC.n5477 9.3005
R36882 VCC.n5478 VCC.n5030 9.3005
R36883 VCC.n5460 VCC.n5030 9.3005
R36884 VCC.n5504 VCC.n5503 9.3005
R36885 VCC.n5520 VCC.n5519 9.3005
R36886 VCC.n5519 VCC.n4996 9.3005
R36887 VCC.n4996 VCC.n4995 9.3005
R36888 VCC.n4998 VCC.n4997 9.3005
R36889 VCC.n5534 VCC.n5533 9.3005
R36890 VCC.n5413 VCC.n5412 9.3005
R36891 VCC.n5576 VCC.n5575 9.3005
R36892 VCC.n5561 VCC.n5560 9.3005
R36893 VCC.n5559 VCC.n5558 9.3005
R36894 VCC.n6031 VCC.n6030 9.3005
R36895 VCC.n6024 VCC.n6023 9.3005
R36896 VCC.n6023 VCC.n6022 9.3005
R36897 VCC.n6022 VCC.n6021 9.3005
R36898 VCC.n6084 VCC.n6083 9.3005
R36899 VCC.n6084 VCC.n5549 9.3005
R36900 VCC.n6088 VCC.n5549 9.3005
R36901 VCC.n6060 VCC.n6059 9.3005
R36902 VCC.n6059 VCC.n6058 9.3005
R36903 VCC.n6058 VCC.n6057 9.3005
R36904 VCC.n6013 VCC.n5600 9.3005
R36905 VCC.n5600 VCC.n5599 9.3005
R36906 VCC.n5971 VCC.n5970 9.3005
R36907 VCC.n5979 VCC.n5978 9.3005
R36908 VCC.n5945 VCC.n5944 9.3005
R36909 VCC.n5934 VCC.n5640 9.3005
R36910 VCC.n5643 VCC.n5642 9.3005
R36911 VCC.n5887 VCC.n5886 9.3005
R36912 VCC.n5886 VCC.n5654 9.3005
R36913 VCC.n5654 VCC.n5653 9.3005
R36914 VCC.n5656 VCC.n5655 9.3005
R36915 VCC.n5902 VCC.n5901 9.3005
R36916 VCC.n5909 VCC.n5649 9.3005
R36917 VCC.n5909 VCC.n5908 9.3005
R36918 VCC.n5908 VCC.n5907 9.3005
R36919 VCC.n5910 VCC.n5650 9.3005
R36920 VCC.n5933 VCC.n5932 9.3005
R36921 VCC.n5937 VCC.n5635 9.3005
R36922 VCC.n5938 VCC.n5937 9.3005
R36923 VCC.n5939 VCC.n5938 9.3005
R36924 VCC.n5630 VCC.n5629 9.3005
R36925 VCC.n5958 VCC.n5618 9.3005
R36926 VCC.n5958 VCC.n5628 9.3005
R36927 VCC.n5628 VCC.n5627 9.3005
R36928 VCC.n5623 VCC.n5621 9.3005
R36929 VCC.n5976 VCC.n5613 9.3005
R36930 VCC.n5976 VCC.n5975 9.3005
R36931 VCC.n5975 VCC.n5974 9.3005
R36932 VCC.n5878 VCC.n5877 9.3005
R36933 VCC.n5879 VCC.n5878 9.3005
R36934 VCC.n5880 VCC.n5879 9.3005
R36935 VCC.n5870 VCC.n5866 9.3005
R36936 VCC.n5872 VCC.n5871 9.3005
R36937 VCC.n5844 VCC.n5843 9.3005
R36938 VCC.n5819 VCC.n5818 9.3005
R36939 VCC.n5707 VCC.n5706 9.3005
R36940 VCC.n5796 VCC.n5795 9.3005
R36941 VCC.n5769 VCC.n5768 9.3005
R36942 VCC.n5769 VCC.n5725 9.3005
R36943 VCC.n5773 VCC.n5725 9.3005
R36944 VCC.n5723 VCC.n5722 9.3005
R36945 VCC.n5779 VCC.n5778 9.3005
R36946 VCC.n5716 VCC.n5715 9.3005
R36947 VCC.n5715 VCC.n5700 9.3005
R36948 VCC.n5700 VCC.n5699 9.3005
R36949 VCC.n5794 VCC.n5714 9.3005
R36950 VCC.n5708 VCC.n5702 9.3005
R36951 VCC.n5697 VCC.n5696 9.3005
R36952 VCC.n5698 VCC.n5697 9.3005
R36953 VCC.n5813 VCC.n5698 9.3005
R36954 VCC.n5691 VCC.n5690 9.3005
R36955 VCC.n5833 VCC.n5680 9.3005
R36956 VCC.n5834 VCC.n5833 9.3005
R36957 VCC.n5835 VCC.n5834 9.3005
R36958 VCC.n5685 VCC.n5683 9.3005
R36959 VCC.n5841 VCC.n5840 9.3005
R36960 VCC.n5760 VCC.n5759 9.3005
R36961 VCC.n5759 VCC.n5758 9.3005
R36962 VCC.n5758 VCC.n5757 9.3005
R36963 VCC.n5742 VCC.n5741 9.3005
R36964 VCC.n5748 VCC.n5747 9.3005
R36965 VCC.n6330 VCC.n6329 9.3005
R36966 VCC.n6299 VCC.n6298 9.3005
R36967 VCC.n6395 VCC.n6394 9.3005
R36968 VCC.n6370 VCC.n6369 9.3005
R36969 VCC.n6258 VCC.n6257 9.3005
R36970 VCC.n6259 VCC.n6253 9.3005
R36971 VCC.n6248 VCC.n6247 9.3005
R36972 VCC.n6249 VCC.n6248 9.3005
R36973 VCC.n6364 VCC.n6249 9.3005
R36974 VCC.n6242 VCC.n6241 9.3005
R36975 VCC.n6384 VCC.n6231 9.3005
R36976 VCC.n6385 VCC.n6384 9.3005
R36977 VCC.n6386 VCC.n6385 9.3005
R36978 VCC.n6236 VCC.n6234 9.3005
R36979 VCC.n6392 VCC.n6391 9.3005
R36980 VCC.n6274 VCC.n6273 9.3005
R36981 VCC.n6311 VCC.n6310 9.3005
R36982 VCC.n6310 VCC.n6309 9.3005
R36983 VCC.n6309 VCC.n6308 9.3005
R36984 VCC.n6293 VCC.n6292 9.3005
R36985 VCC.n6320 VCC.n6319 9.3005
R36986 VCC.n6320 VCC.n6276 9.3005
R36987 VCC.n6324 VCC.n6276 9.3005
R36988 VCC.n6267 VCC.n6266 9.3005
R36989 VCC.n6266 VCC.n6251 9.3005
R36990 VCC.n6251 VCC.n6250 9.3005
R36991 VCC.n6345 VCC.n6265 9.3005
R36992 VCC.n6347 VCC.n6346 9.3005
R36993 VCC.n6454 VCC.n6453 9.3005
R36994 VCC.n6424 VCC.n6423 9.3005
R36995 VCC.n6530 VCC.n6529 9.3005
R36996 VCC.n6497 VCC.n6496 9.3005
R36997 VCC.n6486 VCC.n6192 9.3005
R36998 VCC.n6485 VCC.n6484 9.3005
R36999 VCC.n6182 VCC.n6181 9.3005
R37000 VCC.n6175 VCC.n6173 9.3005
R37001 VCC.n6208 VCC.n6207 9.3005
R37002 VCC.n6422 VCC.n6417 9.3005
R37003 VCC.n6462 VCC.n6202 9.3005
R37004 VCC.n6195 VCC.n6194 9.3005
R37005 VCC.n6489 VCC.n6187 9.3005
R37006 VCC.n6490 VCC.n6489 9.3005
R37007 VCC.n6491 VCC.n6490 9.3005
R37008 VCC.n6510 VCC.n6170 9.3005
R37009 VCC.n6510 VCC.n6180 9.3005
R37010 VCC.n6180 VCC.n6179 9.3005
R37011 VCC.n6527 VCC.n6165 9.3005
R37012 VCC.n6527 VCC.n6526 9.3005
R37013 VCC.n6526 VCC.n6525 9.3005
R37014 VCC.n6430 VCC.n6429 9.3005
R37015 VCC.n6431 VCC.n6430 9.3005
R37016 VCC.n6432 VCC.n6431 9.3005
R37017 VCC.n6439 VCC.n6438 9.3005
R37018 VCC.n6438 VCC.n6206 9.3005
R37019 VCC.n6206 VCC.n6205 9.3005
R37020 VCC.n6461 VCC.n6201 9.3005
R37021 VCC.n6461 VCC.n6460 9.3005
R37022 VCC.n6460 VCC.n6459 9.3005
R37023 VCC.n6620 VCC.n6619 9.3005
R37024 VCC.n6621 VCC.n6620 9.3005
R37025 VCC.n6622 VCC.n6621 9.3005
R37026 VCC.n6566 VCC.n6565 9.3005
R37027 VCC.n6567 VCC.n6566 9.3005
R37028 VCC.n6574 VCC.n6573 9.3005
R37029 VCC.n6587 VCC.n6586 9.3005
R37030 VCC.n6587 VCC.n6139 9.3005
R37031 VCC.n6569 VCC.n6139 9.3005
R37032 VCC.n6613 VCC.n6612 9.3005
R37033 VCC.n6629 VCC.n6628 9.3005
R37034 VCC.n6628 VCC.n6105 9.3005
R37035 VCC.n6105 VCC.n6104 9.3005
R37036 VCC.n6107 VCC.n6106 9.3005
R37037 VCC.n6643 VCC.n6642 9.3005
R37038 VCC.n6522 VCC.n6521 9.3005
R37039 VCC.n6685 VCC.n6684 9.3005
R37040 VCC.n6670 VCC.n6669 9.3005
R37041 VCC.n6668 VCC.n6667 9.3005
R37042 VCC.n7140 VCC.n7139 9.3005
R37043 VCC.n7133 VCC.n7132 9.3005
R37044 VCC.n7132 VCC.n7131 9.3005
R37045 VCC.n7131 VCC.n7130 9.3005
R37046 VCC.n7193 VCC.n7192 9.3005
R37047 VCC.n7193 VCC.n6658 9.3005
R37048 VCC.n7197 VCC.n6658 9.3005
R37049 VCC.n7169 VCC.n7168 9.3005
R37050 VCC.n7168 VCC.n7167 9.3005
R37051 VCC.n7167 VCC.n7166 9.3005
R37052 VCC.n7122 VCC.n6709 9.3005
R37053 VCC.n6709 VCC.n6708 9.3005
R37054 VCC.n7080 VCC.n7079 9.3005
R37055 VCC.n7088 VCC.n7087 9.3005
R37056 VCC.n7054 VCC.n7053 9.3005
R37057 VCC.n7043 VCC.n6749 9.3005
R37058 VCC.n6752 VCC.n6751 9.3005
R37059 VCC.n6996 VCC.n6995 9.3005
R37060 VCC.n6995 VCC.n6763 9.3005
R37061 VCC.n6763 VCC.n6762 9.3005
R37062 VCC.n6765 VCC.n6764 9.3005
R37063 VCC.n7011 VCC.n7010 9.3005
R37064 VCC.n7018 VCC.n6758 9.3005
R37065 VCC.n7018 VCC.n7017 9.3005
R37066 VCC.n7017 VCC.n7016 9.3005
R37067 VCC.n7019 VCC.n6759 9.3005
R37068 VCC.n7042 VCC.n7041 9.3005
R37069 VCC.n7046 VCC.n6744 9.3005
R37070 VCC.n7047 VCC.n7046 9.3005
R37071 VCC.n7048 VCC.n7047 9.3005
R37072 VCC.n6739 VCC.n6738 9.3005
R37073 VCC.n7067 VCC.n6727 9.3005
R37074 VCC.n7067 VCC.n6737 9.3005
R37075 VCC.n6737 VCC.n6736 9.3005
R37076 VCC.n6732 VCC.n6730 9.3005
R37077 VCC.n7085 VCC.n6722 9.3005
R37078 VCC.n7085 VCC.n7084 9.3005
R37079 VCC.n7084 VCC.n7083 9.3005
R37080 VCC.n6987 VCC.n6986 9.3005
R37081 VCC.n6988 VCC.n6987 9.3005
R37082 VCC.n6989 VCC.n6988 9.3005
R37083 VCC.n6979 VCC.n6975 9.3005
R37084 VCC.n6981 VCC.n6980 9.3005
R37085 VCC.n6953 VCC.n6952 9.3005
R37086 VCC.n6928 VCC.n6927 9.3005
R37087 VCC.n6816 VCC.n6815 9.3005
R37088 VCC.n6905 VCC.n6904 9.3005
R37089 VCC.n6878 VCC.n6877 9.3005
R37090 VCC.n6878 VCC.n6834 9.3005
R37091 VCC.n6882 VCC.n6834 9.3005
R37092 VCC.n6832 VCC.n6831 9.3005
R37093 VCC.n6888 VCC.n6887 9.3005
R37094 VCC.n6825 VCC.n6824 9.3005
R37095 VCC.n6824 VCC.n6809 9.3005
R37096 VCC.n6809 VCC.n6808 9.3005
R37097 VCC.n6903 VCC.n6823 9.3005
R37098 VCC.n6817 VCC.n6811 9.3005
R37099 VCC.n6806 VCC.n6805 9.3005
R37100 VCC.n6807 VCC.n6806 9.3005
R37101 VCC.n6922 VCC.n6807 9.3005
R37102 VCC.n6800 VCC.n6799 9.3005
R37103 VCC.n6942 VCC.n6789 9.3005
R37104 VCC.n6943 VCC.n6942 9.3005
R37105 VCC.n6944 VCC.n6943 9.3005
R37106 VCC.n6794 VCC.n6792 9.3005
R37107 VCC.n6950 VCC.n6949 9.3005
R37108 VCC.n6869 VCC.n6868 9.3005
R37109 VCC.n6868 VCC.n6867 9.3005
R37110 VCC.n6867 VCC.n6866 9.3005
R37111 VCC.n6851 VCC.n6850 9.3005
R37112 VCC.n6857 VCC.n6856 9.3005
R37113 VCC.n7439 VCC.n7438 9.3005
R37114 VCC.n7408 VCC.n7407 9.3005
R37115 VCC.n7504 VCC.n7503 9.3005
R37116 VCC.n7479 VCC.n7478 9.3005
R37117 VCC.n7367 VCC.n7366 9.3005
R37118 VCC.n7368 VCC.n7362 9.3005
R37119 VCC.n7357 VCC.n7356 9.3005
R37120 VCC.n7358 VCC.n7357 9.3005
R37121 VCC.n7473 VCC.n7358 9.3005
R37122 VCC.n7351 VCC.n7350 9.3005
R37123 VCC.n7493 VCC.n7340 9.3005
R37124 VCC.n7494 VCC.n7493 9.3005
R37125 VCC.n7495 VCC.n7494 9.3005
R37126 VCC.n7345 VCC.n7343 9.3005
R37127 VCC.n7501 VCC.n7500 9.3005
R37128 VCC.n7383 VCC.n7382 9.3005
R37129 VCC.n7420 VCC.n7419 9.3005
R37130 VCC.n7419 VCC.n7418 9.3005
R37131 VCC.n7418 VCC.n7417 9.3005
R37132 VCC.n7402 VCC.n7401 9.3005
R37133 VCC.n7429 VCC.n7428 9.3005
R37134 VCC.n7429 VCC.n7385 9.3005
R37135 VCC.n7433 VCC.n7385 9.3005
R37136 VCC.n7376 VCC.n7375 9.3005
R37137 VCC.n7375 VCC.n7360 9.3005
R37138 VCC.n7360 VCC.n7359 9.3005
R37139 VCC.n7454 VCC.n7374 9.3005
R37140 VCC.n7456 VCC.n7455 9.3005
R37141 VCC.n7563 VCC.n7562 9.3005
R37142 VCC.n7533 VCC.n7532 9.3005
R37143 VCC.n7639 VCC.n7638 9.3005
R37144 VCC.n7606 VCC.n7605 9.3005
R37145 VCC.n7595 VCC.n7301 9.3005
R37146 VCC.n7594 VCC.n7593 9.3005
R37147 VCC.n7291 VCC.n7290 9.3005
R37148 VCC.n7284 VCC.n7282 9.3005
R37149 VCC.n7317 VCC.n7316 9.3005
R37150 VCC.n7531 VCC.n7526 9.3005
R37151 VCC.n7571 VCC.n7311 9.3005
R37152 VCC.n7304 VCC.n7303 9.3005
R37153 VCC.n7598 VCC.n7296 9.3005
R37154 VCC.n7599 VCC.n7598 9.3005
R37155 VCC.n7600 VCC.n7599 9.3005
R37156 VCC.n7619 VCC.n7279 9.3005
R37157 VCC.n7619 VCC.n7289 9.3005
R37158 VCC.n7289 VCC.n7288 9.3005
R37159 VCC.n7636 VCC.n7274 9.3005
R37160 VCC.n7636 VCC.n7635 9.3005
R37161 VCC.n7635 VCC.n7634 9.3005
R37162 VCC.n7539 VCC.n7538 9.3005
R37163 VCC.n7540 VCC.n7539 9.3005
R37164 VCC.n7541 VCC.n7540 9.3005
R37165 VCC.n7548 VCC.n7547 9.3005
R37166 VCC.n7547 VCC.n7315 9.3005
R37167 VCC.n7315 VCC.n7314 9.3005
R37168 VCC.n7570 VCC.n7310 9.3005
R37169 VCC.n7570 VCC.n7569 9.3005
R37170 VCC.n7569 VCC.n7568 9.3005
R37171 VCC.n7729 VCC.n7728 9.3005
R37172 VCC.n7730 VCC.n7729 9.3005
R37173 VCC.n7731 VCC.n7730 9.3005
R37174 VCC.n7675 VCC.n7674 9.3005
R37175 VCC.n7676 VCC.n7675 9.3005
R37176 VCC.n7683 VCC.n7682 9.3005
R37177 VCC.n7696 VCC.n7695 9.3005
R37178 VCC.n7696 VCC.n7248 9.3005
R37179 VCC.n7678 VCC.n7248 9.3005
R37180 VCC.n7722 VCC.n7721 9.3005
R37181 VCC.n7738 VCC.n7737 9.3005
R37182 VCC.n7737 VCC.n7214 9.3005
R37183 VCC.n7214 VCC.n7213 9.3005
R37184 VCC.n7216 VCC.n7215 9.3005
R37185 VCC.n7752 VCC.n7751 9.3005
R37186 VCC.n7631 VCC.n7630 9.3005
R37187 VCC.n7794 VCC.n7793 9.3005
R37188 VCC.n7779 VCC.n7778 9.3005
R37189 VCC.n7777 VCC.n7776 9.3005
R37190 VCC.n8249 VCC.n8248 9.3005
R37191 VCC.n8242 VCC.n8241 9.3005
R37192 VCC.n8241 VCC.n8240 9.3005
R37193 VCC.n8240 VCC.n8239 9.3005
R37194 VCC.n8302 VCC.n8301 9.3005
R37195 VCC.n8302 VCC.n7767 9.3005
R37196 VCC.n8306 VCC.n7767 9.3005
R37197 VCC.n8278 VCC.n8277 9.3005
R37198 VCC.n8277 VCC.n8276 9.3005
R37199 VCC.n8276 VCC.n8275 9.3005
R37200 VCC.n8231 VCC.n7818 9.3005
R37201 VCC.n7818 VCC.n7817 9.3005
R37202 VCC.n8189 VCC.n8188 9.3005
R37203 VCC.n8197 VCC.n8196 9.3005
R37204 VCC.n8163 VCC.n8162 9.3005
R37205 VCC.n8152 VCC.n7858 9.3005
R37206 VCC.n7861 VCC.n7860 9.3005
R37207 VCC.n8105 VCC.n8104 9.3005
R37208 VCC.n8104 VCC.n7872 9.3005
R37209 VCC.n7872 VCC.n7871 9.3005
R37210 VCC.n7874 VCC.n7873 9.3005
R37211 VCC.n8120 VCC.n8119 9.3005
R37212 VCC.n8127 VCC.n7867 9.3005
R37213 VCC.n8127 VCC.n8126 9.3005
R37214 VCC.n8126 VCC.n8125 9.3005
R37215 VCC.n8128 VCC.n7868 9.3005
R37216 VCC.n8151 VCC.n8150 9.3005
R37217 VCC.n8155 VCC.n7853 9.3005
R37218 VCC.n8156 VCC.n8155 9.3005
R37219 VCC.n8157 VCC.n8156 9.3005
R37220 VCC.n7848 VCC.n7847 9.3005
R37221 VCC.n8176 VCC.n7836 9.3005
R37222 VCC.n8176 VCC.n7846 9.3005
R37223 VCC.n7846 VCC.n7845 9.3005
R37224 VCC.n7841 VCC.n7839 9.3005
R37225 VCC.n8194 VCC.n7831 9.3005
R37226 VCC.n8194 VCC.n8193 9.3005
R37227 VCC.n8193 VCC.n8192 9.3005
R37228 VCC.n8096 VCC.n8095 9.3005
R37229 VCC.n8097 VCC.n8096 9.3005
R37230 VCC.n8098 VCC.n8097 9.3005
R37231 VCC.n8088 VCC.n8084 9.3005
R37232 VCC.n8090 VCC.n8089 9.3005
R37233 VCC.n8062 VCC.n8061 9.3005
R37234 VCC.n8037 VCC.n8036 9.3005
R37235 VCC.n7925 VCC.n7924 9.3005
R37236 VCC.n8014 VCC.n8013 9.3005
R37237 VCC.n7987 VCC.n7986 9.3005
R37238 VCC.n7987 VCC.n7943 9.3005
R37239 VCC.n7991 VCC.n7943 9.3005
R37240 VCC.n7941 VCC.n7940 9.3005
R37241 VCC.n7997 VCC.n7996 9.3005
R37242 VCC.n7934 VCC.n7933 9.3005
R37243 VCC.n7933 VCC.n7918 9.3005
R37244 VCC.n7918 VCC.n7917 9.3005
R37245 VCC.n8012 VCC.n7932 9.3005
R37246 VCC.n7926 VCC.n7920 9.3005
R37247 VCC.n7915 VCC.n7914 9.3005
R37248 VCC.n7916 VCC.n7915 9.3005
R37249 VCC.n8031 VCC.n7916 9.3005
R37250 VCC.n7909 VCC.n7908 9.3005
R37251 VCC.n8051 VCC.n7898 9.3005
R37252 VCC.n8052 VCC.n8051 9.3005
R37253 VCC.n8053 VCC.n8052 9.3005
R37254 VCC.n7903 VCC.n7901 9.3005
R37255 VCC.n8059 VCC.n8058 9.3005
R37256 VCC.n7978 VCC.n7977 9.3005
R37257 VCC.n7977 VCC.n7976 9.3005
R37258 VCC.n7976 VCC.n7975 9.3005
R37259 VCC.n7960 VCC.n7959 9.3005
R37260 VCC.n7966 VCC.n7965 9.3005
R37261 VCC.n8672 VCC.n8671 9.3005
R37262 VCC.n8642 VCC.n8641 9.3005
R37263 VCC.n8748 VCC.n8747 9.3005
R37264 VCC.n8715 VCC.n8714 9.3005
R37265 VCC.n8704 VCC.n8410 9.3005
R37266 VCC.n8703 VCC.n8702 9.3005
R37267 VCC.n8400 VCC.n8399 9.3005
R37268 VCC.n8393 VCC.n8391 9.3005
R37269 VCC.n8426 VCC.n8425 9.3005
R37270 VCC.n8640 VCC.n8635 9.3005
R37271 VCC.n8680 VCC.n8420 9.3005
R37272 VCC.n8413 VCC.n8412 9.3005
R37273 VCC.n8707 VCC.n8405 9.3005
R37274 VCC.n8708 VCC.n8707 9.3005
R37275 VCC.n8709 VCC.n8708 9.3005
R37276 VCC.n8728 VCC.n8388 9.3005
R37277 VCC.n8728 VCC.n8398 9.3005
R37278 VCC.n8398 VCC.n8397 9.3005
R37279 VCC.n8745 VCC.n8383 9.3005
R37280 VCC.n8745 VCC.n8744 9.3005
R37281 VCC.n8744 VCC.n8743 9.3005
R37282 VCC.n8648 VCC.n8647 9.3005
R37283 VCC.n8649 VCC.n8648 9.3005
R37284 VCC.n8650 VCC.n8649 9.3005
R37285 VCC.n8657 VCC.n8656 9.3005
R37286 VCC.n8656 VCC.n8424 9.3005
R37287 VCC.n8424 VCC.n8423 9.3005
R37288 VCC.n8679 VCC.n8419 9.3005
R37289 VCC.n8679 VCC.n8678 9.3005
R37290 VCC.n8678 VCC.n8677 9.3005
R37291 VCC.n8838 VCC.n8837 9.3005
R37292 VCC.n8839 VCC.n8838 9.3005
R37293 VCC.n8840 VCC.n8839 9.3005
R37294 VCC.n8784 VCC.n8783 9.3005
R37295 VCC.n8785 VCC.n8784 9.3005
R37296 VCC.n8792 VCC.n8791 9.3005
R37297 VCC.n8805 VCC.n8804 9.3005
R37298 VCC.n8805 VCC.n8357 9.3005
R37299 VCC.n8787 VCC.n8357 9.3005
R37300 VCC.n8831 VCC.n8830 9.3005
R37301 VCC.n8847 VCC.n8846 9.3005
R37302 VCC.n8846 VCC.n8323 9.3005
R37303 VCC.n8323 VCC.n8322 9.3005
R37304 VCC.n8325 VCC.n8324 9.3005
R37305 VCC.n8861 VCC.n8860 9.3005
R37306 VCC.n8740 VCC.n8739 9.3005
R37307 VCC.n8613 VCC.n8612 9.3005
R37308 VCC.n8588 VCC.n8587 9.3005
R37309 VCC.n8476 VCC.n8475 9.3005
R37310 VCC.n8565 VCC.n8564 9.3005
R37311 VCC.n8538 VCC.n8537 9.3005
R37312 VCC.n8538 VCC.n8494 9.3005
R37313 VCC.n8542 VCC.n8494 9.3005
R37314 VCC.n8492 VCC.n8491 9.3005
R37315 VCC.n8548 VCC.n8547 9.3005
R37316 VCC.n8485 VCC.n8484 9.3005
R37317 VCC.n8484 VCC.n8469 9.3005
R37318 VCC.n8469 VCC.n8468 9.3005
R37319 VCC.n8563 VCC.n8483 9.3005
R37320 VCC.n8477 VCC.n8471 9.3005
R37321 VCC.n8466 VCC.n8465 9.3005
R37322 VCC.n8467 VCC.n8466 9.3005
R37323 VCC.n8582 VCC.n8467 9.3005
R37324 VCC.n8460 VCC.n8459 9.3005
R37325 VCC.n8602 VCC.n8449 9.3005
R37326 VCC.n8603 VCC.n8602 9.3005
R37327 VCC.n8604 VCC.n8603 9.3005
R37328 VCC.n8454 VCC.n8452 9.3005
R37329 VCC.n8610 VCC.n8609 9.3005
R37330 VCC.n8529 VCC.n8528 9.3005
R37331 VCC.n8528 VCC.n8527 9.3005
R37332 VCC.n8527 VCC.n8526 9.3005
R37333 VCC.n8511 VCC.n8510 9.3005
R37334 VCC.n8517 VCC.n8516 9.3005
R37335 VCC.n8903 VCC.n8902 9.3005
R37336 VCC.n8888 VCC.n8887 9.3005
R37337 VCC.n8886 VCC.n8885 9.3005
R37338 VCC.n9358 VCC.n9357 9.3005
R37339 VCC.n9351 VCC.n9350 9.3005
R37340 VCC.n9350 VCC.n9349 9.3005
R37341 VCC.n9349 VCC.n9348 9.3005
R37342 VCC.n9411 VCC.n9410 9.3005
R37343 VCC.n9411 VCC.n8876 9.3005
R37344 VCC.n9415 VCC.n8876 9.3005
R37345 VCC.n9387 VCC.n9386 9.3005
R37346 VCC.n9386 VCC.n9385 9.3005
R37347 VCC.n9385 VCC.n9384 9.3005
R37348 VCC.n9340 VCC.n8927 9.3005
R37349 VCC.n8927 VCC.n8926 9.3005
R37350 VCC.n9298 VCC.n9297 9.3005
R37351 VCC.n9306 VCC.n9305 9.3005
R37352 VCC.n9272 VCC.n9271 9.3005
R37353 VCC.n9261 VCC.n8967 9.3005
R37354 VCC.n8970 VCC.n8969 9.3005
R37355 VCC.n9214 VCC.n9213 9.3005
R37356 VCC.n9213 VCC.n8981 9.3005
R37357 VCC.n8981 VCC.n8980 9.3005
R37358 VCC.n8983 VCC.n8982 9.3005
R37359 VCC.n9229 VCC.n9228 9.3005
R37360 VCC.n9236 VCC.n8976 9.3005
R37361 VCC.n9236 VCC.n9235 9.3005
R37362 VCC.n9235 VCC.n9234 9.3005
R37363 VCC.n9237 VCC.n8977 9.3005
R37364 VCC.n9260 VCC.n9259 9.3005
R37365 VCC.n9264 VCC.n8962 9.3005
R37366 VCC.n9265 VCC.n9264 9.3005
R37367 VCC.n9266 VCC.n9265 9.3005
R37368 VCC.n8957 VCC.n8956 9.3005
R37369 VCC.n9285 VCC.n8945 9.3005
R37370 VCC.n9285 VCC.n8955 9.3005
R37371 VCC.n8955 VCC.n8954 9.3005
R37372 VCC.n8950 VCC.n8948 9.3005
R37373 VCC.n9303 VCC.n8940 9.3005
R37374 VCC.n9303 VCC.n9302 9.3005
R37375 VCC.n9302 VCC.n9301 9.3005
R37376 VCC.n9205 VCC.n9204 9.3005
R37377 VCC.n9206 VCC.n9205 9.3005
R37378 VCC.n9207 VCC.n9206 9.3005
R37379 VCC.n9197 VCC.n9193 9.3005
R37380 VCC.n9199 VCC.n9198 9.3005
R37381 VCC.n9171 VCC.n9170 9.3005
R37382 VCC.n9146 VCC.n9145 9.3005
R37383 VCC.n9034 VCC.n9033 9.3005
R37384 VCC.n9123 VCC.n9122 9.3005
R37385 VCC.n9096 VCC.n9095 9.3005
R37386 VCC.n9096 VCC.n9052 9.3005
R37387 VCC.n9100 VCC.n9052 9.3005
R37388 VCC.n9050 VCC.n9049 9.3005
R37389 VCC.n9106 VCC.n9105 9.3005
R37390 VCC.n9043 VCC.n9042 9.3005
R37391 VCC.n9042 VCC.n9027 9.3005
R37392 VCC.n9027 VCC.n9026 9.3005
R37393 VCC.n9121 VCC.n9041 9.3005
R37394 VCC.n9035 VCC.n9029 9.3005
R37395 VCC.n9024 VCC.n9023 9.3005
R37396 VCC.n9025 VCC.n9024 9.3005
R37397 VCC.n9140 VCC.n9025 9.3005
R37398 VCC.n9018 VCC.n9017 9.3005
R37399 VCC.n9160 VCC.n9007 9.3005
R37400 VCC.n9161 VCC.n9160 9.3005
R37401 VCC.n9162 VCC.n9161 9.3005
R37402 VCC.n9012 VCC.n9010 9.3005
R37403 VCC.n9168 VCC.n9167 9.3005
R37404 VCC.n9087 VCC.n9086 9.3005
R37405 VCC.n9086 VCC.n9085 9.3005
R37406 VCC.n9085 VCC.n9084 9.3005
R37407 VCC.n9069 VCC.n9068 9.3005
R37408 VCC.n9075 VCC.n9074 9.3005
R37409 VCC.n9657 VCC.n9656 9.3005
R37410 VCC.n9626 VCC.n9625 9.3005
R37411 VCC.n9722 VCC.n9721 9.3005
R37412 VCC.n9697 VCC.n9696 9.3005
R37413 VCC.n9585 VCC.n9584 9.3005
R37414 VCC.n9586 VCC.n9580 9.3005
R37415 VCC.n9575 VCC.n9574 9.3005
R37416 VCC.n9576 VCC.n9575 9.3005
R37417 VCC.n9691 VCC.n9576 9.3005
R37418 VCC.n9569 VCC.n9568 9.3005
R37419 VCC.n9711 VCC.n9558 9.3005
R37420 VCC.n9712 VCC.n9711 9.3005
R37421 VCC.n9713 VCC.n9712 9.3005
R37422 VCC.n9563 VCC.n9561 9.3005
R37423 VCC.n9719 VCC.n9718 9.3005
R37424 VCC.n9601 VCC.n9600 9.3005
R37425 VCC.n9638 VCC.n9637 9.3005
R37426 VCC.n9637 VCC.n9636 9.3005
R37427 VCC.n9636 VCC.n9635 9.3005
R37428 VCC.n9620 VCC.n9619 9.3005
R37429 VCC.n9647 VCC.n9646 9.3005
R37430 VCC.n9647 VCC.n9603 9.3005
R37431 VCC.n9651 VCC.n9603 9.3005
R37432 VCC.n9594 VCC.n9593 9.3005
R37433 VCC.n9593 VCC.n9578 9.3005
R37434 VCC.n9578 VCC.n9577 9.3005
R37435 VCC.n9672 VCC.n9592 9.3005
R37436 VCC.n9674 VCC.n9673 9.3005
R37437 VCC.n9781 VCC.n9780 9.3005
R37438 VCC.n9751 VCC.n9750 9.3005
R37439 VCC.n9857 VCC.n9856 9.3005
R37440 VCC.n9824 VCC.n9823 9.3005
R37441 VCC.n9813 VCC.n9519 9.3005
R37442 VCC.n9812 VCC.n9811 9.3005
R37443 VCC.n9509 VCC.n9508 9.3005
R37444 VCC.n9502 VCC.n9500 9.3005
R37445 VCC.n9535 VCC.n9534 9.3005
R37446 VCC.n9749 VCC.n9744 9.3005
R37447 VCC.n9789 VCC.n9529 9.3005
R37448 VCC.n9522 VCC.n9521 9.3005
R37449 VCC.n9816 VCC.n9514 9.3005
R37450 VCC.n9817 VCC.n9816 9.3005
R37451 VCC.n9818 VCC.n9817 9.3005
R37452 VCC.n9837 VCC.n9497 9.3005
R37453 VCC.n9837 VCC.n9507 9.3005
R37454 VCC.n9507 VCC.n9506 9.3005
R37455 VCC.n9854 VCC.n9492 9.3005
R37456 VCC.n9854 VCC.n9853 9.3005
R37457 VCC.n9853 VCC.n9852 9.3005
R37458 VCC.n9757 VCC.n9756 9.3005
R37459 VCC.n9758 VCC.n9757 9.3005
R37460 VCC.n9759 VCC.n9758 9.3005
R37461 VCC.n9766 VCC.n9765 9.3005
R37462 VCC.n9765 VCC.n9533 9.3005
R37463 VCC.n9533 VCC.n9532 9.3005
R37464 VCC.n9788 VCC.n9528 9.3005
R37465 VCC.n9788 VCC.n9787 9.3005
R37466 VCC.n9787 VCC.n9786 9.3005
R37467 VCC.n9947 VCC.n9946 9.3005
R37468 VCC.n9948 VCC.n9947 9.3005
R37469 VCC.n9949 VCC.n9948 9.3005
R37470 VCC.n9893 VCC.n9892 9.3005
R37471 VCC.n9894 VCC.n9893 9.3005
R37472 VCC.n9901 VCC.n9900 9.3005
R37473 VCC.n9914 VCC.n9913 9.3005
R37474 VCC.n9914 VCC.n9466 9.3005
R37475 VCC.n9896 VCC.n9466 9.3005
R37476 VCC.n9940 VCC.n9939 9.3005
R37477 VCC.n9956 VCC.n9955 9.3005
R37478 VCC.n9955 VCC.n9432 9.3005
R37479 VCC.n9432 VCC.n9431 9.3005
R37480 VCC.n9434 VCC.n9433 9.3005
R37481 VCC.n9970 VCC.n9969 9.3005
R37482 VCC.n9849 VCC.n9848 9.3005
R37483 VCC.n10011 VCC.n10010 9.3005
R37484 VCC.n9996 VCC.n9995 9.3005
R37485 VCC.n9994 VCC.n9993 9.3005
R37486 VCC.n10466 VCC.n10465 9.3005
R37487 VCC.n10459 VCC.n10458 9.3005
R37488 VCC.n10458 VCC.n10457 9.3005
R37489 VCC.n10457 VCC.n10456 9.3005
R37490 VCC.n10519 VCC.n10518 9.3005
R37491 VCC.n10519 VCC.n9984 9.3005
R37492 VCC.n10523 VCC.n9984 9.3005
R37493 VCC.n10495 VCC.n10494 9.3005
R37494 VCC.n10494 VCC.n10493 9.3005
R37495 VCC.n10493 VCC.n10492 9.3005
R37496 VCC.n10448 VCC.n10035 9.3005
R37497 VCC.n10035 VCC.n10034 9.3005
R37498 VCC.n10406 VCC.n10405 9.3005
R37499 VCC.n10414 VCC.n10413 9.3005
R37500 VCC.n10380 VCC.n10379 9.3005
R37501 VCC.n10369 VCC.n10075 9.3005
R37502 VCC.n10078 VCC.n10077 9.3005
R37503 VCC.n10322 VCC.n10321 9.3005
R37504 VCC.n10321 VCC.n10089 9.3005
R37505 VCC.n10089 VCC.n10088 9.3005
R37506 VCC.n10091 VCC.n10090 9.3005
R37507 VCC.n10337 VCC.n10336 9.3005
R37508 VCC.n10344 VCC.n10084 9.3005
R37509 VCC.n10344 VCC.n10343 9.3005
R37510 VCC.n10343 VCC.n10342 9.3005
R37511 VCC.n10345 VCC.n10085 9.3005
R37512 VCC.n10368 VCC.n10367 9.3005
R37513 VCC.n10372 VCC.n10070 9.3005
R37514 VCC.n10373 VCC.n10372 9.3005
R37515 VCC.n10374 VCC.n10373 9.3005
R37516 VCC.n10065 VCC.n10064 9.3005
R37517 VCC.n10393 VCC.n10053 9.3005
R37518 VCC.n10393 VCC.n10063 9.3005
R37519 VCC.n10063 VCC.n10062 9.3005
R37520 VCC.n10058 VCC.n10056 9.3005
R37521 VCC.n10411 VCC.n10048 9.3005
R37522 VCC.n10411 VCC.n10410 9.3005
R37523 VCC.n10410 VCC.n10409 9.3005
R37524 VCC.n10313 VCC.n10312 9.3005
R37525 VCC.n10314 VCC.n10313 9.3005
R37526 VCC.n10315 VCC.n10314 9.3005
R37527 VCC.n10305 VCC.n10301 9.3005
R37528 VCC.n10307 VCC.n10306 9.3005
R37529 VCC.n10279 VCC.n10278 9.3005
R37530 VCC.n10254 VCC.n10253 9.3005
R37531 VCC.n10142 VCC.n10141 9.3005
R37532 VCC.n10231 VCC.n10230 9.3005
R37533 VCC.n10204 VCC.n10203 9.3005
R37534 VCC.n10204 VCC.n10160 9.3005
R37535 VCC.n10208 VCC.n10160 9.3005
R37536 VCC.n10158 VCC.n10157 9.3005
R37537 VCC.n10214 VCC.n10213 9.3005
R37538 VCC.n10151 VCC.n10150 9.3005
R37539 VCC.n10150 VCC.n10135 9.3005
R37540 VCC.n10135 VCC.n10134 9.3005
R37541 VCC.n10229 VCC.n10149 9.3005
R37542 VCC.n10143 VCC.n10137 9.3005
R37543 VCC.n10132 VCC.n10131 9.3005
R37544 VCC.n10133 VCC.n10132 9.3005
R37545 VCC.n10248 VCC.n10133 9.3005
R37546 VCC.n10126 VCC.n10125 9.3005
R37547 VCC.n10268 VCC.n10115 9.3005
R37548 VCC.n10269 VCC.n10268 9.3005
R37549 VCC.n10270 VCC.n10269 9.3005
R37550 VCC.n10120 VCC.n10118 9.3005
R37551 VCC.n10276 VCC.n10275 9.3005
R37552 VCC.n10195 VCC.n10194 9.3005
R37553 VCC.n10194 VCC.n10193 9.3005
R37554 VCC.n10193 VCC.n10192 9.3005
R37555 VCC.n10177 VCC.n10176 9.3005
R37556 VCC.n10183 VCC.n10182 9.3005
R37557 VCC.n10764 VCC.n10763 9.3005
R37558 VCC.n10733 VCC.n10732 9.3005
R37559 VCC.n10829 VCC.n10828 9.3005
R37560 VCC.n10804 VCC.n10803 9.3005
R37561 VCC.n10692 VCC.n10691 9.3005
R37562 VCC.n10693 VCC.n10687 9.3005
R37563 VCC.n10682 VCC.n10681 9.3005
R37564 VCC.n10683 VCC.n10682 9.3005
R37565 VCC.n10798 VCC.n10683 9.3005
R37566 VCC.n10676 VCC.n10675 9.3005
R37567 VCC.n10818 VCC.n10665 9.3005
R37568 VCC.n10819 VCC.n10818 9.3005
R37569 VCC.n10820 VCC.n10819 9.3005
R37570 VCC.n10670 VCC.n10668 9.3005
R37571 VCC.n10826 VCC.n10825 9.3005
R37572 VCC.n10708 VCC.n10707 9.3005
R37573 VCC.n10745 VCC.n10744 9.3005
R37574 VCC.n10744 VCC.n10743 9.3005
R37575 VCC.n10743 VCC.n10742 9.3005
R37576 VCC.n10727 VCC.n10726 9.3005
R37577 VCC.n10754 VCC.n10753 9.3005
R37578 VCC.n10754 VCC.n10710 9.3005
R37579 VCC.n10758 VCC.n10710 9.3005
R37580 VCC.n10701 VCC.n10700 9.3005
R37581 VCC.n10700 VCC.n10685 9.3005
R37582 VCC.n10685 VCC.n10684 9.3005
R37583 VCC.n10779 VCC.n10699 9.3005
R37584 VCC.n10781 VCC.n10780 9.3005
R37585 VCC.n10888 VCC.n10887 9.3005
R37586 VCC.n10858 VCC.n10857 9.3005
R37587 VCC.n10964 VCC.n10963 9.3005
R37588 VCC.n10931 VCC.n10930 9.3005
R37589 VCC.n10920 VCC.n10626 9.3005
R37590 VCC.n10919 VCC.n10918 9.3005
R37591 VCC.n10616 VCC.n10615 9.3005
R37592 VCC.n10609 VCC.n10607 9.3005
R37593 VCC.n10642 VCC.n10641 9.3005
R37594 VCC.n10856 VCC.n10851 9.3005
R37595 VCC.n10896 VCC.n10636 9.3005
R37596 VCC.n10629 VCC.n10628 9.3005
R37597 VCC.n10923 VCC.n10621 9.3005
R37598 VCC.n10924 VCC.n10923 9.3005
R37599 VCC.n10925 VCC.n10924 9.3005
R37600 VCC.n10944 VCC.n10604 9.3005
R37601 VCC.n10944 VCC.n10614 9.3005
R37602 VCC.n10614 VCC.n10613 9.3005
R37603 VCC.n10961 VCC.n10599 9.3005
R37604 VCC.n10961 VCC.n10960 9.3005
R37605 VCC.n10960 VCC.n10959 9.3005
R37606 VCC.n10864 VCC.n10863 9.3005
R37607 VCC.n10865 VCC.n10864 9.3005
R37608 VCC.n10866 VCC.n10865 9.3005
R37609 VCC.n10873 VCC.n10872 9.3005
R37610 VCC.n10872 VCC.n10640 9.3005
R37611 VCC.n10640 VCC.n10639 9.3005
R37612 VCC.n10895 VCC.n10635 9.3005
R37613 VCC.n10895 VCC.n10894 9.3005
R37614 VCC.n10894 VCC.n10893 9.3005
R37615 VCC.n11054 VCC.n11053 9.3005
R37616 VCC.n11055 VCC.n11054 9.3005
R37617 VCC.n11056 VCC.n11055 9.3005
R37618 VCC.n11000 VCC.n10999 9.3005
R37619 VCC.n11001 VCC.n11000 9.3005
R37620 VCC.n11008 VCC.n11007 9.3005
R37621 VCC.n11021 VCC.n11020 9.3005
R37622 VCC.n11021 VCC.n10573 9.3005
R37623 VCC.n11003 VCC.n10573 9.3005
R37624 VCC.n11047 VCC.n11046 9.3005
R37625 VCC.n11063 VCC.n11062 9.3005
R37626 VCC.n11062 VCC.n10539 9.3005
R37627 VCC.n10539 VCC.n10538 9.3005
R37628 VCC.n10541 VCC.n10540 9.3005
R37629 VCC.n11077 VCC.n11076 9.3005
R37630 VCC.n10956 VCC.n10955 9.3005
R37631 VCC.n11118 VCC.n11117 9.3005
R37632 VCC.n11103 VCC.n11102 9.3005
R37633 VCC.n11101 VCC.n11100 9.3005
R37634 VCC.n11573 VCC.n11572 9.3005
R37635 VCC.n11566 VCC.n11565 9.3005
R37636 VCC.n11565 VCC.n11564 9.3005
R37637 VCC.n11564 VCC.n11563 9.3005
R37638 VCC.n11626 VCC.n11625 9.3005
R37639 VCC.n11626 VCC.n11091 9.3005
R37640 VCC.n11630 VCC.n11091 9.3005
R37641 VCC.n11602 VCC.n11601 9.3005
R37642 VCC.n11601 VCC.n11600 9.3005
R37643 VCC.n11600 VCC.n11599 9.3005
R37644 VCC.n11555 VCC.n11142 9.3005
R37645 VCC.n11142 VCC.n11141 9.3005
R37646 VCC.n11513 VCC.n11512 9.3005
R37647 VCC.n11521 VCC.n11520 9.3005
R37648 VCC.n11487 VCC.n11486 9.3005
R37649 VCC.n11476 VCC.n11182 9.3005
R37650 VCC.n11185 VCC.n11184 9.3005
R37651 VCC.n11429 VCC.n11428 9.3005
R37652 VCC.n11428 VCC.n11196 9.3005
R37653 VCC.n11196 VCC.n11195 9.3005
R37654 VCC.n11198 VCC.n11197 9.3005
R37655 VCC.n11444 VCC.n11443 9.3005
R37656 VCC.n11451 VCC.n11191 9.3005
R37657 VCC.n11451 VCC.n11450 9.3005
R37658 VCC.n11450 VCC.n11449 9.3005
R37659 VCC.n11452 VCC.n11192 9.3005
R37660 VCC.n11475 VCC.n11474 9.3005
R37661 VCC.n11479 VCC.n11177 9.3005
R37662 VCC.n11480 VCC.n11479 9.3005
R37663 VCC.n11481 VCC.n11480 9.3005
R37664 VCC.n11172 VCC.n11171 9.3005
R37665 VCC.n11500 VCC.n11160 9.3005
R37666 VCC.n11500 VCC.n11170 9.3005
R37667 VCC.n11170 VCC.n11169 9.3005
R37668 VCC.n11165 VCC.n11163 9.3005
R37669 VCC.n11518 VCC.n11155 9.3005
R37670 VCC.n11518 VCC.n11517 9.3005
R37671 VCC.n11517 VCC.n11516 9.3005
R37672 VCC.n11420 VCC.n11419 9.3005
R37673 VCC.n11421 VCC.n11420 9.3005
R37674 VCC.n11422 VCC.n11421 9.3005
R37675 VCC.n11412 VCC.n11408 9.3005
R37676 VCC.n11414 VCC.n11413 9.3005
R37677 VCC.n11386 VCC.n11385 9.3005
R37678 VCC.n11361 VCC.n11360 9.3005
R37679 VCC.n11249 VCC.n11248 9.3005
R37680 VCC.n11338 VCC.n11337 9.3005
R37681 VCC.n11311 VCC.n11310 9.3005
R37682 VCC.n11311 VCC.n11267 9.3005
R37683 VCC.n11315 VCC.n11267 9.3005
R37684 VCC.n11265 VCC.n11264 9.3005
R37685 VCC.n11321 VCC.n11320 9.3005
R37686 VCC.n11258 VCC.n11257 9.3005
R37687 VCC.n11257 VCC.n11242 9.3005
R37688 VCC.n11242 VCC.n11241 9.3005
R37689 VCC.n11336 VCC.n11256 9.3005
R37690 VCC.n11250 VCC.n11244 9.3005
R37691 VCC.n11239 VCC.n11238 9.3005
R37692 VCC.n11240 VCC.n11239 9.3005
R37693 VCC.n11355 VCC.n11240 9.3005
R37694 VCC.n11233 VCC.n11232 9.3005
R37695 VCC.n11375 VCC.n11222 9.3005
R37696 VCC.n11376 VCC.n11375 9.3005
R37697 VCC.n11377 VCC.n11376 9.3005
R37698 VCC.n11227 VCC.n11225 9.3005
R37699 VCC.n11383 VCC.n11382 9.3005
R37700 VCC.n11302 VCC.n11301 9.3005
R37701 VCC.n11301 VCC.n11300 9.3005
R37702 VCC.n11300 VCC.n11299 9.3005
R37703 VCC.n11284 VCC.n11283 9.3005
R37704 VCC.n11290 VCC.n11289 9.3005
R37705 VCC.n11871 VCC.n11870 9.3005
R37706 VCC.n11840 VCC.n11839 9.3005
R37707 VCC.n11936 VCC.n11935 9.3005
R37708 VCC.n11911 VCC.n11910 9.3005
R37709 VCC.n11799 VCC.n11798 9.3005
R37710 VCC.n11800 VCC.n11794 9.3005
R37711 VCC.n11789 VCC.n11788 9.3005
R37712 VCC.n11790 VCC.n11789 9.3005
R37713 VCC.n11905 VCC.n11790 9.3005
R37714 VCC.n11783 VCC.n11782 9.3005
R37715 VCC.n11925 VCC.n11772 9.3005
R37716 VCC.n11926 VCC.n11925 9.3005
R37717 VCC.n11927 VCC.n11926 9.3005
R37718 VCC.n11777 VCC.n11775 9.3005
R37719 VCC.n11933 VCC.n11932 9.3005
R37720 VCC.n11815 VCC.n11814 9.3005
R37721 VCC.n11852 VCC.n11851 9.3005
R37722 VCC.n11851 VCC.n11850 9.3005
R37723 VCC.n11850 VCC.n11849 9.3005
R37724 VCC.n11834 VCC.n11833 9.3005
R37725 VCC.n11861 VCC.n11860 9.3005
R37726 VCC.n11861 VCC.n11817 9.3005
R37727 VCC.n11865 VCC.n11817 9.3005
R37728 VCC.n11808 VCC.n11807 9.3005
R37729 VCC.n11807 VCC.n11792 9.3005
R37730 VCC.n11792 VCC.n11791 9.3005
R37731 VCC.n11886 VCC.n11806 9.3005
R37732 VCC.n11888 VCC.n11887 9.3005
R37733 VCC.n11995 VCC.n11994 9.3005
R37734 VCC.n11965 VCC.n11964 9.3005
R37735 VCC.n12071 VCC.n12070 9.3005
R37736 VCC.n12038 VCC.n12037 9.3005
R37737 VCC.n12027 VCC.n11733 9.3005
R37738 VCC.n12026 VCC.n12025 9.3005
R37739 VCC.n11723 VCC.n11722 9.3005
R37740 VCC.n11716 VCC.n11714 9.3005
R37741 VCC.n11749 VCC.n11748 9.3005
R37742 VCC.n11963 VCC.n11958 9.3005
R37743 VCC.n12003 VCC.n11743 9.3005
R37744 VCC.n11736 VCC.n11735 9.3005
R37745 VCC.n12030 VCC.n11728 9.3005
R37746 VCC.n12031 VCC.n12030 9.3005
R37747 VCC.n12032 VCC.n12031 9.3005
R37748 VCC.n12051 VCC.n11711 9.3005
R37749 VCC.n12051 VCC.n11721 9.3005
R37750 VCC.n11721 VCC.n11720 9.3005
R37751 VCC.n12068 VCC.n11706 9.3005
R37752 VCC.n12068 VCC.n12067 9.3005
R37753 VCC.n12067 VCC.n12066 9.3005
R37754 VCC.n11971 VCC.n11970 9.3005
R37755 VCC.n11972 VCC.n11971 9.3005
R37756 VCC.n11973 VCC.n11972 9.3005
R37757 VCC.n11980 VCC.n11979 9.3005
R37758 VCC.n11979 VCC.n11747 9.3005
R37759 VCC.n11747 VCC.n11746 9.3005
R37760 VCC.n12002 VCC.n11742 9.3005
R37761 VCC.n12002 VCC.n12001 9.3005
R37762 VCC.n12001 VCC.n12000 9.3005
R37763 VCC.n12161 VCC.n12160 9.3005
R37764 VCC.n12162 VCC.n12161 9.3005
R37765 VCC.n12163 VCC.n12162 9.3005
R37766 VCC.n12107 VCC.n12106 9.3005
R37767 VCC.n12108 VCC.n12107 9.3005
R37768 VCC.n12115 VCC.n12114 9.3005
R37769 VCC.n12128 VCC.n12127 9.3005
R37770 VCC.n12128 VCC.n11680 9.3005
R37771 VCC.n12110 VCC.n11680 9.3005
R37772 VCC.n12154 VCC.n12153 9.3005
R37773 VCC.n12170 VCC.n12169 9.3005
R37774 VCC.n12169 VCC.n11646 9.3005
R37775 VCC.n11646 VCC.n11645 9.3005
R37776 VCC.n11648 VCC.n11647 9.3005
R37777 VCC.n12184 VCC.n12183 9.3005
R37778 VCC.n12063 VCC.n12062 9.3005
R37779 VCC.n12225 VCC.n12224 9.3005
R37780 VCC.n12210 VCC.n12209 9.3005
R37781 VCC.n12208 VCC.n12207 9.3005
R37782 VCC.n12680 VCC.n12679 9.3005
R37783 VCC.n12673 VCC.n12672 9.3005
R37784 VCC.n12672 VCC.n12671 9.3005
R37785 VCC.n12671 VCC.n12670 9.3005
R37786 VCC.n12733 VCC.n12732 9.3005
R37787 VCC.n12733 VCC.n12198 9.3005
R37788 VCC.n12737 VCC.n12198 9.3005
R37789 VCC.n12709 VCC.n12708 9.3005
R37790 VCC.n12708 VCC.n12707 9.3005
R37791 VCC.n12707 VCC.n12706 9.3005
R37792 VCC.n12662 VCC.n12249 9.3005
R37793 VCC.n12249 VCC.n12248 9.3005
R37794 VCC.n12620 VCC.n12619 9.3005
R37795 VCC.n12628 VCC.n12627 9.3005
R37796 VCC.n12594 VCC.n12593 9.3005
R37797 VCC.n12583 VCC.n12289 9.3005
R37798 VCC.n12292 VCC.n12291 9.3005
R37799 VCC.n12536 VCC.n12535 9.3005
R37800 VCC.n12535 VCC.n12303 9.3005
R37801 VCC.n12303 VCC.n12302 9.3005
R37802 VCC.n12305 VCC.n12304 9.3005
R37803 VCC.n12551 VCC.n12550 9.3005
R37804 VCC.n12558 VCC.n12298 9.3005
R37805 VCC.n12558 VCC.n12557 9.3005
R37806 VCC.n12557 VCC.n12556 9.3005
R37807 VCC.n12559 VCC.n12299 9.3005
R37808 VCC.n12582 VCC.n12581 9.3005
R37809 VCC.n12586 VCC.n12284 9.3005
R37810 VCC.n12587 VCC.n12586 9.3005
R37811 VCC.n12588 VCC.n12587 9.3005
R37812 VCC.n12279 VCC.n12278 9.3005
R37813 VCC.n12607 VCC.n12267 9.3005
R37814 VCC.n12607 VCC.n12277 9.3005
R37815 VCC.n12277 VCC.n12276 9.3005
R37816 VCC.n12272 VCC.n12270 9.3005
R37817 VCC.n12625 VCC.n12262 9.3005
R37818 VCC.n12625 VCC.n12624 9.3005
R37819 VCC.n12624 VCC.n12623 9.3005
R37820 VCC.n12527 VCC.n12526 9.3005
R37821 VCC.n12528 VCC.n12527 9.3005
R37822 VCC.n12529 VCC.n12528 9.3005
R37823 VCC.n12519 VCC.n12515 9.3005
R37824 VCC.n12521 VCC.n12520 9.3005
R37825 VCC.n12493 VCC.n12492 9.3005
R37826 VCC.n12468 VCC.n12467 9.3005
R37827 VCC.n12356 VCC.n12355 9.3005
R37828 VCC.n12445 VCC.n12444 9.3005
R37829 VCC.n12418 VCC.n12417 9.3005
R37830 VCC.n12418 VCC.n12374 9.3005
R37831 VCC.n12422 VCC.n12374 9.3005
R37832 VCC.n12372 VCC.n12371 9.3005
R37833 VCC.n12428 VCC.n12427 9.3005
R37834 VCC.n12365 VCC.n12364 9.3005
R37835 VCC.n12364 VCC.n12349 9.3005
R37836 VCC.n12349 VCC.n12348 9.3005
R37837 VCC.n12443 VCC.n12363 9.3005
R37838 VCC.n12357 VCC.n12351 9.3005
R37839 VCC.n12346 VCC.n12345 9.3005
R37840 VCC.n12347 VCC.n12346 9.3005
R37841 VCC.n12462 VCC.n12347 9.3005
R37842 VCC.n12340 VCC.n12339 9.3005
R37843 VCC.n12482 VCC.n12329 9.3005
R37844 VCC.n12483 VCC.n12482 9.3005
R37845 VCC.n12484 VCC.n12483 9.3005
R37846 VCC.n12334 VCC.n12332 9.3005
R37847 VCC.n12490 VCC.n12489 9.3005
R37848 VCC.n12409 VCC.n12408 9.3005
R37849 VCC.n12408 VCC.n12407 9.3005
R37850 VCC.n12407 VCC.n12406 9.3005
R37851 VCC.n12391 VCC.n12390 9.3005
R37852 VCC.n12397 VCC.n12396 9.3005
R37853 VCC.n12978 VCC.n12977 9.3005
R37854 VCC.n12947 VCC.n12946 9.3005
R37855 VCC.n13043 VCC.n13042 9.3005
R37856 VCC.n13018 VCC.n13017 9.3005
R37857 VCC.n12906 VCC.n12905 9.3005
R37858 VCC.n12907 VCC.n12901 9.3005
R37859 VCC.n12896 VCC.n12895 9.3005
R37860 VCC.n12897 VCC.n12896 9.3005
R37861 VCC.n13012 VCC.n12897 9.3005
R37862 VCC.n12890 VCC.n12889 9.3005
R37863 VCC.n13032 VCC.n12879 9.3005
R37864 VCC.n13033 VCC.n13032 9.3005
R37865 VCC.n13034 VCC.n13033 9.3005
R37866 VCC.n12884 VCC.n12882 9.3005
R37867 VCC.n13040 VCC.n13039 9.3005
R37868 VCC.n12922 VCC.n12921 9.3005
R37869 VCC.n12959 VCC.n12958 9.3005
R37870 VCC.n12958 VCC.n12957 9.3005
R37871 VCC.n12957 VCC.n12956 9.3005
R37872 VCC.n12941 VCC.n12940 9.3005
R37873 VCC.n12968 VCC.n12967 9.3005
R37874 VCC.n12968 VCC.n12924 9.3005
R37875 VCC.n12972 VCC.n12924 9.3005
R37876 VCC.n12915 VCC.n12914 9.3005
R37877 VCC.n12914 VCC.n12899 9.3005
R37878 VCC.n12899 VCC.n12898 9.3005
R37879 VCC.n12993 VCC.n12913 9.3005
R37880 VCC.n12995 VCC.n12994 9.3005
R37881 VCC.n13102 VCC.n13101 9.3005
R37882 VCC.n13072 VCC.n13071 9.3005
R37883 VCC.n13178 VCC.n13177 9.3005
R37884 VCC.n13145 VCC.n13144 9.3005
R37885 VCC.n13134 VCC.n12840 9.3005
R37886 VCC.n13133 VCC.n13132 9.3005
R37887 VCC.n12830 VCC.n12829 9.3005
R37888 VCC.n12823 VCC.n12821 9.3005
R37889 VCC.n12856 VCC.n12855 9.3005
R37890 VCC.n13070 VCC.n13065 9.3005
R37891 VCC.n13110 VCC.n12850 9.3005
R37892 VCC.n12843 VCC.n12842 9.3005
R37893 VCC.n13137 VCC.n12835 9.3005
R37894 VCC.n13138 VCC.n13137 9.3005
R37895 VCC.n13139 VCC.n13138 9.3005
R37896 VCC.n13158 VCC.n12818 9.3005
R37897 VCC.n13158 VCC.n12828 9.3005
R37898 VCC.n12828 VCC.n12827 9.3005
R37899 VCC.n13175 VCC.n12813 9.3005
R37900 VCC.n13175 VCC.n13174 9.3005
R37901 VCC.n13174 VCC.n13173 9.3005
R37902 VCC.n13078 VCC.n13077 9.3005
R37903 VCC.n13079 VCC.n13078 9.3005
R37904 VCC.n13080 VCC.n13079 9.3005
R37905 VCC.n13087 VCC.n13086 9.3005
R37906 VCC.n13086 VCC.n12854 9.3005
R37907 VCC.n12854 VCC.n12853 9.3005
R37908 VCC.n13109 VCC.n12849 9.3005
R37909 VCC.n13109 VCC.n13108 9.3005
R37910 VCC.n13108 VCC.n13107 9.3005
R37911 VCC.n13268 VCC.n13267 9.3005
R37912 VCC.n13269 VCC.n13268 9.3005
R37913 VCC.n13270 VCC.n13269 9.3005
R37914 VCC.n13214 VCC.n13213 9.3005
R37915 VCC.n13215 VCC.n13214 9.3005
R37916 VCC.n13222 VCC.n13221 9.3005
R37917 VCC.n13235 VCC.n13234 9.3005
R37918 VCC.n13235 VCC.n12787 9.3005
R37919 VCC.n13217 VCC.n12787 9.3005
R37920 VCC.n13261 VCC.n13260 9.3005
R37921 VCC.n13277 VCC.n13276 9.3005
R37922 VCC.n13276 VCC.n12753 9.3005
R37923 VCC.n12753 VCC.n12752 9.3005
R37924 VCC.n12755 VCC.n12754 9.3005
R37925 VCC.n13291 VCC.n13290 9.3005
R37926 VCC.n13170 VCC.n13169 9.3005
R37927 VCC.n13332 VCC.n13331 9.3005
R37928 VCC.n13317 VCC.n13316 9.3005
R37929 VCC.n13315 VCC.n13314 9.3005
R37930 VCC.n13787 VCC.n13786 9.3005
R37931 VCC.n13780 VCC.n13779 9.3005
R37932 VCC.n13779 VCC.n13778 9.3005
R37933 VCC.n13778 VCC.n13777 9.3005
R37934 VCC.n13840 VCC.n13839 9.3005
R37935 VCC.n13840 VCC.n13305 9.3005
R37936 VCC.n13844 VCC.n13305 9.3005
R37937 VCC.n13816 VCC.n13815 9.3005
R37938 VCC.n13815 VCC.n13814 9.3005
R37939 VCC.n13814 VCC.n13813 9.3005
R37940 VCC.n13769 VCC.n13356 9.3005
R37941 VCC.n13356 VCC.n13355 9.3005
R37942 VCC.n13727 VCC.n13726 9.3005
R37943 VCC.n13735 VCC.n13734 9.3005
R37944 VCC.n13701 VCC.n13700 9.3005
R37945 VCC.n13690 VCC.n13396 9.3005
R37946 VCC.n13399 VCC.n13398 9.3005
R37947 VCC.n13643 VCC.n13642 9.3005
R37948 VCC.n13642 VCC.n13410 9.3005
R37949 VCC.n13410 VCC.n13409 9.3005
R37950 VCC.n13412 VCC.n13411 9.3005
R37951 VCC.n13658 VCC.n13657 9.3005
R37952 VCC.n13665 VCC.n13405 9.3005
R37953 VCC.n13665 VCC.n13664 9.3005
R37954 VCC.n13664 VCC.n13663 9.3005
R37955 VCC.n13666 VCC.n13406 9.3005
R37956 VCC.n13689 VCC.n13688 9.3005
R37957 VCC.n13693 VCC.n13391 9.3005
R37958 VCC.n13694 VCC.n13693 9.3005
R37959 VCC.n13695 VCC.n13694 9.3005
R37960 VCC.n13386 VCC.n13385 9.3005
R37961 VCC.n13714 VCC.n13374 9.3005
R37962 VCC.n13714 VCC.n13384 9.3005
R37963 VCC.n13384 VCC.n13383 9.3005
R37964 VCC.n13379 VCC.n13377 9.3005
R37965 VCC.n13732 VCC.n13369 9.3005
R37966 VCC.n13732 VCC.n13731 9.3005
R37967 VCC.n13731 VCC.n13730 9.3005
R37968 VCC.n13634 VCC.n13633 9.3005
R37969 VCC.n13635 VCC.n13634 9.3005
R37970 VCC.n13636 VCC.n13635 9.3005
R37971 VCC.n13626 VCC.n13622 9.3005
R37972 VCC.n13628 VCC.n13627 9.3005
R37973 VCC.n13600 VCC.n13599 9.3005
R37974 VCC.n13575 VCC.n13574 9.3005
R37975 VCC.n13463 VCC.n13462 9.3005
R37976 VCC.n13552 VCC.n13551 9.3005
R37977 VCC.n13525 VCC.n13524 9.3005
R37978 VCC.n13525 VCC.n13481 9.3005
R37979 VCC.n13529 VCC.n13481 9.3005
R37980 VCC.n13479 VCC.n13478 9.3005
R37981 VCC.n13535 VCC.n13534 9.3005
R37982 VCC.n13472 VCC.n13471 9.3005
R37983 VCC.n13471 VCC.n13456 9.3005
R37984 VCC.n13456 VCC.n13455 9.3005
R37985 VCC.n13550 VCC.n13470 9.3005
R37986 VCC.n13464 VCC.n13458 9.3005
R37987 VCC.n13453 VCC.n13452 9.3005
R37988 VCC.n13454 VCC.n13453 9.3005
R37989 VCC.n13569 VCC.n13454 9.3005
R37990 VCC.n13447 VCC.n13446 9.3005
R37991 VCC.n13589 VCC.n13436 9.3005
R37992 VCC.n13590 VCC.n13589 9.3005
R37993 VCC.n13591 VCC.n13590 9.3005
R37994 VCC.n13441 VCC.n13439 9.3005
R37995 VCC.n13597 VCC.n13596 9.3005
R37996 VCC.n13516 VCC.n13515 9.3005
R37997 VCC.n13515 VCC.n13514 9.3005
R37998 VCC.n13514 VCC.n13513 9.3005
R37999 VCC.n13498 VCC.n13497 9.3005
R38000 VCC.n13504 VCC.n13503 9.3005
R38001 VCC.n14085 VCC.n14084 9.3005
R38002 VCC.n14054 VCC.n14053 9.3005
R38003 VCC.n14150 VCC.n14149 9.3005
R38004 VCC.n14125 VCC.n14124 9.3005
R38005 VCC.n14013 VCC.n14012 9.3005
R38006 VCC.n14014 VCC.n14008 9.3005
R38007 VCC.n14003 VCC.n14002 9.3005
R38008 VCC.n14004 VCC.n14003 9.3005
R38009 VCC.n14119 VCC.n14004 9.3005
R38010 VCC.n13997 VCC.n13996 9.3005
R38011 VCC.n14139 VCC.n13986 9.3005
R38012 VCC.n14140 VCC.n14139 9.3005
R38013 VCC.n14141 VCC.n14140 9.3005
R38014 VCC.n13991 VCC.n13989 9.3005
R38015 VCC.n14147 VCC.n14146 9.3005
R38016 VCC.n14029 VCC.n14028 9.3005
R38017 VCC.n14066 VCC.n14065 9.3005
R38018 VCC.n14065 VCC.n14064 9.3005
R38019 VCC.n14064 VCC.n14063 9.3005
R38020 VCC.n14048 VCC.n14047 9.3005
R38021 VCC.n14075 VCC.n14074 9.3005
R38022 VCC.n14075 VCC.n14031 9.3005
R38023 VCC.n14079 VCC.n14031 9.3005
R38024 VCC.n14022 VCC.n14021 9.3005
R38025 VCC.n14021 VCC.n14006 9.3005
R38026 VCC.n14006 VCC.n14005 9.3005
R38027 VCC.n14100 VCC.n14020 9.3005
R38028 VCC.n14102 VCC.n14101 9.3005
R38029 VCC.n14209 VCC.n14208 9.3005
R38030 VCC.n14179 VCC.n14178 9.3005
R38031 VCC.n14285 VCC.n14284 9.3005
R38032 VCC.n14252 VCC.n14251 9.3005
R38033 VCC.n14241 VCC.n13947 9.3005
R38034 VCC.n14240 VCC.n14239 9.3005
R38035 VCC.n13937 VCC.n13936 9.3005
R38036 VCC.n13930 VCC.n13928 9.3005
R38037 VCC.n13963 VCC.n13962 9.3005
R38038 VCC.n14177 VCC.n14172 9.3005
R38039 VCC.n14217 VCC.n13957 9.3005
R38040 VCC.n13950 VCC.n13949 9.3005
R38041 VCC.n14244 VCC.n13942 9.3005
R38042 VCC.n14245 VCC.n14244 9.3005
R38043 VCC.n14246 VCC.n14245 9.3005
R38044 VCC.n14265 VCC.n13925 9.3005
R38045 VCC.n14265 VCC.n13935 9.3005
R38046 VCC.n13935 VCC.n13934 9.3005
R38047 VCC.n14282 VCC.n13920 9.3005
R38048 VCC.n14282 VCC.n14281 9.3005
R38049 VCC.n14281 VCC.n14280 9.3005
R38050 VCC.n14185 VCC.n14184 9.3005
R38051 VCC.n14186 VCC.n14185 9.3005
R38052 VCC.n14187 VCC.n14186 9.3005
R38053 VCC.n14194 VCC.n14193 9.3005
R38054 VCC.n14193 VCC.n13961 9.3005
R38055 VCC.n13961 VCC.n13960 9.3005
R38056 VCC.n14216 VCC.n13956 9.3005
R38057 VCC.n14216 VCC.n14215 9.3005
R38058 VCC.n14215 VCC.n14214 9.3005
R38059 VCC.n14375 VCC.n14374 9.3005
R38060 VCC.n14376 VCC.n14375 9.3005
R38061 VCC.n14377 VCC.n14376 9.3005
R38062 VCC.n14321 VCC.n14320 9.3005
R38063 VCC.n14322 VCC.n14321 9.3005
R38064 VCC.n14329 VCC.n14328 9.3005
R38065 VCC.n14342 VCC.n14341 9.3005
R38066 VCC.n14342 VCC.n13894 9.3005
R38067 VCC.n14324 VCC.n13894 9.3005
R38068 VCC.n14368 VCC.n14367 9.3005
R38069 VCC.n14384 VCC.n14383 9.3005
R38070 VCC.n14383 VCC.n13860 9.3005
R38071 VCC.n13860 VCC.n13859 9.3005
R38072 VCC.n13862 VCC.n13861 9.3005
R38073 VCC.n14398 VCC.n14397 9.3005
R38074 VCC.n14277 VCC.n14276 9.3005
R38075 VCC.n14439 VCC.n14438 9.3005
R38076 VCC.n14424 VCC.n14423 9.3005
R38077 VCC.n14422 VCC.n14421 9.3005
R38078 VCC.n14894 VCC.n14893 9.3005
R38079 VCC.n14887 VCC.n14886 9.3005
R38080 VCC.n14886 VCC.n14885 9.3005
R38081 VCC.n14885 VCC.n14884 9.3005
R38082 VCC.n14947 VCC.n14946 9.3005
R38083 VCC.n14947 VCC.n14412 9.3005
R38084 VCC.n14951 VCC.n14412 9.3005
R38085 VCC.n14923 VCC.n14922 9.3005
R38086 VCC.n14922 VCC.n14921 9.3005
R38087 VCC.n14921 VCC.n14920 9.3005
R38088 VCC.n14876 VCC.n14463 9.3005
R38089 VCC.n14463 VCC.n14462 9.3005
R38090 VCC.n14834 VCC.n14833 9.3005
R38091 VCC.n14842 VCC.n14841 9.3005
R38092 VCC.n14808 VCC.n14807 9.3005
R38093 VCC.n14797 VCC.n14503 9.3005
R38094 VCC.n14506 VCC.n14505 9.3005
R38095 VCC.n14750 VCC.n14749 9.3005
R38096 VCC.n14749 VCC.n14517 9.3005
R38097 VCC.n14517 VCC.n14516 9.3005
R38098 VCC.n14519 VCC.n14518 9.3005
R38099 VCC.n14765 VCC.n14764 9.3005
R38100 VCC.n14772 VCC.n14512 9.3005
R38101 VCC.n14772 VCC.n14771 9.3005
R38102 VCC.n14771 VCC.n14770 9.3005
R38103 VCC.n14773 VCC.n14513 9.3005
R38104 VCC.n14796 VCC.n14795 9.3005
R38105 VCC.n14800 VCC.n14498 9.3005
R38106 VCC.n14801 VCC.n14800 9.3005
R38107 VCC.n14802 VCC.n14801 9.3005
R38108 VCC.n14493 VCC.n14492 9.3005
R38109 VCC.n14821 VCC.n14481 9.3005
R38110 VCC.n14821 VCC.n14491 9.3005
R38111 VCC.n14491 VCC.n14490 9.3005
R38112 VCC.n14486 VCC.n14484 9.3005
R38113 VCC.n14839 VCC.n14476 9.3005
R38114 VCC.n14839 VCC.n14838 9.3005
R38115 VCC.n14838 VCC.n14837 9.3005
R38116 VCC.n14741 VCC.n14740 9.3005
R38117 VCC.n14742 VCC.n14741 9.3005
R38118 VCC.n14743 VCC.n14742 9.3005
R38119 VCC.n14733 VCC.n14729 9.3005
R38120 VCC.n14735 VCC.n14734 9.3005
R38121 VCC.n14707 VCC.n14706 9.3005
R38122 VCC.n14682 VCC.n14681 9.3005
R38123 VCC.n14570 VCC.n14569 9.3005
R38124 VCC.n14659 VCC.n14658 9.3005
R38125 VCC.n14632 VCC.n14631 9.3005
R38126 VCC.n14632 VCC.n14588 9.3005
R38127 VCC.n14636 VCC.n14588 9.3005
R38128 VCC.n14586 VCC.n14585 9.3005
R38129 VCC.n14642 VCC.n14641 9.3005
R38130 VCC.n14579 VCC.n14578 9.3005
R38131 VCC.n14578 VCC.n14563 9.3005
R38132 VCC.n14563 VCC.n14562 9.3005
R38133 VCC.n14657 VCC.n14577 9.3005
R38134 VCC.n14571 VCC.n14565 9.3005
R38135 VCC.n14560 VCC.n14559 9.3005
R38136 VCC.n14561 VCC.n14560 9.3005
R38137 VCC.n14676 VCC.n14561 9.3005
R38138 VCC.n14554 VCC.n14553 9.3005
R38139 VCC.n14696 VCC.n14543 9.3005
R38140 VCC.n14697 VCC.n14696 9.3005
R38141 VCC.n14698 VCC.n14697 9.3005
R38142 VCC.n14548 VCC.n14546 9.3005
R38143 VCC.n14704 VCC.n14703 9.3005
R38144 VCC.n14623 VCC.n14622 9.3005
R38145 VCC.n14622 VCC.n14621 9.3005
R38146 VCC.n14621 VCC.n14620 9.3005
R38147 VCC.n14605 VCC.n14604 9.3005
R38148 VCC.n14611 VCC.n14610 9.3005
R38149 VCC.n15192 VCC.n15191 9.3005
R38150 VCC.n15161 VCC.n15160 9.3005
R38151 VCC.n15257 VCC.n15256 9.3005
R38152 VCC.n15232 VCC.n15231 9.3005
R38153 VCC.n15120 VCC.n15119 9.3005
R38154 VCC.n15121 VCC.n15115 9.3005
R38155 VCC.n15110 VCC.n15109 9.3005
R38156 VCC.n15111 VCC.n15110 9.3005
R38157 VCC.n15226 VCC.n15111 9.3005
R38158 VCC.n15104 VCC.n15103 9.3005
R38159 VCC.n15246 VCC.n15093 9.3005
R38160 VCC.n15247 VCC.n15246 9.3005
R38161 VCC.n15248 VCC.n15247 9.3005
R38162 VCC.n15098 VCC.n15096 9.3005
R38163 VCC.n15254 VCC.n15253 9.3005
R38164 VCC.n15136 VCC.n15135 9.3005
R38165 VCC.n15173 VCC.n15172 9.3005
R38166 VCC.n15172 VCC.n15171 9.3005
R38167 VCC.n15171 VCC.n15170 9.3005
R38168 VCC.n15155 VCC.n15154 9.3005
R38169 VCC.n15182 VCC.n15181 9.3005
R38170 VCC.n15182 VCC.n15138 9.3005
R38171 VCC.n15186 VCC.n15138 9.3005
R38172 VCC.n15129 VCC.n15128 9.3005
R38173 VCC.n15128 VCC.n15113 9.3005
R38174 VCC.n15113 VCC.n15112 9.3005
R38175 VCC.n15207 VCC.n15127 9.3005
R38176 VCC.n15209 VCC.n15208 9.3005
R38177 VCC.n15316 VCC.n15315 9.3005
R38178 VCC.n15286 VCC.n15285 9.3005
R38179 VCC.n15392 VCC.n15391 9.3005
R38180 VCC.n15359 VCC.n15358 9.3005
R38181 VCC.n15348 VCC.n15054 9.3005
R38182 VCC.n15347 VCC.n15346 9.3005
R38183 VCC.n15044 VCC.n15043 9.3005
R38184 VCC.n15037 VCC.n15035 9.3005
R38185 VCC.n15070 VCC.n15069 9.3005
R38186 VCC.n15284 VCC.n15279 9.3005
R38187 VCC.n15324 VCC.n15064 9.3005
R38188 VCC.n15057 VCC.n15056 9.3005
R38189 VCC.n15351 VCC.n15049 9.3005
R38190 VCC.n15352 VCC.n15351 9.3005
R38191 VCC.n15353 VCC.n15352 9.3005
R38192 VCC.n15372 VCC.n15032 9.3005
R38193 VCC.n15372 VCC.n15042 9.3005
R38194 VCC.n15042 VCC.n15041 9.3005
R38195 VCC.n15389 VCC.n15027 9.3005
R38196 VCC.n15389 VCC.n15388 9.3005
R38197 VCC.n15388 VCC.n15387 9.3005
R38198 VCC.n15292 VCC.n15291 9.3005
R38199 VCC.n15293 VCC.n15292 9.3005
R38200 VCC.n15294 VCC.n15293 9.3005
R38201 VCC.n15301 VCC.n15300 9.3005
R38202 VCC.n15300 VCC.n15068 9.3005
R38203 VCC.n15068 VCC.n15067 9.3005
R38204 VCC.n15323 VCC.n15063 9.3005
R38205 VCC.n15323 VCC.n15322 9.3005
R38206 VCC.n15322 VCC.n15321 9.3005
R38207 VCC.n15482 VCC.n15481 9.3005
R38208 VCC.n15483 VCC.n15482 9.3005
R38209 VCC.n15484 VCC.n15483 9.3005
R38210 VCC.n15428 VCC.n15427 9.3005
R38211 VCC.n15429 VCC.n15428 9.3005
R38212 VCC.n15436 VCC.n15435 9.3005
R38213 VCC.n15449 VCC.n15448 9.3005
R38214 VCC.n15449 VCC.n15001 9.3005
R38215 VCC.n15431 VCC.n15001 9.3005
R38216 VCC.n15475 VCC.n15474 9.3005
R38217 VCC.n15491 VCC.n15490 9.3005
R38218 VCC.n15490 VCC.n14967 9.3005
R38219 VCC.n14967 VCC.n14966 9.3005
R38220 VCC.n14969 VCC.n14968 9.3005
R38221 VCC.n15505 VCC.n15504 9.3005
R38222 VCC.n15384 VCC.n15383 9.3005
R38223 VCC.n15546 VCC.n15545 9.3005
R38224 VCC.n15531 VCC.n15530 9.3005
R38225 VCC.n15529 VCC.n15528 9.3005
R38226 VCC.n16001 VCC.n16000 9.3005
R38227 VCC.n15994 VCC.n15993 9.3005
R38228 VCC.n15993 VCC.n15992 9.3005
R38229 VCC.n15992 VCC.n15991 9.3005
R38230 VCC.n16054 VCC.n16053 9.3005
R38231 VCC.n16054 VCC.n15519 9.3005
R38232 VCC.n16058 VCC.n15519 9.3005
R38233 VCC.n16030 VCC.n16029 9.3005
R38234 VCC.n16029 VCC.n16028 9.3005
R38235 VCC.n16028 VCC.n16027 9.3005
R38236 VCC.n15983 VCC.n15570 9.3005
R38237 VCC.n15570 VCC.n15569 9.3005
R38238 VCC.n15941 VCC.n15940 9.3005
R38239 VCC.n15949 VCC.n15948 9.3005
R38240 VCC.n15915 VCC.n15914 9.3005
R38241 VCC.n15904 VCC.n15610 9.3005
R38242 VCC.n15613 VCC.n15612 9.3005
R38243 VCC.n15857 VCC.n15856 9.3005
R38244 VCC.n15856 VCC.n15624 9.3005
R38245 VCC.n15624 VCC.n15623 9.3005
R38246 VCC.n15626 VCC.n15625 9.3005
R38247 VCC.n15872 VCC.n15871 9.3005
R38248 VCC.n15879 VCC.n15619 9.3005
R38249 VCC.n15879 VCC.n15878 9.3005
R38250 VCC.n15878 VCC.n15877 9.3005
R38251 VCC.n15880 VCC.n15620 9.3005
R38252 VCC.n15903 VCC.n15902 9.3005
R38253 VCC.n15907 VCC.n15605 9.3005
R38254 VCC.n15908 VCC.n15907 9.3005
R38255 VCC.n15909 VCC.n15908 9.3005
R38256 VCC.n15600 VCC.n15599 9.3005
R38257 VCC.n15928 VCC.n15588 9.3005
R38258 VCC.n15928 VCC.n15598 9.3005
R38259 VCC.n15598 VCC.n15597 9.3005
R38260 VCC.n15593 VCC.n15591 9.3005
R38261 VCC.n15946 VCC.n15583 9.3005
R38262 VCC.n15946 VCC.n15945 9.3005
R38263 VCC.n15945 VCC.n15944 9.3005
R38264 VCC.n15848 VCC.n15847 9.3005
R38265 VCC.n15849 VCC.n15848 9.3005
R38266 VCC.n15850 VCC.n15849 9.3005
R38267 VCC.n15840 VCC.n15836 9.3005
R38268 VCC.n15842 VCC.n15841 9.3005
R38269 VCC.n15814 VCC.n15813 9.3005
R38270 VCC.n15789 VCC.n15788 9.3005
R38271 VCC.n15677 VCC.n15676 9.3005
R38272 VCC.n15766 VCC.n15765 9.3005
R38273 VCC.n15739 VCC.n15738 9.3005
R38274 VCC.n15739 VCC.n15695 9.3005
R38275 VCC.n15743 VCC.n15695 9.3005
R38276 VCC.n15693 VCC.n15692 9.3005
R38277 VCC.n15749 VCC.n15748 9.3005
R38278 VCC.n15686 VCC.n15685 9.3005
R38279 VCC.n15685 VCC.n15670 9.3005
R38280 VCC.n15670 VCC.n15669 9.3005
R38281 VCC.n15764 VCC.n15684 9.3005
R38282 VCC.n15678 VCC.n15672 9.3005
R38283 VCC.n15667 VCC.n15666 9.3005
R38284 VCC.n15668 VCC.n15667 9.3005
R38285 VCC.n15783 VCC.n15668 9.3005
R38286 VCC.n15661 VCC.n15660 9.3005
R38287 VCC.n15803 VCC.n15650 9.3005
R38288 VCC.n15804 VCC.n15803 9.3005
R38289 VCC.n15805 VCC.n15804 9.3005
R38290 VCC.n15655 VCC.n15653 9.3005
R38291 VCC.n15811 VCC.n15810 9.3005
R38292 VCC.n15730 VCC.n15729 9.3005
R38293 VCC.n15729 VCC.n15728 9.3005
R38294 VCC.n15728 VCC.n15727 9.3005
R38295 VCC.n15712 VCC.n15711 9.3005
R38296 VCC.n15718 VCC.n15717 9.3005
R38297 VCC.n16299 VCC.n16298 9.3005
R38298 VCC.n16268 VCC.n16267 9.3005
R38299 VCC.n16364 VCC.n16363 9.3005
R38300 VCC.n16339 VCC.n16338 9.3005
R38301 VCC.n16227 VCC.n16226 9.3005
R38302 VCC.n16228 VCC.n16222 9.3005
R38303 VCC.n16217 VCC.n16216 9.3005
R38304 VCC.n16218 VCC.n16217 9.3005
R38305 VCC.n16333 VCC.n16218 9.3005
R38306 VCC.n16211 VCC.n16210 9.3005
R38307 VCC.n16353 VCC.n16200 9.3005
R38308 VCC.n16354 VCC.n16353 9.3005
R38309 VCC.n16355 VCC.n16354 9.3005
R38310 VCC.n16205 VCC.n16203 9.3005
R38311 VCC.n16361 VCC.n16360 9.3005
R38312 VCC.n16243 VCC.n16242 9.3005
R38313 VCC.n16280 VCC.n16279 9.3005
R38314 VCC.n16279 VCC.n16278 9.3005
R38315 VCC.n16278 VCC.n16277 9.3005
R38316 VCC.n16262 VCC.n16261 9.3005
R38317 VCC.n16289 VCC.n16288 9.3005
R38318 VCC.n16289 VCC.n16245 9.3005
R38319 VCC.n16293 VCC.n16245 9.3005
R38320 VCC.n16236 VCC.n16235 9.3005
R38321 VCC.n16235 VCC.n16220 9.3005
R38322 VCC.n16220 VCC.n16219 9.3005
R38323 VCC.n16314 VCC.n16234 9.3005
R38324 VCC.n16316 VCC.n16315 9.3005
R38325 VCC.n16423 VCC.n16422 9.3005
R38326 VCC.n16393 VCC.n16392 9.3005
R38327 VCC.n16499 VCC.n16498 9.3005
R38328 VCC.n16466 VCC.n16465 9.3005
R38329 VCC.n16455 VCC.n16161 9.3005
R38330 VCC.n16454 VCC.n16453 9.3005
R38331 VCC.n16151 VCC.n16150 9.3005
R38332 VCC.n16144 VCC.n16142 9.3005
R38333 VCC.n16177 VCC.n16176 9.3005
R38334 VCC.n16391 VCC.n16386 9.3005
R38335 VCC.n16431 VCC.n16171 9.3005
R38336 VCC.n16164 VCC.n16163 9.3005
R38337 VCC.n16458 VCC.n16156 9.3005
R38338 VCC.n16459 VCC.n16458 9.3005
R38339 VCC.n16460 VCC.n16459 9.3005
R38340 VCC.n16479 VCC.n16139 9.3005
R38341 VCC.n16479 VCC.n16149 9.3005
R38342 VCC.n16149 VCC.n16148 9.3005
R38343 VCC.n16496 VCC.n16134 9.3005
R38344 VCC.n16496 VCC.n16495 9.3005
R38345 VCC.n16495 VCC.n16494 9.3005
R38346 VCC.n16399 VCC.n16398 9.3005
R38347 VCC.n16400 VCC.n16399 9.3005
R38348 VCC.n16401 VCC.n16400 9.3005
R38349 VCC.n16408 VCC.n16407 9.3005
R38350 VCC.n16407 VCC.n16175 9.3005
R38351 VCC.n16175 VCC.n16174 9.3005
R38352 VCC.n16430 VCC.n16170 9.3005
R38353 VCC.n16430 VCC.n16429 9.3005
R38354 VCC.n16429 VCC.n16428 9.3005
R38355 VCC.n16589 VCC.n16588 9.3005
R38356 VCC.n16590 VCC.n16589 9.3005
R38357 VCC.n16591 VCC.n16590 9.3005
R38358 VCC.n16535 VCC.n16534 9.3005
R38359 VCC.n16536 VCC.n16535 9.3005
R38360 VCC.n16543 VCC.n16542 9.3005
R38361 VCC.n16556 VCC.n16555 9.3005
R38362 VCC.n16556 VCC.n16108 9.3005
R38363 VCC.n16538 VCC.n16108 9.3005
R38364 VCC.n16582 VCC.n16581 9.3005
R38365 VCC.n16598 VCC.n16597 9.3005
R38366 VCC.n16597 VCC.n16074 9.3005
R38367 VCC.n16074 VCC.n16073 9.3005
R38368 VCC.n16076 VCC.n16075 9.3005
R38369 VCC.n16612 VCC.n16611 9.3005
R38370 VCC.n16491 VCC.n16490 9.3005
R38371 VCC.n16653 VCC.n16652 9.3005
R38372 VCC.n16638 VCC.n16637 9.3005
R38373 VCC.n16636 VCC.n16635 9.3005
R38374 VCC.n17108 VCC.n17107 9.3005
R38375 VCC.n17101 VCC.n17100 9.3005
R38376 VCC.n17100 VCC.n17099 9.3005
R38377 VCC.n17099 VCC.n17098 9.3005
R38378 VCC.n17161 VCC.n17160 9.3005
R38379 VCC.n17161 VCC.n16626 9.3005
R38380 VCC.n17165 VCC.n16626 9.3005
R38381 VCC.n17137 VCC.n17136 9.3005
R38382 VCC.n17136 VCC.n17135 9.3005
R38383 VCC.n17135 VCC.n17134 9.3005
R38384 VCC.n17090 VCC.n16677 9.3005
R38385 VCC.n16677 VCC.n16676 9.3005
R38386 VCC.n17048 VCC.n17047 9.3005
R38387 VCC.n17056 VCC.n17055 9.3005
R38388 VCC.n17022 VCC.n17021 9.3005
R38389 VCC.n17011 VCC.n16717 9.3005
R38390 VCC.n16720 VCC.n16719 9.3005
R38391 VCC.n16964 VCC.n16963 9.3005
R38392 VCC.n16963 VCC.n16731 9.3005
R38393 VCC.n16731 VCC.n16730 9.3005
R38394 VCC.n16733 VCC.n16732 9.3005
R38395 VCC.n16979 VCC.n16978 9.3005
R38396 VCC.n16986 VCC.n16726 9.3005
R38397 VCC.n16986 VCC.n16985 9.3005
R38398 VCC.n16985 VCC.n16984 9.3005
R38399 VCC.n16987 VCC.n16727 9.3005
R38400 VCC.n17010 VCC.n17009 9.3005
R38401 VCC.n17014 VCC.n16712 9.3005
R38402 VCC.n17015 VCC.n17014 9.3005
R38403 VCC.n17016 VCC.n17015 9.3005
R38404 VCC.n16707 VCC.n16706 9.3005
R38405 VCC.n17035 VCC.n16695 9.3005
R38406 VCC.n17035 VCC.n16705 9.3005
R38407 VCC.n16705 VCC.n16704 9.3005
R38408 VCC.n16700 VCC.n16698 9.3005
R38409 VCC.n17053 VCC.n16690 9.3005
R38410 VCC.n17053 VCC.n17052 9.3005
R38411 VCC.n17052 VCC.n17051 9.3005
R38412 VCC.n16955 VCC.n16954 9.3005
R38413 VCC.n16956 VCC.n16955 9.3005
R38414 VCC.n16957 VCC.n16956 9.3005
R38415 VCC.n16947 VCC.n16943 9.3005
R38416 VCC.n16949 VCC.n16948 9.3005
R38417 VCC.n16921 VCC.n16920 9.3005
R38418 VCC.n16896 VCC.n16895 9.3005
R38419 VCC.n16784 VCC.n16783 9.3005
R38420 VCC.n16873 VCC.n16872 9.3005
R38421 VCC.n16846 VCC.n16845 9.3005
R38422 VCC.n16846 VCC.n16802 9.3005
R38423 VCC.n16850 VCC.n16802 9.3005
R38424 VCC.n16800 VCC.n16799 9.3005
R38425 VCC.n16856 VCC.n16855 9.3005
R38426 VCC.n16793 VCC.n16792 9.3005
R38427 VCC.n16792 VCC.n16777 9.3005
R38428 VCC.n16777 VCC.n16776 9.3005
R38429 VCC.n16871 VCC.n16791 9.3005
R38430 VCC.n16785 VCC.n16779 9.3005
R38431 VCC.n16774 VCC.n16773 9.3005
R38432 VCC.n16775 VCC.n16774 9.3005
R38433 VCC.n16890 VCC.n16775 9.3005
R38434 VCC.n16768 VCC.n16767 9.3005
R38435 VCC.n16910 VCC.n16757 9.3005
R38436 VCC.n16911 VCC.n16910 9.3005
R38437 VCC.n16912 VCC.n16911 9.3005
R38438 VCC.n16762 VCC.n16760 9.3005
R38439 VCC.n16918 VCC.n16917 9.3005
R38440 VCC.n16837 VCC.n16836 9.3005
R38441 VCC.n16836 VCC.n16835 9.3005
R38442 VCC.n16835 VCC.n16834 9.3005
R38443 VCC.n16819 VCC.n16818 9.3005
R38444 VCC.n16825 VCC.n16824 9.3005
R38445 VCC.n17343 VCC.n17342 9.3005
R38446 VCC.n17313 VCC.n17312 9.3005
R38447 VCC.n17419 VCC.n17418 9.3005
R38448 VCC.n17386 VCC.n17385 9.3005
R38449 VCC.n17375 VCC.n17268 9.3005
R38450 VCC.n17374 VCC.n17373 9.3005
R38451 VCC.n17258 VCC.n17257 9.3005
R38452 VCC.n17251 VCC.n17249 9.3005
R38453 VCC.n17284 VCC.n17283 9.3005
R38454 VCC.n17311 VCC.n17306 9.3005
R38455 VCC.n17351 VCC.n17278 9.3005
R38456 VCC.n17271 VCC.n17270 9.3005
R38457 VCC.n17378 VCC.n17263 9.3005
R38458 VCC.n17379 VCC.n17378 9.3005
R38459 VCC.n17380 VCC.n17379 9.3005
R38460 VCC.n17399 VCC.n17246 9.3005
R38461 VCC.n17399 VCC.n17256 9.3005
R38462 VCC.n17256 VCC.n17255 9.3005
R38463 VCC.n17416 VCC.n17241 9.3005
R38464 VCC.n17416 VCC.n17415 9.3005
R38465 VCC.n17415 VCC.n17414 9.3005
R38466 VCC.n17319 VCC.n17318 9.3005
R38467 VCC.n17320 VCC.n17319 9.3005
R38468 VCC.n17321 VCC.n17320 9.3005
R38469 VCC.n17328 VCC.n17327 9.3005
R38470 VCC.n17327 VCC.n17282 9.3005
R38471 VCC.n17282 VCC.n17281 9.3005
R38472 VCC.n17350 VCC.n17277 9.3005
R38473 VCC.n17350 VCC.n17349 9.3005
R38474 VCC.n17349 VCC.n17348 9.3005
R38475 VCC.n17509 VCC.n17508 9.3005
R38476 VCC.n17510 VCC.n17509 9.3005
R38477 VCC.n17511 VCC.n17510 9.3005
R38478 VCC.n17455 VCC.n17454 9.3005
R38479 VCC.n17456 VCC.n17455 9.3005
R38480 VCC.n17463 VCC.n17462 9.3005
R38481 VCC.n17476 VCC.n17475 9.3005
R38482 VCC.n17476 VCC.n17215 9.3005
R38483 VCC.n17458 VCC.n17215 9.3005
R38484 VCC.n17502 VCC.n17501 9.3005
R38485 VCC.n17518 VCC.n17517 9.3005
R38486 VCC.n17517 VCC.n17181 9.3005
R38487 VCC.n17181 VCC.n17180 9.3005
R38488 VCC.n17183 VCC.n17182 9.3005
R38489 VCC.n17532 VCC.n17531 9.3005
R38490 VCC.n17411 VCC.n17410 9.3005
R38491 VCC.n210 VCC.n209 9.13511
R38492 VCC.n122 VCC.n120 9.13511
R38493 VCC.n427 VCC.n426 9.13511
R38494 VCC.n762 VCC.n761 9.13511
R38495 VCC.n674 VCC.n672 9.13511
R38496 VCC.n979 VCC.n978 9.13511
R38497 VCC.n1231 VCC.n1229 9.13511
R38498 VCC.n1537 VCC.n1536 9.13511
R38499 VCC.n1320 VCC.n1319 9.13511
R38500 VCC.n1871 VCC.n1870 9.13511
R38501 VCC.n1783 VCC.n1781 9.13511
R38502 VCC.n2088 VCC.n2087 9.13511
R38503 VCC.n2340 VCC.n2338 9.13511
R38504 VCC.n2646 VCC.n2645 9.13511
R38505 VCC.n2429 VCC.n2428 9.13511
R38506 VCC.n2980 VCC.n2979 9.13511
R38507 VCC.n2892 VCC.n2890 9.13511
R38508 VCC.n3197 VCC.n3196 9.13511
R38509 VCC.n3449 VCC.n3447 9.13511
R38510 VCC.n3755 VCC.n3754 9.13511
R38511 VCC.n3538 VCC.n3537 9.13511
R38512 VCC.n4089 VCC.n4088 9.13511
R38513 VCC.n4001 VCC.n3999 9.13511
R38514 VCC.n4306 VCC.n4305 9.13511
R38515 VCC.n4558 VCC.n4556 9.13511
R38516 VCC.n4864 VCC.n4863 9.13511
R38517 VCC.n4647 VCC.n4646 9.13511
R38518 VCC.n5198 VCC.n5197 9.13511
R38519 VCC.n5110 VCC.n5108 9.13511
R38520 VCC.n5415 VCC.n5414 9.13511
R38521 VCC.n5667 VCC.n5665 9.13511
R38522 VCC.n5973 VCC.n5972 9.13511
R38523 VCC.n5756 VCC.n5755 9.13511
R38524 VCC.n6307 VCC.n6306 9.13511
R38525 VCC.n6219 VCC.n6217 9.13511
R38526 VCC.n6524 VCC.n6523 9.13511
R38527 VCC.n6776 VCC.n6774 9.13511
R38528 VCC.n7082 VCC.n7081 9.13511
R38529 VCC.n6865 VCC.n6864 9.13511
R38530 VCC.n7416 VCC.n7415 9.13511
R38531 VCC.n7328 VCC.n7326 9.13511
R38532 VCC.n7633 VCC.n7632 9.13511
R38533 VCC.n7885 VCC.n7883 9.13511
R38534 VCC.n8191 VCC.n8190 9.13511
R38535 VCC.n7974 VCC.n7973 9.13511
R38536 VCC.n8437 VCC.n8435 9.13511
R38537 VCC.n8742 VCC.n8741 9.13511
R38538 VCC.n8525 VCC.n8524 9.13511
R38539 VCC.n8994 VCC.n8992 9.13511
R38540 VCC.n9300 VCC.n9299 9.13511
R38541 VCC.n9083 VCC.n9082 9.13511
R38542 VCC.n9634 VCC.n9633 9.13511
R38543 VCC.n9546 VCC.n9544 9.13511
R38544 VCC.n9851 VCC.n9850 9.13511
R38545 VCC.n10102 VCC.n10100 9.13511
R38546 VCC.n10408 VCC.n10407 9.13511
R38547 VCC.n10191 VCC.n10190 9.13511
R38548 VCC.n10741 VCC.n10740 9.13511
R38549 VCC.n10653 VCC.n10651 9.13511
R38550 VCC.n10958 VCC.n10957 9.13511
R38551 VCC.n11209 VCC.n11207 9.13511
R38552 VCC.n11515 VCC.n11514 9.13511
R38553 VCC.n11298 VCC.n11297 9.13511
R38554 VCC.n11848 VCC.n11847 9.13511
R38555 VCC.n11760 VCC.n11758 9.13511
R38556 VCC.n12065 VCC.n12064 9.13511
R38557 VCC.n12316 VCC.n12314 9.13511
R38558 VCC.n12622 VCC.n12621 9.13511
R38559 VCC.n12405 VCC.n12404 9.13511
R38560 VCC.n12955 VCC.n12954 9.13511
R38561 VCC.n12867 VCC.n12865 9.13511
R38562 VCC.n13172 VCC.n13171 9.13511
R38563 VCC.n13423 VCC.n13421 9.13511
R38564 VCC.n13729 VCC.n13728 9.13511
R38565 VCC.n13512 VCC.n13511 9.13511
R38566 VCC.n14062 VCC.n14061 9.13511
R38567 VCC.n13974 VCC.n13972 9.13511
R38568 VCC.n14279 VCC.n14278 9.13511
R38569 VCC.n14530 VCC.n14528 9.13511
R38570 VCC.n14836 VCC.n14835 9.13511
R38571 VCC.n14619 VCC.n14618 9.13511
R38572 VCC.n15169 VCC.n15168 9.13511
R38573 VCC.n15081 VCC.n15079 9.13511
R38574 VCC.n15386 VCC.n15385 9.13511
R38575 VCC.n15637 VCC.n15635 9.13511
R38576 VCC.n15943 VCC.n15942 9.13511
R38577 VCC.n15726 VCC.n15725 9.13511
R38578 VCC.n16276 VCC.n16275 9.13511
R38579 VCC.n16188 VCC.n16186 9.13511
R38580 VCC.n16493 VCC.n16492 9.13511
R38581 VCC.n16744 VCC.n16742 9.13511
R38582 VCC.n17050 VCC.n17049 9.13511
R38583 VCC.n16833 VCC.n16832 9.13511
R38584 VCC.n17295 VCC.n17293 9.13511
R38585 VCC.n17413 VCC.n17412 9.13511
R38586 VCC.n423 VCC.n56 8.95764
R38587 VCC.n546 VCC.n4 8.95764
R38588 VCC.n975 VCC.n608 8.95764
R38589 VCC.n1100 VCC.n558 8.95764
R38590 VCC.n1533 VCC.n1530 8.95764
R38591 VCC.n1655 VCC.n1654 8.95764
R38592 VCC.n2084 VCC.n1717 8.95764
R38593 VCC.n2209 VCC.n1667 8.95764
R38594 VCC.n2642 VCC.n2639 8.95764
R38595 VCC.n2764 VCC.n2763 8.95764
R38596 VCC.n3193 VCC.n2826 8.95764
R38597 VCC.n3318 VCC.n2776 8.95764
R38598 VCC.n3751 VCC.n3748 8.95764
R38599 VCC.n3873 VCC.n3872 8.95764
R38600 VCC.n4302 VCC.n3935 8.95764
R38601 VCC.n4427 VCC.n3885 8.95764
R38602 VCC.n4860 VCC.n4857 8.95764
R38603 VCC.n4982 VCC.n4981 8.95764
R38604 VCC.n5411 VCC.n5044 8.95764
R38605 VCC.n5536 VCC.n4994 8.95764
R38606 VCC.n5969 VCC.n5966 8.95764
R38607 VCC.n6091 VCC.n6090 8.95764
R38608 VCC.n6520 VCC.n6153 8.95764
R38609 VCC.n6645 VCC.n6103 8.95764
R38610 VCC.n7078 VCC.n7075 8.95764
R38611 VCC.n7200 VCC.n7199 8.95764
R38612 VCC.n7629 VCC.n7262 8.95764
R38613 VCC.n7754 VCC.n7212 8.95764
R38614 VCC.n8187 VCC.n8184 8.95764
R38615 VCC.n8309 VCC.n8308 8.95764
R38616 VCC.n8738 VCC.n8371 8.95764
R38617 VCC.n8863 VCC.n8321 8.95764
R38618 VCC.n9296 VCC.n9293 8.95764
R38619 VCC.n9418 VCC.n9417 8.95764
R38620 VCC.n9847 VCC.n9480 8.95764
R38621 VCC.n9972 VCC.n9430 8.95764
R38622 VCC.n10404 VCC.n10401 8.95764
R38623 VCC.n10526 VCC.n10525 8.95764
R38624 VCC.n10954 VCC.n10587 8.95764
R38625 VCC.n11079 VCC.n10537 8.95764
R38626 VCC.n11511 VCC.n11508 8.95764
R38627 VCC.n11633 VCC.n11632 8.95764
R38628 VCC.n12061 VCC.n11694 8.95764
R38629 VCC.n12186 VCC.n11644 8.95764
R38630 VCC.n12618 VCC.n12615 8.95764
R38631 VCC.n12740 VCC.n12739 8.95764
R38632 VCC.n13168 VCC.n12801 8.95764
R38633 VCC.n13293 VCC.n12751 8.95764
R38634 VCC.n13725 VCC.n13722 8.95764
R38635 VCC.n13847 VCC.n13846 8.95764
R38636 VCC.n14275 VCC.n13908 8.95764
R38637 VCC.n14400 VCC.n13858 8.95764
R38638 VCC.n14832 VCC.n14829 8.95764
R38639 VCC.n14954 VCC.n14953 8.95764
R38640 VCC.n15382 VCC.n15015 8.95764
R38641 VCC.n15507 VCC.n14965 8.95764
R38642 VCC.n15939 VCC.n15936 8.95764
R38643 VCC.n16061 VCC.n16060 8.95764
R38644 VCC.n16489 VCC.n16122 8.95764
R38645 VCC.n16614 VCC.n16072 8.95764
R38646 VCC.n17046 VCC.n17043 8.95764
R38647 VCC.n17168 VCC.n17167 8.95764
R38648 VCC.n17409 VCC.n17229 8.95764
R38649 VCC.n17534 VCC.n17179 8.95764
R38650 VCC.n499 VCC.n40 8.85536
R38651 VCC.n495 VCC.n40 8.85536
R38652 VCC.n1051 VCC.n592 8.85536
R38653 VCC.n1047 VCC.n592 8.85536
R38654 VCC.n1616 VCC.n1144 8.85536
R38655 VCC.n1144 VCC.n1143 8.85536
R38656 VCC.n2160 VCC.n1701 8.85536
R38657 VCC.n2156 VCC.n1701 8.85536
R38658 VCC.n2725 VCC.n2253 8.85536
R38659 VCC.n2253 VCC.n2252 8.85536
R38660 VCC.n3269 VCC.n2810 8.85536
R38661 VCC.n3265 VCC.n2810 8.85536
R38662 VCC.n3834 VCC.n3362 8.85536
R38663 VCC.n3362 VCC.n3361 8.85536
R38664 VCC.n4378 VCC.n3919 8.85536
R38665 VCC.n4374 VCC.n3919 8.85536
R38666 VCC.n4943 VCC.n4471 8.85536
R38667 VCC.n4471 VCC.n4470 8.85536
R38668 VCC.n5487 VCC.n5028 8.85536
R38669 VCC.n5483 VCC.n5028 8.85536
R38670 VCC.n6052 VCC.n5580 8.85536
R38671 VCC.n5580 VCC.n5579 8.85536
R38672 VCC.n6596 VCC.n6137 8.85536
R38673 VCC.n6592 VCC.n6137 8.85536
R38674 VCC.n7161 VCC.n6689 8.85536
R38675 VCC.n6689 VCC.n6688 8.85536
R38676 VCC.n7705 VCC.n7246 8.85536
R38677 VCC.n7701 VCC.n7246 8.85536
R38678 VCC.n8270 VCC.n7798 8.85536
R38679 VCC.n7798 VCC.n7797 8.85536
R38680 VCC.n8814 VCC.n8355 8.85536
R38681 VCC.n8810 VCC.n8355 8.85536
R38682 VCC.n9379 VCC.n8907 8.85536
R38683 VCC.n8907 VCC.n8906 8.85536
R38684 VCC.n9923 VCC.n9464 8.85536
R38685 VCC.n9919 VCC.n9464 8.85536
R38686 VCC.n10487 VCC.n10015 8.85536
R38687 VCC.n10015 VCC.n10014 8.85536
R38688 VCC.n11030 VCC.n10571 8.85536
R38689 VCC.n11026 VCC.n10571 8.85536
R38690 VCC.n11594 VCC.n11122 8.85536
R38691 VCC.n11122 VCC.n11121 8.85536
R38692 VCC.n12137 VCC.n11678 8.85536
R38693 VCC.n12133 VCC.n11678 8.85536
R38694 VCC.n12701 VCC.n12229 8.85536
R38695 VCC.n12229 VCC.n12228 8.85536
R38696 VCC.n13244 VCC.n12785 8.85536
R38697 VCC.n13240 VCC.n12785 8.85536
R38698 VCC.n13808 VCC.n13336 8.85536
R38699 VCC.n13336 VCC.n13335 8.85536
R38700 VCC.n14351 VCC.n13892 8.85536
R38701 VCC.n14347 VCC.n13892 8.85536
R38702 VCC.n14915 VCC.n14443 8.85536
R38703 VCC.n14443 VCC.n14442 8.85536
R38704 VCC.n15458 VCC.n14999 8.85536
R38705 VCC.n15454 VCC.n14999 8.85536
R38706 VCC.n16022 VCC.n15550 8.85536
R38707 VCC.n15550 VCC.n15549 8.85536
R38708 VCC.n16565 VCC.n16106 8.85536
R38709 VCC.n16561 VCC.n16106 8.85536
R38710 VCC.n17129 VCC.n16657 8.85536
R38711 VCC.n16657 VCC.n16656 8.85536
R38712 VCC.n17485 VCC.n17213 8.85536
R38713 VCC.n17481 VCC.n17213 8.85536
R38714 VCC.n295 VCC.n293 8.47776
R38715 VCC.n847 VCC.n845 8.47776
R38716 VCC.n1405 VCC.n1403 8.47776
R38717 VCC.n1956 VCC.n1954 8.47776
R38718 VCC.n2514 VCC.n2512 8.47776
R38719 VCC.n3065 VCC.n3063 8.47776
R38720 VCC.n3623 VCC.n3621 8.47776
R38721 VCC.n4174 VCC.n4172 8.47776
R38722 VCC.n4732 VCC.n4730 8.47776
R38723 VCC.n5283 VCC.n5281 8.47776
R38724 VCC.n5841 VCC.n5839 8.47776
R38725 VCC.n6392 VCC.n6390 8.47776
R38726 VCC.n6950 VCC.n6948 8.47776
R38727 VCC.n7501 VCC.n7499 8.47776
R38728 VCC.n8059 VCC.n8057 8.47776
R38729 VCC.n8610 VCC.n8608 8.47776
R38730 VCC.n9168 VCC.n9166 8.47776
R38731 VCC.n9719 VCC.n9717 8.47776
R38732 VCC.n10276 VCC.n10274 8.47776
R38733 VCC.n10826 VCC.n10824 8.47776
R38734 VCC.n11383 VCC.n11381 8.47776
R38735 VCC.n11933 VCC.n11931 8.47776
R38736 VCC.n12490 VCC.n12488 8.47776
R38737 VCC.n13040 VCC.n13038 8.47776
R38738 VCC.n13597 VCC.n13595 8.47776
R38739 VCC.n14147 VCC.n14145 8.47776
R38740 VCC.n14704 VCC.n14702 8.47776
R38741 VCC.n15254 VCC.n15252 8.47776
R38742 VCC.n15811 VCC.n15809 8.47776
R38743 VCC.n16361 VCC.n16359 8.47776
R38744 VCC.n16918 VCC.n16916 8.47776
R38745 VCC.n471 VCC.n470 7.03754
R38746 VCC.n527 VCC.n5 7.03754
R38747 VCC.n1023 VCC.n1022 7.03754
R38748 VCC.n1079 VCC.n559 7.03754
R38749 VCC.n1580 VCC.n1163 7.03754
R38750 VCC.n1652 VCC.n1651 7.03754
R38751 VCC.n2132 VCC.n2131 7.03754
R38752 VCC.n2188 VCC.n1668 7.03754
R38753 VCC.n2689 VCC.n2272 7.03754
R38754 VCC.n2761 VCC.n2760 7.03754
R38755 VCC.n3241 VCC.n3240 7.03754
R38756 VCC.n3297 VCC.n2777 7.03754
R38757 VCC.n3798 VCC.n3381 7.03754
R38758 VCC.n3870 VCC.n3869 7.03754
R38759 VCC.n4350 VCC.n4349 7.03754
R38760 VCC.n4406 VCC.n3886 7.03754
R38761 VCC.n4907 VCC.n4490 7.03754
R38762 VCC.n4979 VCC.n4978 7.03754
R38763 VCC.n5459 VCC.n5458 7.03754
R38764 VCC.n5515 VCC.n4995 7.03754
R38765 VCC.n6016 VCC.n5599 7.03754
R38766 VCC.n6088 VCC.n6087 7.03754
R38767 VCC.n6568 VCC.n6567 7.03754
R38768 VCC.n6624 VCC.n6104 7.03754
R38769 VCC.n7125 VCC.n6708 7.03754
R38770 VCC.n7197 VCC.n7196 7.03754
R38771 VCC.n7677 VCC.n7676 7.03754
R38772 VCC.n7733 VCC.n7213 7.03754
R38773 VCC.n8234 VCC.n7817 7.03754
R38774 VCC.n8306 VCC.n8305 7.03754
R38775 VCC.n8786 VCC.n8785 7.03754
R38776 VCC.n8842 VCC.n8322 7.03754
R38777 VCC.n9343 VCC.n8926 7.03754
R38778 VCC.n9415 VCC.n9414 7.03754
R38779 VCC.n9895 VCC.n9894 7.03754
R38780 VCC.n9951 VCC.n9431 7.03754
R38781 VCC.n10451 VCC.n10034 7.03754
R38782 VCC.n10523 VCC.n10522 7.03754
R38783 VCC.n11002 VCC.n11001 7.03754
R38784 VCC.n11058 VCC.n10538 7.03754
R38785 VCC.n11558 VCC.n11141 7.03754
R38786 VCC.n11630 VCC.n11629 7.03754
R38787 VCC.n12109 VCC.n12108 7.03754
R38788 VCC.n12165 VCC.n11645 7.03754
R38789 VCC.n12665 VCC.n12248 7.03754
R38790 VCC.n12737 VCC.n12736 7.03754
R38791 VCC.n13216 VCC.n13215 7.03754
R38792 VCC.n13272 VCC.n12752 7.03754
R38793 VCC.n13772 VCC.n13355 7.03754
R38794 VCC.n13844 VCC.n13843 7.03754
R38795 VCC.n14323 VCC.n14322 7.03754
R38796 VCC.n14379 VCC.n13859 7.03754
R38797 VCC.n14879 VCC.n14462 7.03754
R38798 VCC.n14951 VCC.n14950 7.03754
R38799 VCC.n15430 VCC.n15429 7.03754
R38800 VCC.n15486 VCC.n14966 7.03754
R38801 VCC.n15986 VCC.n15569 7.03754
R38802 VCC.n16058 VCC.n16057 7.03754
R38803 VCC.n16537 VCC.n16536 7.03754
R38804 VCC.n16593 VCC.n16073 7.03754
R38805 VCC.n17093 VCC.n16676 7.03754
R38806 VCC.n17165 VCC.n17164 7.03754
R38807 VCC.n17457 VCC.n17456 7.03754
R38808 VCC.n17513 VCC.n17180 7.03754
R38809 VCC.n226 VCC.n181 5.48127
R38810 VCC.n291 VCC.n290 5.48127
R38811 VCC.n337 VCC.n336 5.48127
R38812 VCC.n418 VCC.n417 5.48127
R38813 VCC.n778 VCC.n733 5.48127
R38814 VCC.n843 VCC.n842 5.48127
R38815 VCC.n889 VCC.n888 5.48127
R38816 VCC.n970 VCC.n969 5.48127
R38817 VCC.n1446 VCC.n1445 5.48127
R38818 VCC.n1527 VCC.n1526 5.48127
R38819 VCC.n1336 VCC.n1291 5.48127
R38820 VCC.n1401 VCC.n1400 5.48127
R38821 VCC.n1887 VCC.n1842 5.48127
R38822 VCC.n1952 VCC.n1951 5.48127
R38823 VCC.n1998 VCC.n1997 5.48127
R38824 VCC.n2079 VCC.n2078 5.48127
R38825 VCC.n2555 VCC.n2554 5.48127
R38826 VCC.n2636 VCC.n2635 5.48127
R38827 VCC.n2445 VCC.n2400 5.48127
R38828 VCC.n2510 VCC.n2509 5.48127
R38829 VCC.n2996 VCC.n2951 5.48127
R38830 VCC.n3061 VCC.n3060 5.48127
R38831 VCC.n3107 VCC.n3106 5.48127
R38832 VCC.n3188 VCC.n3187 5.48127
R38833 VCC.n3664 VCC.n3663 5.48127
R38834 VCC.n3745 VCC.n3744 5.48127
R38835 VCC.n3554 VCC.n3509 5.48127
R38836 VCC.n3619 VCC.n3618 5.48127
R38837 VCC.n4105 VCC.n4060 5.48127
R38838 VCC.n4170 VCC.n4169 5.48127
R38839 VCC.n4216 VCC.n4215 5.48127
R38840 VCC.n4297 VCC.n4296 5.48127
R38841 VCC.n4773 VCC.n4772 5.48127
R38842 VCC.n4854 VCC.n4853 5.48127
R38843 VCC.n4663 VCC.n4618 5.48127
R38844 VCC.n4728 VCC.n4727 5.48127
R38845 VCC.n5214 VCC.n5169 5.48127
R38846 VCC.n5279 VCC.n5278 5.48127
R38847 VCC.n5325 VCC.n5324 5.48127
R38848 VCC.n5406 VCC.n5405 5.48127
R38849 VCC.n5882 VCC.n5881 5.48127
R38850 VCC.n5963 VCC.n5962 5.48127
R38851 VCC.n5772 VCC.n5727 5.48127
R38852 VCC.n5837 VCC.n5836 5.48127
R38853 VCC.n6323 VCC.n6278 5.48127
R38854 VCC.n6388 VCC.n6387 5.48127
R38855 VCC.n6434 VCC.n6433 5.48127
R38856 VCC.n6515 VCC.n6514 5.48127
R38857 VCC.n6991 VCC.n6990 5.48127
R38858 VCC.n7072 VCC.n7071 5.48127
R38859 VCC.n6881 VCC.n6836 5.48127
R38860 VCC.n6946 VCC.n6945 5.48127
R38861 VCC.n7432 VCC.n7387 5.48127
R38862 VCC.n7497 VCC.n7496 5.48127
R38863 VCC.n7543 VCC.n7542 5.48127
R38864 VCC.n7624 VCC.n7623 5.48127
R38865 VCC.n8100 VCC.n8099 5.48127
R38866 VCC.n8181 VCC.n8180 5.48127
R38867 VCC.n7990 VCC.n7945 5.48127
R38868 VCC.n8055 VCC.n8054 5.48127
R38869 VCC.n8652 VCC.n8651 5.48127
R38870 VCC.n8733 VCC.n8732 5.48127
R38871 VCC.n8541 VCC.n8496 5.48127
R38872 VCC.n8606 VCC.n8605 5.48127
R38873 VCC.n9209 VCC.n9208 5.48127
R38874 VCC.n9290 VCC.n9289 5.48127
R38875 VCC.n9099 VCC.n9054 5.48127
R38876 VCC.n9164 VCC.n9163 5.48127
R38877 VCC.n9650 VCC.n9605 5.48127
R38878 VCC.n9715 VCC.n9714 5.48127
R38879 VCC.n9761 VCC.n9760 5.48127
R38880 VCC.n9842 VCC.n9841 5.48127
R38881 VCC.n10317 VCC.n10316 5.48127
R38882 VCC.n10398 VCC.n10397 5.48127
R38883 VCC.n10207 VCC.n10162 5.48127
R38884 VCC.n10272 VCC.n10271 5.48127
R38885 VCC.n10757 VCC.n10712 5.48127
R38886 VCC.n10822 VCC.n10821 5.48127
R38887 VCC.n10868 VCC.n10867 5.48127
R38888 VCC.n10949 VCC.n10948 5.48127
R38889 VCC.n11424 VCC.n11423 5.48127
R38890 VCC.n11505 VCC.n11504 5.48127
R38891 VCC.n11314 VCC.n11269 5.48127
R38892 VCC.n11379 VCC.n11378 5.48127
R38893 VCC.n11864 VCC.n11819 5.48127
R38894 VCC.n11929 VCC.n11928 5.48127
R38895 VCC.n11975 VCC.n11974 5.48127
R38896 VCC.n12056 VCC.n12055 5.48127
R38897 VCC.n12531 VCC.n12530 5.48127
R38898 VCC.n12612 VCC.n12611 5.48127
R38899 VCC.n12421 VCC.n12376 5.48127
R38900 VCC.n12486 VCC.n12485 5.48127
R38901 VCC.n12971 VCC.n12926 5.48127
R38902 VCC.n13036 VCC.n13035 5.48127
R38903 VCC.n13082 VCC.n13081 5.48127
R38904 VCC.n13163 VCC.n13162 5.48127
R38905 VCC.n13638 VCC.n13637 5.48127
R38906 VCC.n13719 VCC.n13718 5.48127
R38907 VCC.n13528 VCC.n13483 5.48127
R38908 VCC.n13593 VCC.n13592 5.48127
R38909 VCC.n14078 VCC.n14033 5.48127
R38910 VCC.n14143 VCC.n14142 5.48127
R38911 VCC.n14189 VCC.n14188 5.48127
R38912 VCC.n14270 VCC.n14269 5.48127
R38913 VCC.n14745 VCC.n14744 5.48127
R38914 VCC.n14826 VCC.n14825 5.48127
R38915 VCC.n14635 VCC.n14590 5.48127
R38916 VCC.n14700 VCC.n14699 5.48127
R38917 VCC.n15185 VCC.n15140 5.48127
R38918 VCC.n15250 VCC.n15249 5.48127
R38919 VCC.n15296 VCC.n15295 5.48127
R38920 VCC.n15377 VCC.n15376 5.48127
R38921 VCC.n15852 VCC.n15851 5.48127
R38922 VCC.n15933 VCC.n15932 5.48127
R38923 VCC.n15742 VCC.n15697 5.48127
R38924 VCC.n15807 VCC.n15806 5.48127
R38925 VCC.n16292 VCC.n16247 5.48127
R38926 VCC.n16357 VCC.n16356 5.48127
R38927 VCC.n16403 VCC.n16402 5.48127
R38928 VCC.n16484 VCC.n16483 5.48127
R38929 VCC.n16959 VCC.n16958 5.48127
R38930 VCC.n17040 VCC.n17039 5.48127
R38931 VCC.n16849 VCC.n16804 5.48127
R38932 VCC.n16914 VCC.n16913 5.48127
R38933 VCC.n17323 VCC.n17322 5.48127
R38934 VCC.n17404 VCC.n17403 5.48127
R38935 VCC.n424 VCC.n423 4.88621
R38936 VCC.n976 VCC.n975 4.88621
R38937 VCC.n1534 VCC.n1533 4.88621
R38938 VCC.n2085 VCC.n2084 4.88621
R38939 VCC.n2643 VCC.n2642 4.88621
R38940 VCC.n3194 VCC.n3193 4.88621
R38941 VCC.n3752 VCC.n3751 4.88621
R38942 VCC.n4303 VCC.n4302 4.88621
R38943 VCC.n4861 VCC.n4860 4.88621
R38944 VCC.n5412 VCC.n5411 4.88621
R38945 VCC.n5970 VCC.n5969 4.88621
R38946 VCC.n6521 VCC.n6520 4.88621
R38947 VCC.n7079 VCC.n7078 4.88621
R38948 VCC.n7630 VCC.n7629 4.88621
R38949 VCC.n8188 VCC.n8187 4.88621
R38950 VCC.n8739 VCC.n8738 4.88621
R38951 VCC.n9297 VCC.n9296 4.88621
R38952 VCC.n9848 VCC.n9847 4.88621
R38953 VCC.n10405 VCC.n10404 4.88621
R38954 VCC.n10955 VCC.n10954 4.88621
R38955 VCC.n11512 VCC.n11511 4.88621
R38956 VCC.n12062 VCC.n12061 4.88621
R38957 VCC.n12619 VCC.n12618 4.88621
R38958 VCC.n13169 VCC.n13168 4.88621
R38959 VCC.n13726 VCC.n13725 4.88621
R38960 VCC.n14276 VCC.n14275 4.88621
R38961 VCC.n14833 VCC.n14832 4.88621
R38962 VCC.n15383 VCC.n15382 4.88621
R38963 VCC.n15940 VCC.n15939 4.88621
R38964 VCC.n16490 VCC.n16489 4.88621
R38965 VCC.n17047 VCC.n17046 4.88621
R38966 VCC.n17410 VCC.n17409 4.88621
R38967 VCC.n499 VCC.n39 4.84621
R38968 VCC.n499 VCC.n498 4.84621
R38969 VCC.n1051 VCC.n591 4.84621
R38970 VCC.n1051 VCC.n1050 4.84621
R38971 VCC.n1616 VCC.n1145 4.84621
R38972 VCC.n1617 VCC.n1616 4.84621
R38973 VCC.n2160 VCC.n1700 4.84621
R38974 VCC.n2160 VCC.n2159 4.84621
R38975 VCC.n2725 VCC.n2254 4.84621
R38976 VCC.n2726 VCC.n2725 4.84621
R38977 VCC.n3269 VCC.n2809 4.84621
R38978 VCC.n3269 VCC.n3268 4.84621
R38979 VCC.n3834 VCC.n3363 4.84621
R38980 VCC.n3835 VCC.n3834 4.84621
R38981 VCC.n4378 VCC.n3918 4.84621
R38982 VCC.n4378 VCC.n4377 4.84621
R38983 VCC.n4943 VCC.n4472 4.84621
R38984 VCC.n4944 VCC.n4943 4.84621
R38985 VCC.n5487 VCC.n5027 4.84621
R38986 VCC.n5487 VCC.n5486 4.84621
R38987 VCC.n6052 VCC.n5581 4.84621
R38988 VCC.n6053 VCC.n6052 4.84621
R38989 VCC.n6596 VCC.n6136 4.84621
R38990 VCC.n6596 VCC.n6595 4.84621
R38991 VCC.n7161 VCC.n6690 4.84621
R38992 VCC.n7162 VCC.n7161 4.84621
R38993 VCC.n7705 VCC.n7245 4.84621
R38994 VCC.n7705 VCC.n7704 4.84621
R38995 VCC.n8270 VCC.n7799 4.84621
R38996 VCC.n8271 VCC.n8270 4.84621
R38997 VCC.n8814 VCC.n8354 4.84621
R38998 VCC.n8814 VCC.n8813 4.84621
R38999 VCC.n9379 VCC.n8908 4.84621
R39000 VCC.n9380 VCC.n9379 4.84621
R39001 VCC.n9923 VCC.n9463 4.84621
R39002 VCC.n9923 VCC.n9922 4.84621
R39003 VCC.n10487 VCC.n10016 4.84621
R39004 VCC.n10488 VCC.n10487 4.84621
R39005 VCC.n11030 VCC.n10570 4.84621
R39006 VCC.n11030 VCC.n11029 4.84621
R39007 VCC.n11594 VCC.n11123 4.84621
R39008 VCC.n11595 VCC.n11594 4.84621
R39009 VCC.n12137 VCC.n11677 4.84621
R39010 VCC.n12137 VCC.n12136 4.84621
R39011 VCC.n12701 VCC.n12230 4.84621
R39012 VCC.n12702 VCC.n12701 4.84621
R39013 VCC.n13244 VCC.n12784 4.84621
R39014 VCC.n13244 VCC.n13243 4.84621
R39015 VCC.n13808 VCC.n13337 4.84621
R39016 VCC.n13809 VCC.n13808 4.84621
R39017 VCC.n14351 VCC.n13891 4.84621
R39018 VCC.n14351 VCC.n14350 4.84621
R39019 VCC.n14915 VCC.n14444 4.84621
R39020 VCC.n14916 VCC.n14915 4.84621
R39021 VCC.n15458 VCC.n14998 4.84621
R39022 VCC.n15458 VCC.n15457 4.84621
R39023 VCC.n16022 VCC.n15551 4.84621
R39024 VCC.n16023 VCC.n16022 4.84621
R39025 VCC.n16565 VCC.n16105 4.84621
R39026 VCC.n16565 VCC.n16564 4.84621
R39027 VCC.n17129 VCC.n16658 4.84621
R39028 VCC.n17130 VCC.n17129 4.84621
R39029 VCC.n17485 VCC.n17212 4.84621
R39030 VCC.n17485 VCC.n17484 4.84621
R39031 VCC.n452 VCC.n57 4.6505
R39032 VCC.n1004 VCC.n609 4.6505
R39033 VCC.n1562 VCC.n1165 4.6505
R39034 VCC.n2113 VCC.n1718 4.6505
R39035 VCC.n2671 VCC.n2274 4.6505
R39036 VCC.n3222 VCC.n2827 4.6505
R39037 VCC.n3780 VCC.n3383 4.6505
R39038 VCC.n4331 VCC.n3936 4.6505
R39039 VCC.n4889 VCC.n4492 4.6505
R39040 VCC.n5440 VCC.n5045 4.6505
R39041 VCC.n5998 VCC.n5601 4.6505
R39042 VCC.n6549 VCC.n6154 4.6505
R39043 VCC.n7107 VCC.n6710 4.6505
R39044 VCC.n7658 VCC.n7263 4.6505
R39045 VCC.n8216 VCC.n7819 4.6505
R39046 VCC.n8767 VCC.n8372 4.6505
R39047 VCC.n9325 VCC.n8928 4.6505
R39048 VCC.n9876 VCC.n9481 4.6505
R39049 VCC.n10433 VCC.n10036 4.6505
R39050 VCC.n10983 VCC.n10588 4.6505
R39051 VCC.n11540 VCC.n11143 4.6505
R39052 VCC.n12090 VCC.n11695 4.6505
R39053 VCC.n12647 VCC.n12250 4.6505
R39054 VCC.n13197 VCC.n12802 4.6505
R39055 VCC.n13754 VCC.n13357 4.6505
R39056 VCC.n14304 VCC.n13909 4.6505
R39057 VCC.n14861 VCC.n14464 4.6505
R39058 VCC.n15411 VCC.n15016 4.6505
R39059 VCC.n15968 VCC.n15571 4.6505
R39060 VCC.n16518 VCC.n16123 4.6505
R39061 VCC.n17075 VCC.n16678 4.6505
R39062 VCC.n17438 VCC.n17230 4.6505
R39063 VCC.n215 VCC.n192 4.51211
R39064 VCC.n767 VCC.n744 4.51211
R39065 VCC.n1325 VCC.n1302 4.51211
R39066 VCC.n1876 VCC.n1853 4.51211
R39067 VCC.n2434 VCC.n2411 4.51211
R39068 VCC.n2985 VCC.n2962 4.51211
R39069 VCC.n3543 VCC.n3520 4.51211
R39070 VCC.n4094 VCC.n4071 4.51211
R39071 VCC.n4652 VCC.n4629 4.51211
R39072 VCC.n5203 VCC.n5180 4.51211
R39073 VCC.n5761 VCC.n5738 4.51211
R39074 VCC.n6312 VCC.n6289 4.51211
R39075 VCC.n6870 VCC.n6847 4.51211
R39076 VCC.n7421 VCC.n7398 4.51211
R39077 VCC.n7979 VCC.n7956 4.51211
R39078 VCC.n8530 VCC.n8507 4.51211
R39079 VCC.n9088 VCC.n9065 4.51211
R39080 VCC.n9639 VCC.n9616 4.51211
R39081 VCC.n10196 VCC.n10173 4.51211
R39082 VCC.n10746 VCC.n10723 4.51211
R39083 VCC.n11303 VCC.n11280 4.51211
R39084 VCC.n11853 VCC.n11830 4.51211
R39085 VCC.n12410 VCC.n12387 4.51211
R39086 VCC.n12960 VCC.n12937 4.51211
R39087 VCC.n13517 VCC.n13494 4.51211
R39088 VCC.n14067 VCC.n14044 4.51211
R39089 VCC.n14624 VCC.n14601 4.51211
R39090 VCC.n15174 VCC.n15151 4.51211
R39091 VCC.n15731 VCC.n15708 4.51211
R39092 VCC.n16281 VCC.n16258 4.51211
R39093 VCC.n16838 VCC.n16815 4.51211
R39094 VCC.n314 VCC.n125 4.51121
R39095 VCC.n866 VCC.n677 4.51121
R39096 VCC.n1424 VCC.n1234 4.51121
R39097 VCC.n1975 VCC.n1786 4.51121
R39098 VCC.n2533 VCC.n2343 4.51121
R39099 VCC.n3084 VCC.n2895 4.51121
R39100 VCC.n3642 VCC.n3452 4.51121
R39101 VCC.n4193 VCC.n4004 4.51121
R39102 VCC.n4751 VCC.n4561 4.51121
R39103 VCC.n5302 VCC.n5113 4.51121
R39104 VCC.n5860 VCC.n5670 4.51121
R39105 VCC.n6411 VCC.n6222 4.51121
R39106 VCC.n6969 VCC.n6779 4.51121
R39107 VCC.n7520 VCC.n7331 4.51121
R39108 VCC.n8078 VCC.n7888 4.51121
R39109 VCC.n8629 VCC.n8440 4.51121
R39110 VCC.n9187 VCC.n8997 4.51121
R39111 VCC.n9738 VCC.n9549 4.51121
R39112 VCC.n10295 VCC.n10105 4.51121
R39113 VCC.n10845 VCC.n10656 4.51121
R39114 VCC.n11402 VCC.n11212 4.51121
R39115 VCC.n11952 VCC.n11763 4.51121
R39116 VCC.n12509 VCC.n12319 4.51121
R39117 VCC.n13059 VCC.n12870 4.51121
R39118 VCC.n13616 VCC.n13426 4.51121
R39119 VCC.n14166 VCC.n13977 4.51121
R39120 VCC.n14723 VCC.n14533 4.51121
R39121 VCC.n15273 VCC.n15084 4.51121
R39122 VCC.n15830 VCC.n15640 4.51121
R39123 VCC.n16380 VCC.n16191 4.51121
R39124 VCC.n16937 VCC.n16747 4.51121
R39125 VCC.n17300 VCC.n17298 4.51121
R39126 VCC.n301 VCC.n135 4.5005
R39127 VCC.n300 VCC.n299 4.5005
R39128 VCC.n204 VCC.n203 4.5005
R39129 VCC.n200 VCC.n197 4.5005
R39130 VCC.n236 VCC.n175 4.5005
R39131 VCC.n246 VCC.n245 4.5005
R39132 VCC.n247 VCC.n246 4.5005
R39133 VCC.n199 VCC.n198 4.5005
R39134 VCC.n221 VCC.n174 4.5005
R39135 VCC.n221 VCC.n184 4.5005
R39136 VCC.n206 VCC.n205 4.5005
R39137 VCC.n207 VCC.n206 4.5005
R39138 VCC.n251 VCC.n166 4.5005
R39139 VCC.n251 VCC.n155 4.5005
R39140 VCC.n312 VCC.n311 4.5005
R39141 VCC.n276 VCC.n275 4.5005
R39142 VCC.n274 VCC.n146 4.5005
R39143 VCC.n254 VCC.n167 4.5005
R39144 VCC.n262 VCC.n261 4.5005
R39145 VCC.n263 VCC.n262 4.5005
R39146 VCC.n158 VCC.n148 4.5005
R39147 VCC.n159 VCC.n158 4.5005
R39148 VCC.n284 VCC.n283 4.5005
R39149 VCC.n285 VCC.n284 4.5005
R39150 VCC.n303 VCC.n302 4.5005
R39151 VCC.n138 VCC.n136 4.5005
R39152 VCC.n296 VCC.n138 4.5005
R39153 VCC.n239 VCC.n238 4.5005
R39154 VCC.n436 VCC.n74 4.5005
R39155 VCC.n435 VCC.n434 4.5005
R39156 VCC.n329 VCC.n328 4.5005
R39157 VCC.n324 VCC.n321 4.5005
R39158 VCC.n353 VCC.n352 4.5005
R39159 VCC.n323 VCC.n322 4.5005
R39160 VCC.n447 VCC.n446 4.5005
R39161 VCC.n403 VCC.n402 4.5005
R39162 VCC.n401 VCC.n86 4.5005
R39163 VCC.n438 VCC.n437 4.5005
R39164 VCC.n355 VCC.n354 4.5005
R39165 VCC.n368 VCC.n367 4.5005
R39166 VCC.n367 VCC.n366 4.5005
R39167 VCC.n117 VCC.n113 4.5005
R39168 VCC.n340 VCC.n117 4.5005
R39169 VCC.n331 VCC.n330 4.5005
R39170 VCC.n331 VCC.n124 4.5005
R39171 VCC.n383 VCC.n382 4.5005
R39172 VCC.n384 VCC.n383 4.5005
R39173 VCC.n375 VCC.n96 4.5005
R39174 VCC.n386 VCC.n96 4.5005
R39175 VCC.n390 VCC.n88 4.5005
R39176 VCC.n391 VCC.n390 4.5005
R39177 VCC.n411 VCC.n410 4.5005
R39178 VCC.n412 VCC.n411 4.5005
R39179 VCC.n77 VCC.n75 4.5005
R39180 VCC.n431 VCC.n77 4.5005
R39181 VCC.n540 VCC.n9 4.5005
R39182 VCC.n542 VCC.n541 4.5005
R39183 VCC.n519 VCC.n27 4.5005
R39184 VCC.n53 VCC.n51 4.5005
R39185 VCC.n60 VCC.n58 4.5005
R39186 VCC.n451 VCC.n450 4.5005
R39187 VCC.n456 VCC.n455 4.5005
R39188 VCC.n462 VCC.n50 4.5005
R39189 VCC.n48 VCC.n47 4.5005
R39190 VCC.n518 VCC.n517 4.5005
R39191 VCC.n509 VCC.n31 4.5005
R39192 VCC.n521 VCC.n520 4.5005
R39193 VCC.n521 VCC.n25 4.5005
R39194 VCC.n29 VCC.n16 4.5005
R39195 VCC.n17 VCC.n10 4.5005
R39196 VCC.n19 VCC.n18 4.5005
R39197 VCC.n530 VCC.n19 4.5005
R39198 VCC.n508 VCC.n507 4.5005
R39199 VCC.n38 VCC.n36 4.5005
R39200 VCC.n46 VCC.n44 4.5005
R39201 VCC.n44 VCC.n43 4.5005
R39202 VCC.n479 VCC.n478 4.5005
R39203 VCC.n467 VCC.n466 4.5005
R39204 VCC.n454 VCC.n453 4.5005
R39205 VCC.n551 VCC.n550 4.5005
R39206 VCC.n853 VCC.n687 4.5005
R39207 VCC.n852 VCC.n851 4.5005
R39208 VCC.n756 VCC.n755 4.5005
R39209 VCC.n752 VCC.n749 4.5005
R39210 VCC.n788 VCC.n727 4.5005
R39211 VCC.n798 VCC.n797 4.5005
R39212 VCC.n799 VCC.n798 4.5005
R39213 VCC.n751 VCC.n750 4.5005
R39214 VCC.n773 VCC.n726 4.5005
R39215 VCC.n773 VCC.n736 4.5005
R39216 VCC.n758 VCC.n757 4.5005
R39217 VCC.n759 VCC.n758 4.5005
R39218 VCC.n803 VCC.n718 4.5005
R39219 VCC.n803 VCC.n707 4.5005
R39220 VCC.n864 VCC.n863 4.5005
R39221 VCC.n828 VCC.n827 4.5005
R39222 VCC.n826 VCC.n698 4.5005
R39223 VCC.n806 VCC.n719 4.5005
R39224 VCC.n814 VCC.n813 4.5005
R39225 VCC.n815 VCC.n814 4.5005
R39226 VCC.n710 VCC.n700 4.5005
R39227 VCC.n711 VCC.n710 4.5005
R39228 VCC.n836 VCC.n835 4.5005
R39229 VCC.n837 VCC.n836 4.5005
R39230 VCC.n855 VCC.n854 4.5005
R39231 VCC.n690 VCC.n688 4.5005
R39232 VCC.n848 VCC.n690 4.5005
R39233 VCC.n791 VCC.n790 4.5005
R39234 VCC.n988 VCC.n626 4.5005
R39235 VCC.n987 VCC.n986 4.5005
R39236 VCC.n881 VCC.n880 4.5005
R39237 VCC.n876 VCC.n873 4.5005
R39238 VCC.n905 VCC.n904 4.5005
R39239 VCC.n875 VCC.n874 4.5005
R39240 VCC.n999 VCC.n998 4.5005
R39241 VCC.n955 VCC.n954 4.5005
R39242 VCC.n953 VCC.n638 4.5005
R39243 VCC.n990 VCC.n989 4.5005
R39244 VCC.n907 VCC.n906 4.5005
R39245 VCC.n920 VCC.n919 4.5005
R39246 VCC.n919 VCC.n918 4.5005
R39247 VCC.n669 VCC.n665 4.5005
R39248 VCC.n892 VCC.n669 4.5005
R39249 VCC.n883 VCC.n882 4.5005
R39250 VCC.n883 VCC.n676 4.5005
R39251 VCC.n935 VCC.n934 4.5005
R39252 VCC.n936 VCC.n935 4.5005
R39253 VCC.n927 VCC.n648 4.5005
R39254 VCC.n938 VCC.n648 4.5005
R39255 VCC.n942 VCC.n640 4.5005
R39256 VCC.n943 VCC.n942 4.5005
R39257 VCC.n963 VCC.n962 4.5005
R39258 VCC.n964 VCC.n963 4.5005
R39259 VCC.n629 VCC.n627 4.5005
R39260 VCC.n983 VCC.n629 4.5005
R39261 VCC.n569 VCC.n564 4.5005
R39262 VCC.n1096 VCC.n1095 4.5005
R39263 VCC.n1006 VCC.n1005 4.5005
R39264 VCC.n612 VCC.n610 4.5005
R39265 VCC.n1031 VCC.n1030 4.5005
R39266 VCC.n598 VCC.n596 4.5005
R39267 VCC.n596 VCC.n595 4.5005
R39268 VCC.n600 VCC.n599 4.5005
R39269 VCC.n1014 VCC.n602 4.5005
R39270 VCC.n1019 VCC.n1018 4.5005
R39271 VCC.n1003 VCC.n1002 4.5005
R39272 VCC.n1008 VCC.n1007 4.5005
R39273 VCC.n571 VCC.n570 4.5005
R39274 VCC.n1082 VCC.n571 4.5005
R39275 VCC.n1070 VCC.n1069 4.5005
R39276 VCC.n581 VCC.n568 4.5005
R39277 VCC.n1060 VCC.n1059 4.5005
R39278 VCC.n590 VCC.n588 4.5005
R39279 VCC.n1061 VCC.n583 4.5005
R39280 VCC.n1071 VCC.n579 4.5005
R39281 VCC.n1073 VCC.n1072 4.5005
R39282 VCC.n1073 VCC.n577 4.5005
R39283 VCC.n1094 VCC.n563 4.5005
R39284 VCC.n1105 VCC.n1104 4.5005
R39285 VCC.n605 VCC.n603 4.5005
R39286 VCC.n1564 VCC.n1166 4.5005
R39287 VCC.n1567 VCC.n1566 4.5005
R39288 VCC.n1641 VCC.n1121 4.5005
R39289 VCC.n1643 VCC.n1642 4.5005
R39290 VCC.n1138 VCC.n1137 4.5005
R39291 VCC.n1158 VCC.n1156 4.5005
R39292 VCC.n1168 VCC.n1155 4.5005
R39293 VCC.n1597 VCC.n1596 4.5005
R39294 VCC.n1606 VCC.n1605 4.5005
R39295 VCC.n1149 VCC.n1148 4.5005
R39296 VCC.n1129 VCC.n1128 4.5005
R39297 VCC.n1632 VCC.n1631 4.5005
R39298 VCC.n1644 VCC.n1119 4.5005
R39299 VCC.n1133 VCC.n1131 4.5005
R39300 VCC.n1604 VCC.n1603 4.5005
R39301 VCC.n1565 VCC.n1563 4.5005
R39302 VCC.n1561 VCC.n1560 4.5005
R39303 VCC.n1576 VCC.n1167 4.5005
R39304 VCC.n1646 VCC.n1645 4.5005
R39305 VCC.n1646 VCC.n1117 4.5005
R39306 VCC.n1136 VCC.n1134 4.5005
R39307 VCC.n1141 VCC.n1134 4.5005
R39308 VCC.n1592 VCC.n1591 4.5005
R39309 VCC.n1593 VCC.n1592 4.5005
R39310 VCC.n1659 VCC.n1658 4.5005
R39311 VCC.n1546 VCC.n1183 4.5005
R39312 VCC.n1545 VCC.n1544 4.5005
R39313 VCC.n1510 VCC.n1195 4.5005
R39314 VCC.n1464 VCC.n1463 4.5005
R39315 VCC.n1438 VCC.n1437 4.5005
R39316 VCC.n1433 VCC.n1429 4.5005
R39317 VCC.n1439 VCC.n1235 4.5005
R39318 VCC.n1235 VCC.n1233 4.5005
R39319 VCC.n1557 VCC.n1556 4.5005
R39320 VCC.n1512 VCC.n1511 4.5005
R39321 VCC.n1432 VCC.n1431 4.5005
R39322 VCC.n1226 VCC.n1222 4.5005
R39323 VCC.n1449 VCC.n1226 4.5005
R39324 VCC.n1462 VCC.n1461 4.5005
R39325 VCC.n1477 VCC.n1476 4.5005
R39326 VCC.n1476 VCC.n1475 4.5005
R39327 VCC.n1492 VCC.n1491 4.5005
R39328 VCC.n1493 VCC.n1492 4.5005
R39329 VCC.n1484 VCC.n1205 4.5005
R39330 VCC.n1495 VCC.n1205 4.5005
R39331 VCC.n1499 VCC.n1197 4.5005
R39332 VCC.n1500 VCC.n1499 4.5005
R39333 VCC.n1520 VCC.n1519 4.5005
R39334 VCC.n1521 VCC.n1520 4.5005
R39335 VCC.n1548 VCC.n1547 4.5005
R39336 VCC.n1186 VCC.n1184 4.5005
R39337 VCC.n1541 VCC.n1186 4.5005
R39338 VCC.n1411 VCC.n1245 4.5005
R39339 VCC.n1410 VCC.n1409 4.5005
R39340 VCC.n1384 VCC.n1256 4.5005
R39341 VCC.n1349 VCC.n1348 4.5005
R39342 VCC.n1314 VCC.n1313 4.5005
R39343 VCC.n1310 VCC.n1307 4.5005
R39344 VCC.n1316 VCC.n1315 4.5005
R39345 VCC.n1317 VCC.n1316 4.5005
R39346 VCC.n1422 VCC.n1421 4.5005
R39347 VCC.n1386 VCC.n1385 4.5005
R39348 VCC.n1309 VCC.n1308 4.5005
R39349 VCC.n1331 VCC.n1284 4.5005
R39350 VCC.n1331 VCC.n1294 4.5005
R39351 VCC.n1346 VCC.n1285 4.5005
R39352 VCC.n1356 VCC.n1355 4.5005
R39353 VCC.n1357 VCC.n1356 4.5005
R39354 VCC.n1361 VCC.n1276 4.5005
R39355 VCC.n1361 VCC.n1265 4.5005
R39356 VCC.n1364 VCC.n1277 4.5005
R39357 VCC.n1372 VCC.n1371 4.5005
R39358 VCC.n1373 VCC.n1372 4.5005
R39359 VCC.n1268 VCC.n1258 4.5005
R39360 VCC.n1269 VCC.n1268 4.5005
R39361 VCC.n1394 VCC.n1393 4.5005
R39362 VCC.n1395 VCC.n1394 4.5005
R39363 VCC.n1413 VCC.n1412 4.5005
R39364 VCC.n1248 VCC.n1246 4.5005
R39365 VCC.n1406 VCC.n1248 4.5005
R39366 VCC.n1962 VCC.n1796 4.5005
R39367 VCC.n1961 VCC.n1960 4.5005
R39368 VCC.n1865 VCC.n1864 4.5005
R39369 VCC.n1861 VCC.n1858 4.5005
R39370 VCC.n1897 VCC.n1836 4.5005
R39371 VCC.n1907 VCC.n1906 4.5005
R39372 VCC.n1908 VCC.n1907 4.5005
R39373 VCC.n1860 VCC.n1859 4.5005
R39374 VCC.n1882 VCC.n1835 4.5005
R39375 VCC.n1882 VCC.n1845 4.5005
R39376 VCC.n1867 VCC.n1866 4.5005
R39377 VCC.n1868 VCC.n1867 4.5005
R39378 VCC.n1912 VCC.n1827 4.5005
R39379 VCC.n1912 VCC.n1816 4.5005
R39380 VCC.n1973 VCC.n1972 4.5005
R39381 VCC.n1937 VCC.n1936 4.5005
R39382 VCC.n1935 VCC.n1807 4.5005
R39383 VCC.n1915 VCC.n1828 4.5005
R39384 VCC.n1923 VCC.n1922 4.5005
R39385 VCC.n1924 VCC.n1923 4.5005
R39386 VCC.n1819 VCC.n1809 4.5005
R39387 VCC.n1820 VCC.n1819 4.5005
R39388 VCC.n1945 VCC.n1944 4.5005
R39389 VCC.n1946 VCC.n1945 4.5005
R39390 VCC.n1964 VCC.n1963 4.5005
R39391 VCC.n1799 VCC.n1797 4.5005
R39392 VCC.n1957 VCC.n1799 4.5005
R39393 VCC.n1900 VCC.n1899 4.5005
R39394 VCC.n2097 VCC.n1735 4.5005
R39395 VCC.n2096 VCC.n2095 4.5005
R39396 VCC.n1990 VCC.n1989 4.5005
R39397 VCC.n1985 VCC.n1982 4.5005
R39398 VCC.n2014 VCC.n2013 4.5005
R39399 VCC.n1984 VCC.n1983 4.5005
R39400 VCC.n2108 VCC.n2107 4.5005
R39401 VCC.n2064 VCC.n2063 4.5005
R39402 VCC.n2062 VCC.n1747 4.5005
R39403 VCC.n2099 VCC.n2098 4.5005
R39404 VCC.n2016 VCC.n2015 4.5005
R39405 VCC.n2029 VCC.n2028 4.5005
R39406 VCC.n2028 VCC.n2027 4.5005
R39407 VCC.n1778 VCC.n1774 4.5005
R39408 VCC.n2001 VCC.n1778 4.5005
R39409 VCC.n1992 VCC.n1991 4.5005
R39410 VCC.n1992 VCC.n1785 4.5005
R39411 VCC.n2044 VCC.n2043 4.5005
R39412 VCC.n2045 VCC.n2044 4.5005
R39413 VCC.n2036 VCC.n1757 4.5005
R39414 VCC.n2047 VCC.n1757 4.5005
R39415 VCC.n2051 VCC.n1749 4.5005
R39416 VCC.n2052 VCC.n2051 4.5005
R39417 VCC.n2072 VCC.n2071 4.5005
R39418 VCC.n2073 VCC.n2072 4.5005
R39419 VCC.n1738 VCC.n1736 4.5005
R39420 VCC.n2092 VCC.n1738 4.5005
R39421 VCC.n1678 VCC.n1673 4.5005
R39422 VCC.n2205 VCC.n2204 4.5005
R39423 VCC.n2115 VCC.n2114 4.5005
R39424 VCC.n1721 VCC.n1719 4.5005
R39425 VCC.n2140 VCC.n2139 4.5005
R39426 VCC.n1707 VCC.n1705 4.5005
R39427 VCC.n1705 VCC.n1704 4.5005
R39428 VCC.n1709 VCC.n1708 4.5005
R39429 VCC.n2123 VCC.n1711 4.5005
R39430 VCC.n2128 VCC.n2127 4.5005
R39431 VCC.n2112 VCC.n2111 4.5005
R39432 VCC.n2117 VCC.n2116 4.5005
R39433 VCC.n1680 VCC.n1679 4.5005
R39434 VCC.n2191 VCC.n1680 4.5005
R39435 VCC.n2179 VCC.n2178 4.5005
R39436 VCC.n1690 VCC.n1677 4.5005
R39437 VCC.n2169 VCC.n2168 4.5005
R39438 VCC.n1699 VCC.n1697 4.5005
R39439 VCC.n2170 VCC.n1692 4.5005
R39440 VCC.n2180 VCC.n1688 4.5005
R39441 VCC.n2182 VCC.n2181 4.5005
R39442 VCC.n2182 VCC.n1686 4.5005
R39443 VCC.n2203 VCC.n1672 4.5005
R39444 VCC.n2214 VCC.n2213 4.5005
R39445 VCC.n1714 VCC.n1712 4.5005
R39446 VCC.n2673 VCC.n2275 4.5005
R39447 VCC.n2676 VCC.n2675 4.5005
R39448 VCC.n2750 VCC.n2230 4.5005
R39449 VCC.n2752 VCC.n2751 4.5005
R39450 VCC.n2247 VCC.n2246 4.5005
R39451 VCC.n2267 VCC.n2265 4.5005
R39452 VCC.n2277 VCC.n2264 4.5005
R39453 VCC.n2706 VCC.n2705 4.5005
R39454 VCC.n2715 VCC.n2714 4.5005
R39455 VCC.n2258 VCC.n2257 4.5005
R39456 VCC.n2238 VCC.n2237 4.5005
R39457 VCC.n2741 VCC.n2740 4.5005
R39458 VCC.n2753 VCC.n2228 4.5005
R39459 VCC.n2242 VCC.n2240 4.5005
R39460 VCC.n2713 VCC.n2712 4.5005
R39461 VCC.n2674 VCC.n2672 4.5005
R39462 VCC.n2670 VCC.n2669 4.5005
R39463 VCC.n2685 VCC.n2276 4.5005
R39464 VCC.n2755 VCC.n2754 4.5005
R39465 VCC.n2755 VCC.n2226 4.5005
R39466 VCC.n2245 VCC.n2243 4.5005
R39467 VCC.n2250 VCC.n2243 4.5005
R39468 VCC.n2701 VCC.n2700 4.5005
R39469 VCC.n2702 VCC.n2701 4.5005
R39470 VCC.n2768 VCC.n2767 4.5005
R39471 VCC.n2655 VCC.n2292 4.5005
R39472 VCC.n2654 VCC.n2653 4.5005
R39473 VCC.n2619 VCC.n2304 4.5005
R39474 VCC.n2573 VCC.n2572 4.5005
R39475 VCC.n2547 VCC.n2546 4.5005
R39476 VCC.n2542 VCC.n2538 4.5005
R39477 VCC.n2548 VCC.n2344 4.5005
R39478 VCC.n2344 VCC.n2342 4.5005
R39479 VCC.n2666 VCC.n2665 4.5005
R39480 VCC.n2621 VCC.n2620 4.5005
R39481 VCC.n2541 VCC.n2540 4.5005
R39482 VCC.n2335 VCC.n2331 4.5005
R39483 VCC.n2558 VCC.n2335 4.5005
R39484 VCC.n2571 VCC.n2570 4.5005
R39485 VCC.n2586 VCC.n2585 4.5005
R39486 VCC.n2585 VCC.n2584 4.5005
R39487 VCC.n2601 VCC.n2600 4.5005
R39488 VCC.n2602 VCC.n2601 4.5005
R39489 VCC.n2593 VCC.n2314 4.5005
R39490 VCC.n2604 VCC.n2314 4.5005
R39491 VCC.n2608 VCC.n2306 4.5005
R39492 VCC.n2609 VCC.n2608 4.5005
R39493 VCC.n2629 VCC.n2628 4.5005
R39494 VCC.n2630 VCC.n2629 4.5005
R39495 VCC.n2657 VCC.n2656 4.5005
R39496 VCC.n2295 VCC.n2293 4.5005
R39497 VCC.n2650 VCC.n2295 4.5005
R39498 VCC.n2520 VCC.n2354 4.5005
R39499 VCC.n2519 VCC.n2518 4.5005
R39500 VCC.n2493 VCC.n2365 4.5005
R39501 VCC.n2458 VCC.n2457 4.5005
R39502 VCC.n2423 VCC.n2422 4.5005
R39503 VCC.n2419 VCC.n2416 4.5005
R39504 VCC.n2425 VCC.n2424 4.5005
R39505 VCC.n2426 VCC.n2425 4.5005
R39506 VCC.n2531 VCC.n2530 4.5005
R39507 VCC.n2495 VCC.n2494 4.5005
R39508 VCC.n2418 VCC.n2417 4.5005
R39509 VCC.n2440 VCC.n2393 4.5005
R39510 VCC.n2440 VCC.n2403 4.5005
R39511 VCC.n2455 VCC.n2394 4.5005
R39512 VCC.n2465 VCC.n2464 4.5005
R39513 VCC.n2466 VCC.n2465 4.5005
R39514 VCC.n2470 VCC.n2385 4.5005
R39515 VCC.n2470 VCC.n2374 4.5005
R39516 VCC.n2473 VCC.n2386 4.5005
R39517 VCC.n2481 VCC.n2480 4.5005
R39518 VCC.n2482 VCC.n2481 4.5005
R39519 VCC.n2377 VCC.n2367 4.5005
R39520 VCC.n2378 VCC.n2377 4.5005
R39521 VCC.n2503 VCC.n2502 4.5005
R39522 VCC.n2504 VCC.n2503 4.5005
R39523 VCC.n2522 VCC.n2521 4.5005
R39524 VCC.n2357 VCC.n2355 4.5005
R39525 VCC.n2515 VCC.n2357 4.5005
R39526 VCC.n3071 VCC.n2905 4.5005
R39527 VCC.n3070 VCC.n3069 4.5005
R39528 VCC.n2974 VCC.n2973 4.5005
R39529 VCC.n2970 VCC.n2967 4.5005
R39530 VCC.n3006 VCC.n2945 4.5005
R39531 VCC.n3016 VCC.n3015 4.5005
R39532 VCC.n3017 VCC.n3016 4.5005
R39533 VCC.n2969 VCC.n2968 4.5005
R39534 VCC.n2991 VCC.n2944 4.5005
R39535 VCC.n2991 VCC.n2954 4.5005
R39536 VCC.n2976 VCC.n2975 4.5005
R39537 VCC.n2977 VCC.n2976 4.5005
R39538 VCC.n3021 VCC.n2936 4.5005
R39539 VCC.n3021 VCC.n2925 4.5005
R39540 VCC.n3082 VCC.n3081 4.5005
R39541 VCC.n3046 VCC.n3045 4.5005
R39542 VCC.n3044 VCC.n2916 4.5005
R39543 VCC.n3024 VCC.n2937 4.5005
R39544 VCC.n3032 VCC.n3031 4.5005
R39545 VCC.n3033 VCC.n3032 4.5005
R39546 VCC.n2928 VCC.n2918 4.5005
R39547 VCC.n2929 VCC.n2928 4.5005
R39548 VCC.n3054 VCC.n3053 4.5005
R39549 VCC.n3055 VCC.n3054 4.5005
R39550 VCC.n3073 VCC.n3072 4.5005
R39551 VCC.n2908 VCC.n2906 4.5005
R39552 VCC.n3066 VCC.n2908 4.5005
R39553 VCC.n3009 VCC.n3008 4.5005
R39554 VCC.n3206 VCC.n2844 4.5005
R39555 VCC.n3205 VCC.n3204 4.5005
R39556 VCC.n3099 VCC.n3098 4.5005
R39557 VCC.n3094 VCC.n3091 4.5005
R39558 VCC.n3123 VCC.n3122 4.5005
R39559 VCC.n3093 VCC.n3092 4.5005
R39560 VCC.n3217 VCC.n3216 4.5005
R39561 VCC.n3173 VCC.n3172 4.5005
R39562 VCC.n3171 VCC.n2856 4.5005
R39563 VCC.n3208 VCC.n3207 4.5005
R39564 VCC.n3125 VCC.n3124 4.5005
R39565 VCC.n3138 VCC.n3137 4.5005
R39566 VCC.n3137 VCC.n3136 4.5005
R39567 VCC.n2887 VCC.n2883 4.5005
R39568 VCC.n3110 VCC.n2887 4.5005
R39569 VCC.n3101 VCC.n3100 4.5005
R39570 VCC.n3101 VCC.n2894 4.5005
R39571 VCC.n3153 VCC.n3152 4.5005
R39572 VCC.n3154 VCC.n3153 4.5005
R39573 VCC.n3145 VCC.n2866 4.5005
R39574 VCC.n3156 VCC.n2866 4.5005
R39575 VCC.n3160 VCC.n2858 4.5005
R39576 VCC.n3161 VCC.n3160 4.5005
R39577 VCC.n3181 VCC.n3180 4.5005
R39578 VCC.n3182 VCC.n3181 4.5005
R39579 VCC.n2847 VCC.n2845 4.5005
R39580 VCC.n3201 VCC.n2847 4.5005
R39581 VCC.n2787 VCC.n2782 4.5005
R39582 VCC.n3314 VCC.n3313 4.5005
R39583 VCC.n3224 VCC.n3223 4.5005
R39584 VCC.n2830 VCC.n2828 4.5005
R39585 VCC.n3249 VCC.n3248 4.5005
R39586 VCC.n2816 VCC.n2814 4.5005
R39587 VCC.n2814 VCC.n2813 4.5005
R39588 VCC.n2818 VCC.n2817 4.5005
R39589 VCC.n3232 VCC.n2820 4.5005
R39590 VCC.n3237 VCC.n3236 4.5005
R39591 VCC.n3221 VCC.n3220 4.5005
R39592 VCC.n3226 VCC.n3225 4.5005
R39593 VCC.n2789 VCC.n2788 4.5005
R39594 VCC.n3300 VCC.n2789 4.5005
R39595 VCC.n3288 VCC.n3287 4.5005
R39596 VCC.n2799 VCC.n2786 4.5005
R39597 VCC.n3278 VCC.n3277 4.5005
R39598 VCC.n2808 VCC.n2806 4.5005
R39599 VCC.n3279 VCC.n2801 4.5005
R39600 VCC.n3289 VCC.n2797 4.5005
R39601 VCC.n3291 VCC.n3290 4.5005
R39602 VCC.n3291 VCC.n2795 4.5005
R39603 VCC.n3312 VCC.n2781 4.5005
R39604 VCC.n3323 VCC.n3322 4.5005
R39605 VCC.n2823 VCC.n2821 4.5005
R39606 VCC.n3782 VCC.n3384 4.5005
R39607 VCC.n3785 VCC.n3784 4.5005
R39608 VCC.n3859 VCC.n3339 4.5005
R39609 VCC.n3861 VCC.n3860 4.5005
R39610 VCC.n3356 VCC.n3355 4.5005
R39611 VCC.n3376 VCC.n3374 4.5005
R39612 VCC.n3386 VCC.n3373 4.5005
R39613 VCC.n3815 VCC.n3814 4.5005
R39614 VCC.n3824 VCC.n3823 4.5005
R39615 VCC.n3367 VCC.n3366 4.5005
R39616 VCC.n3347 VCC.n3346 4.5005
R39617 VCC.n3850 VCC.n3849 4.5005
R39618 VCC.n3862 VCC.n3337 4.5005
R39619 VCC.n3351 VCC.n3349 4.5005
R39620 VCC.n3822 VCC.n3821 4.5005
R39621 VCC.n3783 VCC.n3781 4.5005
R39622 VCC.n3779 VCC.n3778 4.5005
R39623 VCC.n3794 VCC.n3385 4.5005
R39624 VCC.n3864 VCC.n3863 4.5005
R39625 VCC.n3864 VCC.n3335 4.5005
R39626 VCC.n3354 VCC.n3352 4.5005
R39627 VCC.n3359 VCC.n3352 4.5005
R39628 VCC.n3810 VCC.n3809 4.5005
R39629 VCC.n3811 VCC.n3810 4.5005
R39630 VCC.n3877 VCC.n3876 4.5005
R39631 VCC.n3764 VCC.n3401 4.5005
R39632 VCC.n3763 VCC.n3762 4.5005
R39633 VCC.n3728 VCC.n3413 4.5005
R39634 VCC.n3682 VCC.n3681 4.5005
R39635 VCC.n3656 VCC.n3655 4.5005
R39636 VCC.n3651 VCC.n3647 4.5005
R39637 VCC.n3657 VCC.n3453 4.5005
R39638 VCC.n3453 VCC.n3451 4.5005
R39639 VCC.n3775 VCC.n3774 4.5005
R39640 VCC.n3730 VCC.n3729 4.5005
R39641 VCC.n3650 VCC.n3649 4.5005
R39642 VCC.n3444 VCC.n3440 4.5005
R39643 VCC.n3667 VCC.n3444 4.5005
R39644 VCC.n3680 VCC.n3679 4.5005
R39645 VCC.n3695 VCC.n3694 4.5005
R39646 VCC.n3694 VCC.n3693 4.5005
R39647 VCC.n3710 VCC.n3709 4.5005
R39648 VCC.n3711 VCC.n3710 4.5005
R39649 VCC.n3702 VCC.n3423 4.5005
R39650 VCC.n3713 VCC.n3423 4.5005
R39651 VCC.n3717 VCC.n3415 4.5005
R39652 VCC.n3718 VCC.n3717 4.5005
R39653 VCC.n3738 VCC.n3737 4.5005
R39654 VCC.n3739 VCC.n3738 4.5005
R39655 VCC.n3766 VCC.n3765 4.5005
R39656 VCC.n3404 VCC.n3402 4.5005
R39657 VCC.n3759 VCC.n3404 4.5005
R39658 VCC.n3629 VCC.n3463 4.5005
R39659 VCC.n3628 VCC.n3627 4.5005
R39660 VCC.n3602 VCC.n3474 4.5005
R39661 VCC.n3567 VCC.n3566 4.5005
R39662 VCC.n3532 VCC.n3531 4.5005
R39663 VCC.n3528 VCC.n3525 4.5005
R39664 VCC.n3534 VCC.n3533 4.5005
R39665 VCC.n3535 VCC.n3534 4.5005
R39666 VCC.n3640 VCC.n3639 4.5005
R39667 VCC.n3604 VCC.n3603 4.5005
R39668 VCC.n3527 VCC.n3526 4.5005
R39669 VCC.n3549 VCC.n3502 4.5005
R39670 VCC.n3549 VCC.n3512 4.5005
R39671 VCC.n3564 VCC.n3503 4.5005
R39672 VCC.n3574 VCC.n3573 4.5005
R39673 VCC.n3575 VCC.n3574 4.5005
R39674 VCC.n3579 VCC.n3494 4.5005
R39675 VCC.n3579 VCC.n3483 4.5005
R39676 VCC.n3582 VCC.n3495 4.5005
R39677 VCC.n3590 VCC.n3589 4.5005
R39678 VCC.n3591 VCC.n3590 4.5005
R39679 VCC.n3486 VCC.n3476 4.5005
R39680 VCC.n3487 VCC.n3486 4.5005
R39681 VCC.n3612 VCC.n3611 4.5005
R39682 VCC.n3613 VCC.n3612 4.5005
R39683 VCC.n3631 VCC.n3630 4.5005
R39684 VCC.n3466 VCC.n3464 4.5005
R39685 VCC.n3624 VCC.n3466 4.5005
R39686 VCC.n4180 VCC.n4014 4.5005
R39687 VCC.n4179 VCC.n4178 4.5005
R39688 VCC.n4083 VCC.n4082 4.5005
R39689 VCC.n4079 VCC.n4076 4.5005
R39690 VCC.n4115 VCC.n4054 4.5005
R39691 VCC.n4125 VCC.n4124 4.5005
R39692 VCC.n4126 VCC.n4125 4.5005
R39693 VCC.n4078 VCC.n4077 4.5005
R39694 VCC.n4100 VCC.n4053 4.5005
R39695 VCC.n4100 VCC.n4063 4.5005
R39696 VCC.n4085 VCC.n4084 4.5005
R39697 VCC.n4086 VCC.n4085 4.5005
R39698 VCC.n4130 VCC.n4045 4.5005
R39699 VCC.n4130 VCC.n4034 4.5005
R39700 VCC.n4191 VCC.n4190 4.5005
R39701 VCC.n4155 VCC.n4154 4.5005
R39702 VCC.n4153 VCC.n4025 4.5005
R39703 VCC.n4133 VCC.n4046 4.5005
R39704 VCC.n4141 VCC.n4140 4.5005
R39705 VCC.n4142 VCC.n4141 4.5005
R39706 VCC.n4037 VCC.n4027 4.5005
R39707 VCC.n4038 VCC.n4037 4.5005
R39708 VCC.n4163 VCC.n4162 4.5005
R39709 VCC.n4164 VCC.n4163 4.5005
R39710 VCC.n4182 VCC.n4181 4.5005
R39711 VCC.n4017 VCC.n4015 4.5005
R39712 VCC.n4175 VCC.n4017 4.5005
R39713 VCC.n4118 VCC.n4117 4.5005
R39714 VCC.n4315 VCC.n3953 4.5005
R39715 VCC.n4314 VCC.n4313 4.5005
R39716 VCC.n4208 VCC.n4207 4.5005
R39717 VCC.n4203 VCC.n4200 4.5005
R39718 VCC.n4232 VCC.n4231 4.5005
R39719 VCC.n4202 VCC.n4201 4.5005
R39720 VCC.n4326 VCC.n4325 4.5005
R39721 VCC.n4282 VCC.n4281 4.5005
R39722 VCC.n4280 VCC.n3965 4.5005
R39723 VCC.n4317 VCC.n4316 4.5005
R39724 VCC.n4234 VCC.n4233 4.5005
R39725 VCC.n4247 VCC.n4246 4.5005
R39726 VCC.n4246 VCC.n4245 4.5005
R39727 VCC.n3996 VCC.n3992 4.5005
R39728 VCC.n4219 VCC.n3996 4.5005
R39729 VCC.n4210 VCC.n4209 4.5005
R39730 VCC.n4210 VCC.n4003 4.5005
R39731 VCC.n4262 VCC.n4261 4.5005
R39732 VCC.n4263 VCC.n4262 4.5005
R39733 VCC.n4254 VCC.n3975 4.5005
R39734 VCC.n4265 VCC.n3975 4.5005
R39735 VCC.n4269 VCC.n3967 4.5005
R39736 VCC.n4270 VCC.n4269 4.5005
R39737 VCC.n4290 VCC.n4289 4.5005
R39738 VCC.n4291 VCC.n4290 4.5005
R39739 VCC.n3956 VCC.n3954 4.5005
R39740 VCC.n4310 VCC.n3956 4.5005
R39741 VCC.n3896 VCC.n3891 4.5005
R39742 VCC.n4423 VCC.n4422 4.5005
R39743 VCC.n4333 VCC.n4332 4.5005
R39744 VCC.n3939 VCC.n3937 4.5005
R39745 VCC.n4358 VCC.n4357 4.5005
R39746 VCC.n3925 VCC.n3923 4.5005
R39747 VCC.n3923 VCC.n3922 4.5005
R39748 VCC.n3927 VCC.n3926 4.5005
R39749 VCC.n4341 VCC.n3929 4.5005
R39750 VCC.n4346 VCC.n4345 4.5005
R39751 VCC.n4330 VCC.n4329 4.5005
R39752 VCC.n4335 VCC.n4334 4.5005
R39753 VCC.n3898 VCC.n3897 4.5005
R39754 VCC.n4409 VCC.n3898 4.5005
R39755 VCC.n4397 VCC.n4396 4.5005
R39756 VCC.n3908 VCC.n3895 4.5005
R39757 VCC.n4387 VCC.n4386 4.5005
R39758 VCC.n3917 VCC.n3915 4.5005
R39759 VCC.n4388 VCC.n3910 4.5005
R39760 VCC.n4398 VCC.n3906 4.5005
R39761 VCC.n4400 VCC.n4399 4.5005
R39762 VCC.n4400 VCC.n3904 4.5005
R39763 VCC.n4421 VCC.n3890 4.5005
R39764 VCC.n4432 VCC.n4431 4.5005
R39765 VCC.n3932 VCC.n3930 4.5005
R39766 VCC.n4891 VCC.n4493 4.5005
R39767 VCC.n4894 VCC.n4893 4.5005
R39768 VCC.n4968 VCC.n4448 4.5005
R39769 VCC.n4970 VCC.n4969 4.5005
R39770 VCC.n4465 VCC.n4464 4.5005
R39771 VCC.n4485 VCC.n4483 4.5005
R39772 VCC.n4495 VCC.n4482 4.5005
R39773 VCC.n4924 VCC.n4923 4.5005
R39774 VCC.n4933 VCC.n4932 4.5005
R39775 VCC.n4476 VCC.n4475 4.5005
R39776 VCC.n4456 VCC.n4455 4.5005
R39777 VCC.n4959 VCC.n4958 4.5005
R39778 VCC.n4971 VCC.n4446 4.5005
R39779 VCC.n4460 VCC.n4458 4.5005
R39780 VCC.n4931 VCC.n4930 4.5005
R39781 VCC.n4892 VCC.n4890 4.5005
R39782 VCC.n4888 VCC.n4887 4.5005
R39783 VCC.n4903 VCC.n4494 4.5005
R39784 VCC.n4973 VCC.n4972 4.5005
R39785 VCC.n4973 VCC.n4444 4.5005
R39786 VCC.n4463 VCC.n4461 4.5005
R39787 VCC.n4468 VCC.n4461 4.5005
R39788 VCC.n4919 VCC.n4918 4.5005
R39789 VCC.n4920 VCC.n4919 4.5005
R39790 VCC.n4986 VCC.n4985 4.5005
R39791 VCC.n4873 VCC.n4510 4.5005
R39792 VCC.n4872 VCC.n4871 4.5005
R39793 VCC.n4837 VCC.n4522 4.5005
R39794 VCC.n4791 VCC.n4790 4.5005
R39795 VCC.n4765 VCC.n4764 4.5005
R39796 VCC.n4760 VCC.n4756 4.5005
R39797 VCC.n4766 VCC.n4562 4.5005
R39798 VCC.n4562 VCC.n4560 4.5005
R39799 VCC.n4884 VCC.n4883 4.5005
R39800 VCC.n4839 VCC.n4838 4.5005
R39801 VCC.n4759 VCC.n4758 4.5005
R39802 VCC.n4553 VCC.n4549 4.5005
R39803 VCC.n4776 VCC.n4553 4.5005
R39804 VCC.n4789 VCC.n4788 4.5005
R39805 VCC.n4804 VCC.n4803 4.5005
R39806 VCC.n4803 VCC.n4802 4.5005
R39807 VCC.n4819 VCC.n4818 4.5005
R39808 VCC.n4820 VCC.n4819 4.5005
R39809 VCC.n4811 VCC.n4532 4.5005
R39810 VCC.n4822 VCC.n4532 4.5005
R39811 VCC.n4826 VCC.n4524 4.5005
R39812 VCC.n4827 VCC.n4826 4.5005
R39813 VCC.n4847 VCC.n4846 4.5005
R39814 VCC.n4848 VCC.n4847 4.5005
R39815 VCC.n4875 VCC.n4874 4.5005
R39816 VCC.n4513 VCC.n4511 4.5005
R39817 VCC.n4868 VCC.n4513 4.5005
R39818 VCC.n4738 VCC.n4572 4.5005
R39819 VCC.n4737 VCC.n4736 4.5005
R39820 VCC.n4711 VCC.n4583 4.5005
R39821 VCC.n4676 VCC.n4675 4.5005
R39822 VCC.n4641 VCC.n4640 4.5005
R39823 VCC.n4637 VCC.n4634 4.5005
R39824 VCC.n4643 VCC.n4642 4.5005
R39825 VCC.n4644 VCC.n4643 4.5005
R39826 VCC.n4749 VCC.n4748 4.5005
R39827 VCC.n4713 VCC.n4712 4.5005
R39828 VCC.n4636 VCC.n4635 4.5005
R39829 VCC.n4658 VCC.n4611 4.5005
R39830 VCC.n4658 VCC.n4621 4.5005
R39831 VCC.n4673 VCC.n4612 4.5005
R39832 VCC.n4683 VCC.n4682 4.5005
R39833 VCC.n4684 VCC.n4683 4.5005
R39834 VCC.n4688 VCC.n4603 4.5005
R39835 VCC.n4688 VCC.n4592 4.5005
R39836 VCC.n4691 VCC.n4604 4.5005
R39837 VCC.n4699 VCC.n4698 4.5005
R39838 VCC.n4700 VCC.n4699 4.5005
R39839 VCC.n4595 VCC.n4585 4.5005
R39840 VCC.n4596 VCC.n4595 4.5005
R39841 VCC.n4721 VCC.n4720 4.5005
R39842 VCC.n4722 VCC.n4721 4.5005
R39843 VCC.n4740 VCC.n4739 4.5005
R39844 VCC.n4575 VCC.n4573 4.5005
R39845 VCC.n4733 VCC.n4575 4.5005
R39846 VCC.n5289 VCC.n5123 4.5005
R39847 VCC.n5288 VCC.n5287 4.5005
R39848 VCC.n5192 VCC.n5191 4.5005
R39849 VCC.n5188 VCC.n5185 4.5005
R39850 VCC.n5224 VCC.n5163 4.5005
R39851 VCC.n5234 VCC.n5233 4.5005
R39852 VCC.n5235 VCC.n5234 4.5005
R39853 VCC.n5187 VCC.n5186 4.5005
R39854 VCC.n5209 VCC.n5162 4.5005
R39855 VCC.n5209 VCC.n5172 4.5005
R39856 VCC.n5194 VCC.n5193 4.5005
R39857 VCC.n5195 VCC.n5194 4.5005
R39858 VCC.n5239 VCC.n5154 4.5005
R39859 VCC.n5239 VCC.n5143 4.5005
R39860 VCC.n5300 VCC.n5299 4.5005
R39861 VCC.n5264 VCC.n5263 4.5005
R39862 VCC.n5262 VCC.n5134 4.5005
R39863 VCC.n5242 VCC.n5155 4.5005
R39864 VCC.n5250 VCC.n5249 4.5005
R39865 VCC.n5251 VCC.n5250 4.5005
R39866 VCC.n5146 VCC.n5136 4.5005
R39867 VCC.n5147 VCC.n5146 4.5005
R39868 VCC.n5272 VCC.n5271 4.5005
R39869 VCC.n5273 VCC.n5272 4.5005
R39870 VCC.n5291 VCC.n5290 4.5005
R39871 VCC.n5126 VCC.n5124 4.5005
R39872 VCC.n5284 VCC.n5126 4.5005
R39873 VCC.n5227 VCC.n5226 4.5005
R39874 VCC.n5424 VCC.n5062 4.5005
R39875 VCC.n5423 VCC.n5422 4.5005
R39876 VCC.n5317 VCC.n5316 4.5005
R39877 VCC.n5312 VCC.n5309 4.5005
R39878 VCC.n5341 VCC.n5340 4.5005
R39879 VCC.n5311 VCC.n5310 4.5005
R39880 VCC.n5435 VCC.n5434 4.5005
R39881 VCC.n5391 VCC.n5390 4.5005
R39882 VCC.n5389 VCC.n5074 4.5005
R39883 VCC.n5426 VCC.n5425 4.5005
R39884 VCC.n5343 VCC.n5342 4.5005
R39885 VCC.n5356 VCC.n5355 4.5005
R39886 VCC.n5355 VCC.n5354 4.5005
R39887 VCC.n5105 VCC.n5101 4.5005
R39888 VCC.n5328 VCC.n5105 4.5005
R39889 VCC.n5319 VCC.n5318 4.5005
R39890 VCC.n5319 VCC.n5112 4.5005
R39891 VCC.n5371 VCC.n5370 4.5005
R39892 VCC.n5372 VCC.n5371 4.5005
R39893 VCC.n5363 VCC.n5084 4.5005
R39894 VCC.n5374 VCC.n5084 4.5005
R39895 VCC.n5378 VCC.n5076 4.5005
R39896 VCC.n5379 VCC.n5378 4.5005
R39897 VCC.n5399 VCC.n5398 4.5005
R39898 VCC.n5400 VCC.n5399 4.5005
R39899 VCC.n5065 VCC.n5063 4.5005
R39900 VCC.n5419 VCC.n5065 4.5005
R39901 VCC.n5005 VCC.n5000 4.5005
R39902 VCC.n5532 VCC.n5531 4.5005
R39903 VCC.n5442 VCC.n5441 4.5005
R39904 VCC.n5048 VCC.n5046 4.5005
R39905 VCC.n5467 VCC.n5466 4.5005
R39906 VCC.n5034 VCC.n5032 4.5005
R39907 VCC.n5032 VCC.n5031 4.5005
R39908 VCC.n5036 VCC.n5035 4.5005
R39909 VCC.n5450 VCC.n5038 4.5005
R39910 VCC.n5455 VCC.n5454 4.5005
R39911 VCC.n5439 VCC.n5438 4.5005
R39912 VCC.n5444 VCC.n5443 4.5005
R39913 VCC.n5007 VCC.n5006 4.5005
R39914 VCC.n5518 VCC.n5007 4.5005
R39915 VCC.n5506 VCC.n5505 4.5005
R39916 VCC.n5017 VCC.n5004 4.5005
R39917 VCC.n5496 VCC.n5495 4.5005
R39918 VCC.n5026 VCC.n5024 4.5005
R39919 VCC.n5497 VCC.n5019 4.5005
R39920 VCC.n5507 VCC.n5015 4.5005
R39921 VCC.n5509 VCC.n5508 4.5005
R39922 VCC.n5509 VCC.n5013 4.5005
R39923 VCC.n5530 VCC.n4999 4.5005
R39924 VCC.n5541 VCC.n5540 4.5005
R39925 VCC.n5041 VCC.n5039 4.5005
R39926 VCC.n6000 VCC.n5602 4.5005
R39927 VCC.n6003 VCC.n6002 4.5005
R39928 VCC.n6077 VCC.n5557 4.5005
R39929 VCC.n6079 VCC.n6078 4.5005
R39930 VCC.n5574 VCC.n5573 4.5005
R39931 VCC.n5594 VCC.n5592 4.5005
R39932 VCC.n5604 VCC.n5591 4.5005
R39933 VCC.n6033 VCC.n6032 4.5005
R39934 VCC.n6042 VCC.n6041 4.5005
R39935 VCC.n5585 VCC.n5584 4.5005
R39936 VCC.n5565 VCC.n5564 4.5005
R39937 VCC.n6068 VCC.n6067 4.5005
R39938 VCC.n6080 VCC.n5555 4.5005
R39939 VCC.n5569 VCC.n5567 4.5005
R39940 VCC.n6040 VCC.n6039 4.5005
R39941 VCC.n6001 VCC.n5999 4.5005
R39942 VCC.n5997 VCC.n5996 4.5005
R39943 VCC.n6012 VCC.n5603 4.5005
R39944 VCC.n6082 VCC.n6081 4.5005
R39945 VCC.n6082 VCC.n5553 4.5005
R39946 VCC.n5572 VCC.n5570 4.5005
R39947 VCC.n5577 VCC.n5570 4.5005
R39948 VCC.n6028 VCC.n6027 4.5005
R39949 VCC.n6029 VCC.n6028 4.5005
R39950 VCC.n6095 VCC.n6094 4.5005
R39951 VCC.n5982 VCC.n5619 4.5005
R39952 VCC.n5981 VCC.n5980 4.5005
R39953 VCC.n5946 VCC.n5631 4.5005
R39954 VCC.n5900 VCC.n5899 4.5005
R39955 VCC.n5874 VCC.n5873 4.5005
R39956 VCC.n5869 VCC.n5865 4.5005
R39957 VCC.n5875 VCC.n5671 4.5005
R39958 VCC.n5671 VCC.n5669 4.5005
R39959 VCC.n5993 VCC.n5992 4.5005
R39960 VCC.n5948 VCC.n5947 4.5005
R39961 VCC.n5868 VCC.n5867 4.5005
R39962 VCC.n5662 VCC.n5658 4.5005
R39963 VCC.n5885 VCC.n5662 4.5005
R39964 VCC.n5898 VCC.n5897 4.5005
R39965 VCC.n5913 VCC.n5912 4.5005
R39966 VCC.n5912 VCC.n5911 4.5005
R39967 VCC.n5928 VCC.n5927 4.5005
R39968 VCC.n5929 VCC.n5928 4.5005
R39969 VCC.n5920 VCC.n5641 4.5005
R39970 VCC.n5931 VCC.n5641 4.5005
R39971 VCC.n5935 VCC.n5633 4.5005
R39972 VCC.n5936 VCC.n5935 4.5005
R39973 VCC.n5956 VCC.n5955 4.5005
R39974 VCC.n5957 VCC.n5956 4.5005
R39975 VCC.n5984 VCC.n5983 4.5005
R39976 VCC.n5622 VCC.n5620 4.5005
R39977 VCC.n5977 VCC.n5622 4.5005
R39978 VCC.n5847 VCC.n5681 4.5005
R39979 VCC.n5846 VCC.n5845 4.5005
R39980 VCC.n5820 VCC.n5692 4.5005
R39981 VCC.n5785 VCC.n5784 4.5005
R39982 VCC.n5750 VCC.n5749 4.5005
R39983 VCC.n5746 VCC.n5743 4.5005
R39984 VCC.n5752 VCC.n5751 4.5005
R39985 VCC.n5753 VCC.n5752 4.5005
R39986 VCC.n5858 VCC.n5857 4.5005
R39987 VCC.n5822 VCC.n5821 4.5005
R39988 VCC.n5745 VCC.n5744 4.5005
R39989 VCC.n5767 VCC.n5720 4.5005
R39990 VCC.n5767 VCC.n5730 4.5005
R39991 VCC.n5782 VCC.n5721 4.5005
R39992 VCC.n5792 VCC.n5791 4.5005
R39993 VCC.n5793 VCC.n5792 4.5005
R39994 VCC.n5797 VCC.n5712 4.5005
R39995 VCC.n5797 VCC.n5701 4.5005
R39996 VCC.n5800 VCC.n5713 4.5005
R39997 VCC.n5808 VCC.n5807 4.5005
R39998 VCC.n5809 VCC.n5808 4.5005
R39999 VCC.n5704 VCC.n5694 4.5005
R40000 VCC.n5705 VCC.n5704 4.5005
R40001 VCC.n5830 VCC.n5829 4.5005
R40002 VCC.n5831 VCC.n5830 4.5005
R40003 VCC.n5849 VCC.n5848 4.5005
R40004 VCC.n5684 VCC.n5682 4.5005
R40005 VCC.n5842 VCC.n5684 4.5005
R40006 VCC.n6398 VCC.n6232 4.5005
R40007 VCC.n6397 VCC.n6396 4.5005
R40008 VCC.n6301 VCC.n6300 4.5005
R40009 VCC.n6297 VCC.n6294 4.5005
R40010 VCC.n6333 VCC.n6272 4.5005
R40011 VCC.n6343 VCC.n6342 4.5005
R40012 VCC.n6344 VCC.n6343 4.5005
R40013 VCC.n6296 VCC.n6295 4.5005
R40014 VCC.n6318 VCC.n6271 4.5005
R40015 VCC.n6318 VCC.n6281 4.5005
R40016 VCC.n6303 VCC.n6302 4.5005
R40017 VCC.n6304 VCC.n6303 4.5005
R40018 VCC.n6348 VCC.n6263 4.5005
R40019 VCC.n6348 VCC.n6252 4.5005
R40020 VCC.n6409 VCC.n6408 4.5005
R40021 VCC.n6373 VCC.n6372 4.5005
R40022 VCC.n6371 VCC.n6243 4.5005
R40023 VCC.n6351 VCC.n6264 4.5005
R40024 VCC.n6359 VCC.n6358 4.5005
R40025 VCC.n6360 VCC.n6359 4.5005
R40026 VCC.n6255 VCC.n6245 4.5005
R40027 VCC.n6256 VCC.n6255 4.5005
R40028 VCC.n6381 VCC.n6380 4.5005
R40029 VCC.n6382 VCC.n6381 4.5005
R40030 VCC.n6400 VCC.n6399 4.5005
R40031 VCC.n6235 VCC.n6233 4.5005
R40032 VCC.n6393 VCC.n6235 4.5005
R40033 VCC.n6336 VCC.n6335 4.5005
R40034 VCC.n6533 VCC.n6171 4.5005
R40035 VCC.n6532 VCC.n6531 4.5005
R40036 VCC.n6426 VCC.n6425 4.5005
R40037 VCC.n6421 VCC.n6418 4.5005
R40038 VCC.n6450 VCC.n6449 4.5005
R40039 VCC.n6420 VCC.n6419 4.5005
R40040 VCC.n6544 VCC.n6543 4.5005
R40041 VCC.n6500 VCC.n6499 4.5005
R40042 VCC.n6498 VCC.n6183 4.5005
R40043 VCC.n6535 VCC.n6534 4.5005
R40044 VCC.n6452 VCC.n6451 4.5005
R40045 VCC.n6465 VCC.n6464 4.5005
R40046 VCC.n6464 VCC.n6463 4.5005
R40047 VCC.n6214 VCC.n6210 4.5005
R40048 VCC.n6437 VCC.n6214 4.5005
R40049 VCC.n6428 VCC.n6427 4.5005
R40050 VCC.n6428 VCC.n6221 4.5005
R40051 VCC.n6480 VCC.n6479 4.5005
R40052 VCC.n6481 VCC.n6480 4.5005
R40053 VCC.n6472 VCC.n6193 4.5005
R40054 VCC.n6483 VCC.n6193 4.5005
R40055 VCC.n6487 VCC.n6185 4.5005
R40056 VCC.n6488 VCC.n6487 4.5005
R40057 VCC.n6508 VCC.n6507 4.5005
R40058 VCC.n6509 VCC.n6508 4.5005
R40059 VCC.n6174 VCC.n6172 4.5005
R40060 VCC.n6528 VCC.n6174 4.5005
R40061 VCC.n6114 VCC.n6109 4.5005
R40062 VCC.n6641 VCC.n6640 4.5005
R40063 VCC.n6551 VCC.n6550 4.5005
R40064 VCC.n6157 VCC.n6155 4.5005
R40065 VCC.n6576 VCC.n6575 4.5005
R40066 VCC.n6143 VCC.n6141 4.5005
R40067 VCC.n6141 VCC.n6140 4.5005
R40068 VCC.n6145 VCC.n6144 4.5005
R40069 VCC.n6559 VCC.n6147 4.5005
R40070 VCC.n6564 VCC.n6563 4.5005
R40071 VCC.n6548 VCC.n6547 4.5005
R40072 VCC.n6553 VCC.n6552 4.5005
R40073 VCC.n6116 VCC.n6115 4.5005
R40074 VCC.n6627 VCC.n6116 4.5005
R40075 VCC.n6615 VCC.n6614 4.5005
R40076 VCC.n6126 VCC.n6113 4.5005
R40077 VCC.n6605 VCC.n6604 4.5005
R40078 VCC.n6135 VCC.n6133 4.5005
R40079 VCC.n6606 VCC.n6128 4.5005
R40080 VCC.n6616 VCC.n6124 4.5005
R40081 VCC.n6618 VCC.n6617 4.5005
R40082 VCC.n6618 VCC.n6122 4.5005
R40083 VCC.n6639 VCC.n6108 4.5005
R40084 VCC.n6650 VCC.n6649 4.5005
R40085 VCC.n6150 VCC.n6148 4.5005
R40086 VCC.n7109 VCC.n6711 4.5005
R40087 VCC.n7112 VCC.n7111 4.5005
R40088 VCC.n7186 VCC.n6666 4.5005
R40089 VCC.n7188 VCC.n7187 4.5005
R40090 VCC.n6683 VCC.n6682 4.5005
R40091 VCC.n6703 VCC.n6701 4.5005
R40092 VCC.n6713 VCC.n6700 4.5005
R40093 VCC.n7142 VCC.n7141 4.5005
R40094 VCC.n7151 VCC.n7150 4.5005
R40095 VCC.n6694 VCC.n6693 4.5005
R40096 VCC.n6674 VCC.n6673 4.5005
R40097 VCC.n7177 VCC.n7176 4.5005
R40098 VCC.n7189 VCC.n6664 4.5005
R40099 VCC.n6678 VCC.n6676 4.5005
R40100 VCC.n7149 VCC.n7148 4.5005
R40101 VCC.n7110 VCC.n7108 4.5005
R40102 VCC.n7106 VCC.n7105 4.5005
R40103 VCC.n7121 VCC.n6712 4.5005
R40104 VCC.n7191 VCC.n7190 4.5005
R40105 VCC.n7191 VCC.n6662 4.5005
R40106 VCC.n6681 VCC.n6679 4.5005
R40107 VCC.n6686 VCC.n6679 4.5005
R40108 VCC.n7137 VCC.n7136 4.5005
R40109 VCC.n7138 VCC.n7137 4.5005
R40110 VCC.n7204 VCC.n7203 4.5005
R40111 VCC.n7091 VCC.n6728 4.5005
R40112 VCC.n7090 VCC.n7089 4.5005
R40113 VCC.n7055 VCC.n6740 4.5005
R40114 VCC.n7009 VCC.n7008 4.5005
R40115 VCC.n6983 VCC.n6982 4.5005
R40116 VCC.n6978 VCC.n6974 4.5005
R40117 VCC.n6984 VCC.n6780 4.5005
R40118 VCC.n6780 VCC.n6778 4.5005
R40119 VCC.n7102 VCC.n7101 4.5005
R40120 VCC.n7057 VCC.n7056 4.5005
R40121 VCC.n6977 VCC.n6976 4.5005
R40122 VCC.n6771 VCC.n6767 4.5005
R40123 VCC.n6994 VCC.n6771 4.5005
R40124 VCC.n7007 VCC.n7006 4.5005
R40125 VCC.n7022 VCC.n7021 4.5005
R40126 VCC.n7021 VCC.n7020 4.5005
R40127 VCC.n7037 VCC.n7036 4.5005
R40128 VCC.n7038 VCC.n7037 4.5005
R40129 VCC.n7029 VCC.n6750 4.5005
R40130 VCC.n7040 VCC.n6750 4.5005
R40131 VCC.n7044 VCC.n6742 4.5005
R40132 VCC.n7045 VCC.n7044 4.5005
R40133 VCC.n7065 VCC.n7064 4.5005
R40134 VCC.n7066 VCC.n7065 4.5005
R40135 VCC.n7093 VCC.n7092 4.5005
R40136 VCC.n6731 VCC.n6729 4.5005
R40137 VCC.n7086 VCC.n6731 4.5005
R40138 VCC.n6956 VCC.n6790 4.5005
R40139 VCC.n6955 VCC.n6954 4.5005
R40140 VCC.n6929 VCC.n6801 4.5005
R40141 VCC.n6894 VCC.n6893 4.5005
R40142 VCC.n6859 VCC.n6858 4.5005
R40143 VCC.n6855 VCC.n6852 4.5005
R40144 VCC.n6861 VCC.n6860 4.5005
R40145 VCC.n6862 VCC.n6861 4.5005
R40146 VCC.n6967 VCC.n6966 4.5005
R40147 VCC.n6931 VCC.n6930 4.5005
R40148 VCC.n6854 VCC.n6853 4.5005
R40149 VCC.n6876 VCC.n6829 4.5005
R40150 VCC.n6876 VCC.n6839 4.5005
R40151 VCC.n6891 VCC.n6830 4.5005
R40152 VCC.n6901 VCC.n6900 4.5005
R40153 VCC.n6902 VCC.n6901 4.5005
R40154 VCC.n6906 VCC.n6821 4.5005
R40155 VCC.n6906 VCC.n6810 4.5005
R40156 VCC.n6909 VCC.n6822 4.5005
R40157 VCC.n6917 VCC.n6916 4.5005
R40158 VCC.n6918 VCC.n6917 4.5005
R40159 VCC.n6813 VCC.n6803 4.5005
R40160 VCC.n6814 VCC.n6813 4.5005
R40161 VCC.n6939 VCC.n6938 4.5005
R40162 VCC.n6940 VCC.n6939 4.5005
R40163 VCC.n6958 VCC.n6957 4.5005
R40164 VCC.n6793 VCC.n6791 4.5005
R40165 VCC.n6951 VCC.n6793 4.5005
R40166 VCC.n7507 VCC.n7341 4.5005
R40167 VCC.n7506 VCC.n7505 4.5005
R40168 VCC.n7410 VCC.n7409 4.5005
R40169 VCC.n7406 VCC.n7403 4.5005
R40170 VCC.n7442 VCC.n7381 4.5005
R40171 VCC.n7452 VCC.n7451 4.5005
R40172 VCC.n7453 VCC.n7452 4.5005
R40173 VCC.n7405 VCC.n7404 4.5005
R40174 VCC.n7427 VCC.n7380 4.5005
R40175 VCC.n7427 VCC.n7390 4.5005
R40176 VCC.n7412 VCC.n7411 4.5005
R40177 VCC.n7413 VCC.n7412 4.5005
R40178 VCC.n7457 VCC.n7372 4.5005
R40179 VCC.n7457 VCC.n7361 4.5005
R40180 VCC.n7518 VCC.n7517 4.5005
R40181 VCC.n7482 VCC.n7481 4.5005
R40182 VCC.n7480 VCC.n7352 4.5005
R40183 VCC.n7460 VCC.n7373 4.5005
R40184 VCC.n7468 VCC.n7467 4.5005
R40185 VCC.n7469 VCC.n7468 4.5005
R40186 VCC.n7364 VCC.n7354 4.5005
R40187 VCC.n7365 VCC.n7364 4.5005
R40188 VCC.n7490 VCC.n7489 4.5005
R40189 VCC.n7491 VCC.n7490 4.5005
R40190 VCC.n7509 VCC.n7508 4.5005
R40191 VCC.n7344 VCC.n7342 4.5005
R40192 VCC.n7502 VCC.n7344 4.5005
R40193 VCC.n7445 VCC.n7444 4.5005
R40194 VCC.n7642 VCC.n7280 4.5005
R40195 VCC.n7641 VCC.n7640 4.5005
R40196 VCC.n7535 VCC.n7534 4.5005
R40197 VCC.n7530 VCC.n7527 4.5005
R40198 VCC.n7559 VCC.n7558 4.5005
R40199 VCC.n7529 VCC.n7528 4.5005
R40200 VCC.n7653 VCC.n7652 4.5005
R40201 VCC.n7609 VCC.n7608 4.5005
R40202 VCC.n7607 VCC.n7292 4.5005
R40203 VCC.n7644 VCC.n7643 4.5005
R40204 VCC.n7561 VCC.n7560 4.5005
R40205 VCC.n7574 VCC.n7573 4.5005
R40206 VCC.n7573 VCC.n7572 4.5005
R40207 VCC.n7323 VCC.n7319 4.5005
R40208 VCC.n7546 VCC.n7323 4.5005
R40209 VCC.n7537 VCC.n7536 4.5005
R40210 VCC.n7537 VCC.n7330 4.5005
R40211 VCC.n7589 VCC.n7588 4.5005
R40212 VCC.n7590 VCC.n7589 4.5005
R40213 VCC.n7581 VCC.n7302 4.5005
R40214 VCC.n7592 VCC.n7302 4.5005
R40215 VCC.n7596 VCC.n7294 4.5005
R40216 VCC.n7597 VCC.n7596 4.5005
R40217 VCC.n7617 VCC.n7616 4.5005
R40218 VCC.n7618 VCC.n7617 4.5005
R40219 VCC.n7283 VCC.n7281 4.5005
R40220 VCC.n7637 VCC.n7283 4.5005
R40221 VCC.n7223 VCC.n7218 4.5005
R40222 VCC.n7750 VCC.n7749 4.5005
R40223 VCC.n7660 VCC.n7659 4.5005
R40224 VCC.n7266 VCC.n7264 4.5005
R40225 VCC.n7685 VCC.n7684 4.5005
R40226 VCC.n7252 VCC.n7250 4.5005
R40227 VCC.n7250 VCC.n7249 4.5005
R40228 VCC.n7254 VCC.n7253 4.5005
R40229 VCC.n7668 VCC.n7256 4.5005
R40230 VCC.n7673 VCC.n7672 4.5005
R40231 VCC.n7657 VCC.n7656 4.5005
R40232 VCC.n7662 VCC.n7661 4.5005
R40233 VCC.n7225 VCC.n7224 4.5005
R40234 VCC.n7736 VCC.n7225 4.5005
R40235 VCC.n7724 VCC.n7723 4.5005
R40236 VCC.n7235 VCC.n7222 4.5005
R40237 VCC.n7714 VCC.n7713 4.5005
R40238 VCC.n7244 VCC.n7242 4.5005
R40239 VCC.n7715 VCC.n7237 4.5005
R40240 VCC.n7725 VCC.n7233 4.5005
R40241 VCC.n7727 VCC.n7726 4.5005
R40242 VCC.n7727 VCC.n7231 4.5005
R40243 VCC.n7748 VCC.n7217 4.5005
R40244 VCC.n7759 VCC.n7758 4.5005
R40245 VCC.n7259 VCC.n7257 4.5005
R40246 VCC.n8218 VCC.n7820 4.5005
R40247 VCC.n8221 VCC.n8220 4.5005
R40248 VCC.n8295 VCC.n7775 4.5005
R40249 VCC.n8297 VCC.n8296 4.5005
R40250 VCC.n7792 VCC.n7791 4.5005
R40251 VCC.n7812 VCC.n7810 4.5005
R40252 VCC.n7822 VCC.n7809 4.5005
R40253 VCC.n8251 VCC.n8250 4.5005
R40254 VCC.n8260 VCC.n8259 4.5005
R40255 VCC.n7803 VCC.n7802 4.5005
R40256 VCC.n7783 VCC.n7782 4.5005
R40257 VCC.n8286 VCC.n8285 4.5005
R40258 VCC.n8298 VCC.n7773 4.5005
R40259 VCC.n7787 VCC.n7785 4.5005
R40260 VCC.n8258 VCC.n8257 4.5005
R40261 VCC.n8219 VCC.n8217 4.5005
R40262 VCC.n8215 VCC.n8214 4.5005
R40263 VCC.n8230 VCC.n7821 4.5005
R40264 VCC.n8300 VCC.n8299 4.5005
R40265 VCC.n8300 VCC.n7771 4.5005
R40266 VCC.n7790 VCC.n7788 4.5005
R40267 VCC.n7795 VCC.n7788 4.5005
R40268 VCC.n8246 VCC.n8245 4.5005
R40269 VCC.n8247 VCC.n8246 4.5005
R40270 VCC.n8313 VCC.n8312 4.5005
R40271 VCC.n8200 VCC.n7837 4.5005
R40272 VCC.n8199 VCC.n8198 4.5005
R40273 VCC.n8164 VCC.n7849 4.5005
R40274 VCC.n8118 VCC.n8117 4.5005
R40275 VCC.n8092 VCC.n8091 4.5005
R40276 VCC.n8087 VCC.n8083 4.5005
R40277 VCC.n8093 VCC.n7889 4.5005
R40278 VCC.n7889 VCC.n7887 4.5005
R40279 VCC.n8211 VCC.n8210 4.5005
R40280 VCC.n8166 VCC.n8165 4.5005
R40281 VCC.n8086 VCC.n8085 4.5005
R40282 VCC.n7880 VCC.n7876 4.5005
R40283 VCC.n8103 VCC.n7880 4.5005
R40284 VCC.n8116 VCC.n8115 4.5005
R40285 VCC.n8131 VCC.n8130 4.5005
R40286 VCC.n8130 VCC.n8129 4.5005
R40287 VCC.n8146 VCC.n8145 4.5005
R40288 VCC.n8147 VCC.n8146 4.5005
R40289 VCC.n8138 VCC.n7859 4.5005
R40290 VCC.n8149 VCC.n7859 4.5005
R40291 VCC.n8153 VCC.n7851 4.5005
R40292 VCC.n8154 VCC.n8153 4.5005
R40293 VCC.n8174 VCC.n8173 4.5005
R40294 VCC.n8175 VCC.n8174 4.5005
R40295 VCC.n8202 VCC.n8201 4.5005
R40296 VCC.n7840 VCC.n7838 4.5005
R40297 VCC.n8195 VCC.n7840 4.5005
R40298 VCC.n8065 VCC.n7899 4.5005
R40299 VCC.n8064 VCC.n8063 4.5005
R40300 VCC.n8038 VCC.n7910 4.5005
R40301 VCC.n8003 VCC.n8002 4.5005
R40302 VCC.n7968 VCC.n7967 4.5005
R40303 VCC.n7964 VCC.n7961 4.5005
R40304 VCC.n7970 VCC.n7969 4.5005
R40305 VCC.n7971 VCC.n7970 4.5005
R40306 VCC.n8076 VCC.n8075 4.5005
R40307 VCC.n8040 VCC.n8039 4.5005
R40308 VCC.n7963 VCC.n7962 4.5005
R40309 VCC.n7985 VCC.n7938 4.5005
R40310 VCC.n7985 VCC.n7948 4.5005
R40311 VCC.n8000 VCC.n7939 4.5005
R40312 VCC.n8010 VCC.n8009 4.5005
R40313 VCC.n8011 VCC.n8010 4.5005
R40314 VCC.n8015 VCC.n7930 4.5005
R40315 VCC.n8015 VCC.n7919 4.5005
R40316 VCC.n8018 VCC.n7931 4.5005
R40317 VCC.n8026 VCC.n8025 4.5005
R40318 VCC.n8027 VCC.n8026 4.5005
R40319 VCC.n7922 VCC.n7912 4.5005
R40320 VCC.n7923 VCC.n7922 4.5005
R40321 VCC.n8048 VCC.n8047 4.5005
R40322 VCC.n8049 VCC.n8048 4.5005
R40323 VCC.n8067 VCC.n8066 4.5005
R40324 VCC.n7902 VCC.n7900 4.5005
R40325 VCC.n8060 VCC.n7902 4.5005
R40326 VCC.n8751 VCC.n8389 4.5005
R40327 VCC.n8750 VCC.n8749 4.5005
R40328 VCC.n8644 VCC.n8643 4.5005
R40329 VCC.n8639 VCC.n8636 4.5005
R40330 VCC.n8668 VCC.n8667 4.5005
R40331 VCC.n8638 VCC.n8637 4.5005
R40332 VCC.n8762 VCC.n8761 4.5005
R40333 VCC.n8718 VCC.n8717 4.5005
R40334 VCC.n8716 VCC.n8401 4.5005
R40335 VCC.n8753 VCC.n8752 4.5005
R40336 VCC.n8670 VCC.n8669 4.5005
R40337 VCC.n8683 VCC.n8682 4.5005
R40338 VCC.n8682 VCC.n8681 4.5005
R40339 VCC.n8432 VCC.n8428 4.5005
R40340 VCC.n8655 VCC.n8432 4.5005
R40341 VCC.n8646 VCC.n8645 4.5005
R40342 VCC.n8646 VCC.n8439 4.5005
R40343 VCC.n8698 VCC.n8697 4.5005
R40344 VCC.n8699 VCC.n8698 4.5005
R40345 VCC.n8690 VCC.n8411 4.5005
R40346 VCC.n8701 VCC.n8411 4.5005
R40347 VCC.n8705 VCC.n8403 4.5005
R40348 VCC.n8706 VCC.n8705 4.5005
R40349 VCC.n8726 VCC.n8725 4.5005
R40350 VCC.n8727 VCC.n8726 4.5005
R40351 VCC.n8392 VCC.n8390 4.5005
R40352 VCC.n8746 VCC.n8392 4.5005
R40353 VCC.n8332 VCC.n8327 4.5005
R40354 VCC.n8859 VCC.n8858 4.5005
R40355 VCC.n8769 VCC.n8768 4.5005
R40356 VCC.n8375 VCC.n8373 4.5005
R40357 VCC.n8794 VCC.n8793 4.5005
R40358 VCC.n8361 VCC.n8359 4.5005
R40359 VCC.n8359 VCC.n8358 4.5005
R40360 VCC.n8363 VCC.n8362 4.5005
R40361 VCC.n8777 VCC.n8365 4.5005
R40362 VCC.n8782 VCC.n8781 4.5005
R40363 VCC.n8766 VCC.n8765 4.5005
R40364 VCC.n8771 VCC.n8770 4.5005
R40365 VCC.n8334 VCC.n8333 4.5005
R40366 VCC.n8845 VCC.n8334 4.5005
R40367 VCC.n8833 VCC.n8832 4.5005
R40368 VCC.n8344 VCC.n8331 4.5005
R40369 VCC.n8823 VCC.n8822 4.5005
R40370 VCC.n8353 VCC.n8351 4.5005
R40371 VCC.n8824 VCC.n8346 4.5005
R40372 VCC.n8834 VCC.n8342 4.5005
R40373 VCC.n8836 VCC.n8835 4.5005
R40374 VCC.n8836 VCC.n8340 4.5005
R40375 VCC.n8857 VCC.n8326 4.5005
R40376 VCC.n8868 VCC.n8867 4.5005
R40377 VCC.n8368 VCC.n8366 4.5005
R40378 VCC.n8616 VCC.n8450 4.5005
R40379 VCC.n8615 VCC.n8614 4.5005
R40380 VCC.n8589 VCC.n8461 4.5005
R40381 VCC.n8554 VCC.n8553 4.5005
R40382 VCC.n8519 VCC.n8518 4.5005
R40383 VCC.n8515 VCC.n8512 4.5005
R40384 VCC.n8521 VCC.n8520 4.5005
R40385 VCC.n8522 VCC.n8521 4.5005
R40386 VCC.n8627 VCC.n8626 4.5005
R40387 VCC.n8591 VCC.n8590 4.5005
R40388 VCC.n8514 VCC.n8513 4.5005
R40389 VCC.n8536 VCC.n8489 4.5005
R40390 VCC.n8536 VCC.n8499 4.5005
R40391 VCC.n8551 VCC.n8490 4.5005
R40392 VCC.n8561 VCC.n8560 4.5005
R40393 VCC.n8562 VCC.n8561 4.5005
R40394 VCC.n8566 VCC.n8481 4.5005
R40395 VCC.n8566 VCC.n8470 4.5005
R40396 VCC.n8569 VCC.n8482 4.5005
R40397 VCC.n8577 VCC.n8576 4.5005
R40398 VCC.n8578 VCC.n8577 4.5005
R40399 VCC.n8473 VCC.n8463 4.5005
R40400 VCC.n8474 VCC.n8473 4.5005
R40401 VCC.n8599 VCC.n8598 4.5005
R40402 VCC.n8600 VCC.n8599 4.5005
R40403 VCC.n8618 VCC.n8617 4.5005
R40404 VCC.n8453 VCC.n8451 4.5005
R40405 VCC.n8611 VCC.n8453 4.5005
R40406 VCC.n9327 VCC.n8929 4.5005
R40407 VCC.n9330 VCC.n9329 4.5005
R40408 VCC.n9404 VCC.n8884 4.5005
R40409 VCC.n9406 VCC.n9405 4.5005
R40410 VCC.n8901 VCC.n8900 4.5005
R40411 VCC.n8921 VCC.n8919 4.5005
R40412 VCC.n8931 VCC.n8918 4.5005
R40413 VCC.n9360 VCC.n9359 4.5005
R40414 VCC.n9369 VCC.n9368 4.5005
R40415 VCC.n8912 VCC.n8911 4.5005
R40416 VCC.n8892 VCC.n8891 4.5005
R40417 VCC.n9395 VCC.n9394 4.5005
R40418 VCC.n9407 VCC.n8882 4.5005
R40419 VCC.n8896 VCC.n8894 4.5005
R40420 VCC.n9367 VCC.n9366 4.5005
R40421 VCC.n9328 VCC.n9326 4.5005
R40422 VCC.n9324 VCC.n9323 4.5005
R40423 VCC.n9339 VCC.n8930 4.5005
R40424 VCC.n9409 VCC.n9408 4.5005
R40425 VCC.n9409 VCC.n8880 4.5005
R40426 VCC.n8899 VCC.n8897 4.5005
R40427 VCC.n8904 VCC.n8897 4.5005
R40428 VCC.n9355 VCC.n9354 4.5005
R40429 VCC.n9356 VCC.n9355 4.5005
R40430 VCC.n9422 VCC.n9421 4.5005
R40431 VCC.n9309 VCC.n8946 4.5005
R40432 VCC.n9308 VCC.n9307 4.5005
R40433 VCC.n9273 VCC.n8958 4.5005
R40434 VCC.n9227 VCC.n9226 4.5005
R40435 VCC.n9201 VCC.n9200 4.5005
R40436 VCC.n9196 VCC.n9192 4.5005
R40437 VCC.n9202 VCC.n8998 4.5005
R40438 VCC.n8998 VCC.n8996 4.5005
R40439 VCC.n9320 VCC.n9319 4.5005
R40440 VCC.n9275 VCC.n9274 4.5005
R40441 VCC.n9195 VCC.n9194 4.5005
R40442 VCC.n8989 VCC.n8985 4.5005
R40443 VCC.n9212 VCC.n8989 4.5005
R40444 VCC.n9225 VCC.n9224 4.5005
R40445 VCC.n9240 VCC.n9239 4.5005
R40446 VCC.n9239 VCC.n9238 4.5005
R40447 VCC.n9255 VCC.n9254 4.5005
R40448 VCC.n9256 VCC.n9255 4.5005
R40449 VCC.n9247 VCC.n8968 4.5005
R40450 VCC.n9258 VCC.n8968 4.5005
R40451 VCC.n9262 VCC.n8960 4.5005
R40452 VCC.n9263 VCC.n9262 4.5005
R40453 VCC.n9283 VCC.n9282 4.5005
R40454 VCC.n9284 VCC.n9283 4.5005
R40455 VCC.n9311 VCC.n9310 4.5005
R40456 VCC.n8949 VCC.n8947 4.5005
R40457 VCC.n9304 VCC.n8949 4.5005
R40458 VCC.n9174 VCC.n9008 4.5005
R40459 VCC.n9173 VCC.n9172 4.5005
R40460 VCC.n9147 VCC.n9019 4.5005
R40461 VCC.n9112 VCC.n9111 4.5005
R40462 VCC.n9077 VCC.n9076 4.5005
R40463 VCC.n9073 VCC.n9070 4.5005
R40464 VCC.n9079 VCC.n9078 4.5005
R40465 VCC.n9080 VCC.n9079 4.5005
R40466 VCC.n9185 VCC.n9184 4.5005
R40467 VCC.n9149 VCC.n9148 4.5005
R40468 VCC.n9072 VCC.n9071 4.5005
R40469 VCC.n9094 VCC.n9047 4.5005
R40470 VCC.n9094 VCC.n9057 4.5005
R40471 VCC.n9109 VCC.n9048 4.5005
R40472 VCC.n9119 VCC.n9118 4.5005
R40473 VCC.n9120 VCC.n9119 4.5005
R40474 VCC.n9124 VCC.n9039 4.5005
R40475 VCC.n9124 VCC.n9028 4.5005
R40476 VCC.n9127 VCC.n9040 4.5005
R40477 VCC.n9135 VCC.n9134 4.5005
R40478 VCC.n9136 VCC.n9135 4.5005
R40479 VCC.n9031 VCC.n9021 4.5005
R40480 VCC.n9032 VCC.n9031 4.5005
R40481 VCC.n9157 VCC.n9156 4.5005
R40482 VCC.n9158 VCC.n9157 4.5005
R40483 VCC.n9176 VCC.n9175 4.5005
R40484 VCC.n9011 VCC.n9009 4.5005
R40485 VCC.n9169 VCC.n9011 4.5005
R40486 VCC.n9725 VCC.n9559 4.5005
R40487 VCC.n9724 VCC.n9723 4.5005
R40488 VCC.n9628 VCC.n9627 4.5005
R40489 VCC.n9624 VCC.n9621 4.5005
R40490 VCC.n9660 VCC.n9599 4.5005
R40491 VCC.n9670 VCC.n9669 4.5005
R40492 VCC.n9671 VCC.n9670 4.5005
R40493 VCC.n9623 VCC.n9622 4.5005
R40494 VCC.n9645 VCC.n9598 4.5005
R40495 VCC.n9645 VCC.n9608 4.5005
R40496 VCC.n9630 VCC.n9629 4.5005
R40497 VCC.n9631 VCC.n9630 4.5005
R40498 VCC.n9675 VCC.n9590 4.5005
R40499 VCC.n9675 VCC.n9579 4.5005
R40500 VCC.n9736 VCC.n9735 4.5005
R40501 VCC.n9700 VCC.n9699 4.5005
R40502 VCC.n9698 VCC.n9570 4.5005
R40503 VCC.n9678 VCC.n9591 4.5005
R40504 VCC.n9686 VCC.n9685 4.5005
R40505 VCC.n9687 VCC.n9686 4.5005
R40506 VCC.n9582 VCC.n9572 4.5005
R40507 VCC.n9583 VCC.n9582 4.5005
R40508 VCC.n9708 VCC.n9707 4.5005
R40509 VCC.n9709 VCC.n9708 4.5005
R40510 VCC.n9727 VCC.n9726 4.5005
R40511 VCC.n9562 VCC.n9560 4.5005
R40512 VCC.n9720 VCC.n9562 4.5005
R40513 VCC.n9663 VCC.n9662 4.5005
R40514 VCC.n9860 VCC.n9498 4.5005
R40515 VCC.n9859 VCC.n9858 4.5005
R40516 VCC.n9753 VCC.n9752 4.5005
R40517 VCC.n9748 VCC.n9745 4.5005
R40518 VCC.n9777 VCC.n9776 4.5005
R40519 VCC.n9747 VCC.n9746 4.5005
R40520 VCC.n9871 VCC.n9870 4.5005
R40521 VCC.n9827 VCC.n9826 4.5005
R40522 VCC.n9825 VCC.n9510 4.5005
R40523 VCC.n9862 VCC.n9861 4.5005
R40524 VCC.n9779 VCC.n9778 4.5005
R40525 VCC.n9792 VCC.n9791 4.5005
R40526 VCC.n9791 VCC.n9790 4.5005
R40527 VCC.n9541 VCC.n9537 4.5005
R40528 VCC.n9764 VCC.n9541 4.5005
R40529 VCC.n9755 VCC.n9754 4.5005
R40530 VCC.n9755 VCC.n9548 4.5005
R40531 VCC.n9807 VCC.n9806 4.5005
R40532 VCC.n9808 VCC.n9807 4.5005
R40533 VCC.n9799 VCC.n9520 4.5005
R40534 VCC.n9810 VCC.n9520 4.5005
R40535 VCC.n9814 VCC.n9512 4.5005
R40536 VCC.n9815 VCC.n9814 4.5005
R40537 VCC.n9835 VCC.n9834 4.5005
R40538 VCC.n9836 VCC.n9835 4.5005
R40539 VCC.n9501 VCC.n9499 4.5005
R40540 VCC.n9855 VCC.n9501 4.5005
R40541 VCC.n9441 VCC.n9436 4.5005
R40542 VCC.n9968 VCC.n9967 4.5005
R40543 VCC.n9878 VCC.n9877 4.5005
R40544 VCC.n9484 VCC.n9482 4.5005
R40545 VCC.n9903 VCC.n9902 4.5005
R40546 VCC.n9470 VCC.n9468 4.5005
R40547 VCC.n9468 VCC.n9467 4.5005
R40548 VCC.n9472 VCC.n9471 4.5005
R40549 VCC.n9886 VCC.n9474 4.5005
R40550 VCC.n9891 VCC.n9890 4.5005
R40551 VCC.n9875 VCC.n9874 4.5005
R40552 VCC.n9880 VCC.n9879 4.5005
R40553 VCC.n9443 VCC.n9442 4.5005
R40554 VCC.n9954 VCC.n9443 4.5005
R40555 VCC.n9942 VCC.n9941 4.5005
R40556 VCC.n9453 VCC.n9440 4.5005
R40557 VCC.n9932 VCC.n9931 4.5005
R40558 VCC.n9462 VCC.n9460 4.5005
R40559 VCC.n9933 VCC.n9455 4.5005
R40560 VCC.n9943 VCC.n9451 4.5005
R40561 VCC.n9945 VCC.n9944 4.5005
R40562 VCC.n9945 VCC.n9449 4.5005
R40563 VCC.n9966 VCC.n9435 4.5005
R40564 VCC.n9977 VCC.n9976 4.5005
R40565 VCC.n9477 VCC.n9475 4.5005
R40566 VCC.n10435 VCC.n10037 4.5005
R40567 VCC.n10438 VCC.n10437 4.5005
R40568 VCC.n10512 VCC.n9992 4.5005
R40569 VCC.n10514 VCC.n10513 4.5005
R40570 VCC.n10009 VCC.n10008 4.5005
R40571 VCC.n10029 VCC.n10027 4.5005
R40572 VCC.n10039 VCC.n10026 4.5005
R40573 VCC.n10468 VCC.n10467 4.5005
R40574 VCC.n10477 VCC.n10476 4.5005
R40575 VCC.n10020 VCC.n10019 4.5005
R40576 VCC.n10000 VCC.n9999 4.5005
R40577 VCC.n10503 VCC.n10502 4.5005
R40578 VCC.n10515 VCC.n9990 4.5005
R40579 VCC.n10004 VCC.n10002 4.5005
R40580 VCC.n10475 VCC.n10474 4.5005
R40581 VCC.n10436 VCC.n10434 4.5005
R40582 VCC.n10432 VCC.n10431 4.5005
R40583 VCC.n10447 VCC.n10038 4.5005
R40584 VCC.n10517 VCC.n10516 4.5005
R40585 VCC.n10517 VCC.n9988 4.5005
R40586 VCC.n10007 VCC.n10005 4.5005
R40587 VCC.n10012 VCC.n10005 4.5005
R40588 VCC.n10463 VCC.n10462 4.5005
R40589 VCC.n10464 VCC.n10463 4.5005
R40590 VCC.n10530 VCC.n10529 4.5005
R40591 VCC.n10417 VCC.n10054 4.5005
R40592 VCC.n10416 VCC.n10415 4.5005
R40593 VCC.n10381 VCC.n10066 4.5005
R40594 VCC.n10335 VCC.n10334 4.5005
R40595 VCC.n10309 VCC.n10308 4.5005
R40596 VCC.n10304 VCC.n10300 4.5005
R40597 VCC.n10310 VCC.n10106 4.5005
R40598 VCC.n10106 VCC.n10104 4.5005
R40599 VCC.n10428 VCC.n10427 4.5005
R40600 VCC.n10383 VCC.n10382 4.5005
R40601 VCC.n10303 VCC.n10302 4.5005
R40602 VCC.n10097 VCC.n10093 4.5005
R40603 VCC.n10320 VCC.n10097 4.5005
R40604 VCC.n10333 VCC.n10332 4.5005
R40605 VCC.n10348 VCC.n10347 4.5005
R40606 VCC.n10347 VCC.n10346 4.5005
R40607 VCC.n10363 VCC.n10362 4.5005
R40608 VCC.n10364 VCC.n10363 4.5005
R40609 VCC.n10355 VCC.n10076 4.5005
R40610 VCC.n10366 VCC.n10076 4.5005
R40611 VCC.n10370 VCC.n10068 4.5005
R40612 VCC.n10371 VCC.n10370 4.5005
R40613 VCC.n10391 VCC.n10390 4.5005
R40614 VCC.n10392 VCC.n10391 4.5005
R40615 VCC.n10419 VCC.n10418 4.5005
R40616 VCC.n10057 VCC.n10055 4.5005
R40617 VCC.n10412 VCC.n10057 4.5005
R40618 VCC.n10282 VCC.n10116 4.5005
R40619 VCC.n10281 VCC.n10280 4.5005
R40620 VCC.n10255 VCC.n10127 4.5005
R40621 VCC.n10220 VCC.n10219 4.5005
R40622 VCC.n10185 VCC.n10184 4.5005
R40623 VCC.n10181 VCC.n10178 4.5005
R40624 VCC.n10187 VCC.n10186 4.5005
R40625 VCC.n10188 VCC.n10187 4.5005
R40626 VCC.n10293 VCC.n10292 4.5005
R40627 VCC.n10257 VCC.n10256 4.5005
R40628 VCC.n10180 VCC.n10179 4.5005
R40629 VCC.n10202 VCC.n10155 4.5005
R40630 VCC.n10202 VCC.n10165 4.5005
R40631 VCC.n10217 VCC.n10156 4.5005
R40632 VCC.n10227 VCC.n10226 4.5005
R40633 VCC.n10228 VCC.n10227 4.5005
R40634 VCC.n10232 VCC.n10147 4.5005
R40635 VCC.n10232 VCC.n10136 4.5005
R40636 VCC.n10235 VCC.n10148 4.5005
R40637 VCC.n10243 VCC.n10242 4.5005
R40638 VCC.n10244 VCC.n10243 4.5005
R40639 VCC.n10139 VCC.n10129 4.5005
R40640 VCC.n10140 VCC.n10139 4.5005
R40641 VCC.n10265 VCC.n10264 4.5005
R40642 VCC.n10266 VCC.n10265 4.5005
R40643 VCC.n10284 VCC.n10283 4.5005
R40644 VCC.n10119 VCC.n10117 4.5005
R40645 VCC.n10277 VCC.n10119 4.5005
R40646 VCC.n10832 VCC.n10666 4.5005
R40647 VCC.n10831 VCC.n10830 4.5005
R40648 VCC.n10735 VCC.n10734 4.5005
R40649 VCC.n10731 VCC.n10728 4.5005
R40650 VCC.n10767 VCC.n10706 4.5005
R40651 VCC.n10777 VCC.n10776 4.5005
R40652 VCC.n10778 VCC.n10777 4.5005
R40653 VCC.n10730 VCC.n10729 4.5005
R40654 VCC.n10752 VCC.n10705 4.5005
R40655 VCC.n10752 VCC.n10715 4.5005
R40656 VCC.n10737 VCC.n10736 4.5005
R40657 VCC.n10738 VCC.n10737 4.5005
R40658 VCC.n10782 VCC.n10697 4.5005
R40659 VCC.n10782 VCC.n10686 4.5005
R40660 VCC.n10843 VCC.n10842 4.5005
R40661 VCC.n10807 VCC.n10806 4.5005
R40662 VCC.n10805 VCC.n10677 4.5005
R40663 VCC.n10785 VCC.n10698 4.5005
R40664 VCC.n10793 VCC.n10792 4.5005
R40665 VCC.n10794 VCC.n10793 4.5005
R40666 VCC.n10689 VCC.n10679 4.5005
R40667 VCC.n10690 VCC.n10689 4.5005
R40668 VCC.n10815 VCC.n10814 4.5005
R40669 VCC.n10816 VCC.n10815 4.5005
R40670 VCC.n10834 VCC.n10833 4.5005
R40671 VCC.n10669 VCC.n10667 4.5005
R40672 VCC.n10827 VCC.n10669 4.5005
R40673 VCC.n10770 VCC.n10769 4.5005
R40674 VCC.n10967 VCC.n10605 4.5005
R40675 VCC.n10966 VCC.n10965 4.5005
R40676 VCC.n10860 VCC.n10859 4.5005
R40677 VCC.n10855 VCC.n10852 4.5005
R40678 VCC.n10884 VCC.n10883 4.5005
R40679 VCC.n10854 VCC.n10853 4.5005
R40680 VCC.n10978 VCC.n10977 4.5005
R40681 VCC.n10934 VCC.n10933 4.5005
R40682 VCC.n10932 VCC.n10617 4.5005
R40683 VCC.n10969 VCC.n10968 4.5005
R40684 VCC.n10886 VCC.n10885 4.5005
R40685 VCC.n10899 VCC.n10898 4.5005
R40686 VCC.n10898 VCC.n10897 4.5005
R40687 VCC.n10648 VCC.n10644 4.5005
R40688 VCC.n10871 VCC.n10648 4.5005
R40689 VCC.n10862 VCC.n10861 4.5005
R40690 VCC.n10862 VCC.n10655 4.5005
R40691 VCC.n10914 VCC.n10913 4.5005
R40692 VCC.n10915 VCC.n10914 4.5005
R40693 VCC.n10906 VCC.n10627 4.5005
R40694 VCC.n10917 VCC.n10627 4.5005
R40695 VCC.n10921 VCC.n10619 4.5005
R40696 VCC.n10922 VCC.n10921 4.5005
R40697 VCC.n10942 VCC.n10941 4.5005
R40698 VCC.n10943 VCC.n10942 4.5005
R40699 VCC.n10608 VCC.n10606 4.5005
R40700 VCC.n10962 VCC.n10608 4.5005
R40701 VCC.n10548 VCC.n10543 4.5005
R40702 VCC.n11075 VCC.n11074 4.5005
R40703 VCC.n10985 VCC.n10984 4.5005
R40704 VCC.n10591 VCC.n10589 4.5005
R40705 VCC.n11010 VCC.n11009 4.5005
R40706 VCC.n10577 VCC.n10575 4.5005
R40707 VCC.n10575 VCC.n10574 4.5005
R40708 VCC.n10579 VCC.n10578 4.5005
R40709 VCC.n10993 VCC.n10581 4.5005
R40710 VCC.n10998 VCC.n10997 4.5005
R40711 VCC.n10982 VCC.n10981 4.5005
R40712 VCC.n10987 VCC.n10986 4.5005
R40713 VCC.n10550 VCC.n10549 4.5005
R40714 VCC.n11061 VCC.n10550 4.5005
R40715 VCC.n11049 VCC.n11048 4.5005
R40716 VCC.n10560 VCC.n10547 4.5005
R40717 VCC.n11039 VCC.n11038 4.5005
R40718 VCC.n10569 VCC.n10567 4.5005
R40719 VCC.n11040 VCC.n10562 4.5005
R40720 VCC.n11050 VCC.n10558 4.5005
R40721 VCC.n11052 VCC.n11051 4.5005
R40722 VCC.n11052 VCC.n10556 4.5005
R40723 VCC.n11073 VCC.n10542 4.5005
R40724 VCC.n11084 VCC.n11083 4.5005
R40725 VCC.n10584 VCC.n10582 4.5005
R40726 VCC.n11542 VCC.n11144 4.5005
R40727 VCC.n11545 VCC.n11544 4.5005
R40728 VCC.n11619 VCC.n11099 4.5005
R40729 VCC.n11621 VCC.n11620 4.5005
R40730 VCC.n11116 VCC.n11115 4.5005
R40731 VCC.n11136 VCC.n11134 4.5005
R40732 VCC.n11146 VCC.n11133 4.5005
R40733 VCC.n11575 VCC.n11574 4.5005
R40734 VCC.n11584 VCC.n11583 4.5005
R40735 VCC.n11127 VCC.n11126 4.5005
R40736 VCC.n11107 VCC.n11106 4.5005
R40737 VCC.n11610 VCC.n11609 4.5005
R40738 VCC.n11622 VCC.n11097 4.5005
R40739 VCC.n11111 VCC.n11109 4.5005
R40740 VCC.n11582 VCC.n11581 4.5005
R40741 VCC.n11543 VCC.n11541 4.5005
R40742 VCC.n11539 VCC.n11538 4.5005
R40743 VCC.n11554 VCC.n11145 4.5005
R40744 VCC.n11624 VCC.n11623 4.5005
R40745 VCC.n11624 VCC.n11095 4.5005
R40746 VCC.n11114 VCC.n11112 4.5005
R40747 VCC.n11119 VCC.n11112 4.5005
R40748 VCC.n11570 VCC.n11569 4.5005
R40749 VCC.n11571 VCC.n11570 4.5005
R40750 VCC.n11637 VCC.n11636 4.5005
R40751 VCC.n11524 VCC.n11161 4.5005
R40752 VCC.n11523 VCC.n11522 4.5005
R40753 VCC.n11488 VCC.n11173 4.5005
R40754 VCC.n11442 VCC.n11441 4.5005
R40755 VCC.n11416 VCC.n11415 4.5005
R40756 VCC.n11411 VCC.n11407 4.5005
R40757 VCC.n11417 VCC.n11213 4.5005
R40758 VCC.n11213 VCC.n11211 4.5005
R40759 VCC.n11535 VCC.n11534 4.5005
R40760 VCC.n11490 VCC.n11489 4.5005
R40761 VCC.n11410 VCC.n11409 4.5005
R40762 VCC.n11204 VCC.n11200 4.5005
R40763 VCC.n11427 VCC.n11204 4.5005
R40764 VCC.n11440 VCC.n11439 4.5005
R40765 VCC.n11455 VCC.n11454 4.5005
R40766 VCC.n11454 VCC.n11453 4.5005
R40767 VCC.n11470 VCC.n11469 4.5005
R40768 VCC.n11471 VCC.n11470 4.5005
R40769 VCC.n11462 VCC.n11183 4.5005
R40770 VCC.n11473 VCC.n11183 4.5005
R40771 VCC.n11477 VCC.n11175 4.5005
R40772 VCC.n11478 VCC.n11477 4.5005
R40773 VCC.n11498 VCC.n11497 4.5005
R40774 VCC.n11499 VCC.n11498 4.5005
R40775 VCC.n11526 VCC.n11525 4.5005
R40776 VCC.n11164 VCC.n11162 4.5005
R40777 VCC.n11519 VCC.n11164 4.5005
R40778 VCC.n11389 VCC.n11223 4.5005
R40779 VCC.n11388 VCC.n11387 4.5005
R40780 VCC.n11362 VCC.n11234 4.5005
R40781 VCC.n11327 VCC.n11326 4.5005
R40782 VCC.n11292 VCC.n11291 4.5005
R40783 VCC.n11288 VCC.n11285 4.5005
R40784 VCC.n11294 VCC.n11293 4.5005
R40785 VCC.n11295 VCC.n11294 4.5005
R40786 VCC.n11400 VCC.n11399 4.5005
R40787 VCC.n11364 VCC.n11363 4.5005
R40788 VCC.n11287 VCC.n11286 4.5005
R40789 VCC.n11309 VCC.n11262 4.5005
R40790 VCC.n11309 VCC.n11272 4.5005
R40791 VCC.n11324 VCC.n11263 4.5005
R40792 VCC.n11334 VCC.n11333 4.5005
R40793 VCC.n11335 VCC.n11334 4.5005
R40794 VCC.n11339 VCC.n11254 4.5005
R40795 VCC.n11339 VCC.n11243 4.5005
R40796 VCC.n11342 VCC.n11255 4.5005
R40797 VCC.n11350 VCC.n11349 4.5005
R40798 VCC.n11351 VCC.n11350 4.5005
R40799 VCC.n11246 VCC.n11236 4.5005
R40800 VCC.n11247 VCC.n11246 4.5005
R40801 VCC.n11372 VCC.n11371 4.5005
R40802 VCC.n11373 VCC.n11372 4.5005
R40803 VCC.n11391 VCC.n11390 4.5005
R40804 VCC.n11226 VCC.n11224 4.5005
R40805 VCC.n11384 VCC.n11226 4.5005
R40806 VCC.n11939 VCC.n11773 4.5005
R40807 VCC.n11938 VCC.n11937 4.5005
R40808 VCC.n11842 VCC.n11841 4.5005
R40809 VCC.n11838 VCC.n11835 4.5005
R40810 VCC.n11874 VCC.n11813 4.5005
R40811 VCC.n11884 VCC.n11883 4.5005
R40812 VCC.n11885 VCC.n11884 4.5005
R40813 VCC.n11837 VCC.n11836 4.5005
R40814 VCC.n11859 VCC.n11812 4.5005
R40815 VCC.n11859 VCC.n11822 4.5005
R40816 VCC.n11844 VCC.n11843 4.5005
R40817 VCC.n11845 VCC.n11844 4.5005
R40818 VCC.n11889 VCC.n11804 4.5005
R40819 VCC.n11889 VCC.n11793 4.5005
R40820 VCC.n11950 VCC.n11949 4.5005
R40821 VCC.n11914 VCC.n11913 4.5005
R40822 VCC.n11912 VCC.n11784 4.5005
R40823 VCC.n11892 VCC.n11805 4.5005
R40824 VCC.n11900 VCC.n11899 4.5005
R40825 VCC.n11901 VCC.n11900 4.5005
R40826 VCC.n11796 VCC.n11786 4.5005
R40827 VCC.n11797 VCC.n11796 4.5005
R40828 VCC.n11922 VCC.n11921 4.5005
R40829 VCC.n11923 VCC.n11922 4.5005
R40830 VCC.n11941 VCC.n11940 4.5005
R40831 VCC.n11776 VCC.n11774 4.5005
R40832 VCC.n11934 VCC.n11776 4.5005
R40833 VCC.n11877 VCC.n11876 4.5005
R40834 VCC.n12074 VCC.n11712 4.5005
R40835 VCC.n12073 VCC.n12072 4.5005
R40836 VCC.n11967 VCC.n11966 4.5005
R40837 VCC.n11962 VCC.n11959 4.5005
R40838 VCC.n11991 VCC.n11990 4.5005
R40839 VCC.n11961 VCC.n11960 4.5005
R40840 VCC.n12085 VCC.n12084 4.5005
R40841 VCC.n12041 VCC.n12040 4.5005
R40842 VCC.n12039 VCC.n11724 4.5005
R40843 VCC.n12076 VCC.n12075 4.5005
R40844 VCC.n11993 VCC.n11992 4.5005
R40845 VCC.n12006 VCC.n12005 4.5005
R40846 VCC.n12005 VCC.n12004 4.5005
R40847 VCC.n11755 VCC.n11751 4.5005
R40848 VCC.n11978 VCC.n11755 4.5005
R40849 VCC.n11969 VCC.n11968 4.5005
R40850 VCC.n11969 VCC.n11762 4.5005
R40851 VCC.n12021 VCC.n12020 4.5005
R40852 VCC.n12022 VCC.n12021 4.5005
R40853 VCC.n12013 VCC.n11734 4.5005
R40854 VCC.n12024 VCC.n11734 4.5005
R40855 VCC.n12028 VCC.n11726 4.5005
R40856 VCC.n12029 VCC.n12028 4.5005
R40857 VCC.n12049 VCC.n12048 4.5005
R40858 VCC.n12050 VCC.n12049 4.5005
R40859 VCC.n11715 VCC.n11713 4.5005
R40860 VCC.n12069 VCC.n11715 4.5005
R40861 VCC.n11655 VCC.n11650 4.5005
R40862 VCC.n12182 VCC.n12181 4.5005
R40863 VCC.n12092 VCC.n12091 4.5005
R40864 VCC.n11698 VCC.n11696 4.5005
R40865 VCC.n12117 VCC.n12116 4.5005
R40866 VCC.n11684 VCC.n11682 4.5005
R40867 VCC.n11682 VCC.n11681 4.5005
R40868 VCC.n11686 VCC.n11685 4.5005
R40869 VCC.n12100 VCC.n11688 4.5005
R40870 VCC.n12105 VCC.n12104 4.5005
R40871 VCC.n12089 VCC.n12088 4.5005
R40872 VCC.n12094 VCC.n12093 4.5005
R40873 VCC.n11657 VCC.n11656 4.5005
R40874 VCC.n12168 VCC.n11657 4.5005
R40875 VCC.n12156 VCC.n12155 4.5005
R40876 VCC.n11667 VCC.n11654 4.5005
R40877 VCC.n12146 VCC.n12145 4.5005
R40878 VCC.n11676 VCC.n11674 4.5005
R40879 VCC.n12147 VCC.n11669 4.5005
R40880 VCC.n12157 VCC.n11665 4.5005
R40881 VCC.n12159 VCC.n12158 4.5005
R40882 VCC.n12159 VCC.n11663 4.5005
R40883 VCC.n12180 VCC.n11649 4.5005
R40884 VCC.n12191 VCC.n12190 4.5005
R40885 VCC.n11691 VCC.n11689 4.5005
R40886 VCC.n12649 VCC.n12251 4.5005
R40887 VCC.n12652 VCC.n12651 4.5005
R40888 VCC.n12726 VCC.n12206 4.5005
R40889 VCC.n12728 VCC.n12727 4.5005
R40890 VCC.n12223 VCC.n12222 4.5005
R40891 VCC.n12243 VCC.n12241 4.5005
R40892 VCC.n12253 VCC.n12240 4.5005
R40893 VCC.n12682 VCC.n12681 4.5005
R40894 VCC.n12691 VCC.n12690 4.5005
R40895 VCC.n12234 VCC.n12233 4.5005
R40896 VCC.n12214 VCC.n12213 4.5005
R40897 VCC.n12717 VCC.n12716 4.5005
R40898 VCC.n12729 VCC.n12204 4.5005
R40899 VCC.n12218 VCC.n12216 4.5005
R40900 VCC.n12689 VCC.n12688 4.5005
R40901 VCC.n12650 VCC.n12648 4.5005
R40902 VCC.n12646 VCC.n12645 4.5005
R40903 VCC.n12661 VCC.n12252 4.5005
R40904 VCC.n12731 VCC.n12730 4.5005
R40905 VCC.n12731 VCC.n12202 4.5005
R40906 VCC.n12221 VCC.n12219 4.5005
R40907 VCC.n12226 VCC.n12219 4.5005
R40908 VCC.n12677 VCC.n12676 4.5005
R40909 VCC.n12678 VCC.n12677 4.5005
R40910 VCC.n12744 VCC.n12743 4.5005
R40911 VCC.n12631 VCC.n12268 4.5005
R40912 VCC.n12630 VCC.n12629 4.5005
R40913 VCC.n12595 VCC.n12280 4.5005
R40914 VCC.n12549 VCC.n12548 4.5005
R40915 VCC.n12523 VCC.n12522 4.5005
R40916 VCC.n12518 VCC.n12514 4.5005
R40917 VCC.n12524 VCC.n12320 4.5005
R40918 VCC.n12320 VCC.n12318 4.5005
R40919 VCC.n12642 VCC.n12641 4.5005
R40920 VCC.n12597 VCC.n12596 4.5005
R40921 VCC.n12517 VCC.n12516 4.5005
R40922 VCC.n12311 VCC.n12307 4.5005
R40923 VCC.n12534 VCC.n12311 4.5005
R40924 VCC.n12547 VCC.n12546 4.5005
R40925 VCC.n12562 VCC.n12561 4.5005
R40926 VCC.n12561 VCC.n12560 4.5005
R40927 VCC.n12577 VCC.n12576 4.5005
R40928 VCC.n12578 VCC.n12577 4.5005
R40929 VCC.n12569 VCC.n12290 4.5005
R40930 VCC.n12580 VCC.n12290 4.5005
R40931 VCC.n12584 VCC.n12282 4.5005
R40932 VCC.n12585 VCC.n12584 4.5005
R40933 VCC.n12605 VCC.n12604 4.5005
R40934 VCC.n12606 VCC.n12605 4.5005
R40935 VCC.n12633 VCC.n12632 4.5005
R40936 VCC.n12271 VCC.n12269 4.5005
R40937 VCC.n12626 VCC.n12271 4.5005
R40938 VCC.n12496 VCC.n12330 4.5005
R40939 VCC.n12495 VCC.n12494 4.5005
R40940 VCC.n12469 VCC.n12341 4.5005
R40941 VCC.n12434 VCC.n12433 4.5005
R40942 VCC.n12399 VCC.n12398 4.5005
R40943 VCC.n12395 VCC.n12392 4.5005
R40944 VCC.n12401 VCC.n12400 4.5005
R40945 VCC.n12402 VCC.n12401 4.5005
R40946 VCC.n12507 VCC.n12506 4.5005
R40947 VCC.n12471 VCC.n12470 4.5005
R40948 VCC.n12394 VCC.n12393 4.5005
R40949 VCC.n12416 VCC.n12369 4.5005
R40950 VCC.n12416 VCC.n12379 4.5005
R40951 VCC.n12431 VCC.n12370 4.5005
R40952 VCC.n12441 VCC.n12440 4.5005
R40953 VCC.n12442 VCC.n12441 4.5005
R40954 VCC.n12446 VCC.n12361 4.5005
R40955 VCC.n12446 VCC.n12350 4.5005
R40956 VCC.n12449 VCC.n12362 4.5005
R40957 VCC.n12457 VCC.n12456 4.5005
R40958 VCC.n12458 VCC.n12457 4.5005
R40959 VCC.n12353 VCC.n12343 4.5005
R40960 VCC.n12354 VCC.n12353 4.5005
R40961 VCC.n12479 VCC.n12478 4.5005
R40962 VCC.n12480 VCC.n12479 4.5005
R40963 VCC.n12498 VCC.n12497 4.5005
R40964 VCC.n12333 VCC.n12331 4.5005
R40965 VCC.n12491 VCC.n12333 4.5005
R40966 VCC.n13046 VCC.n12880 4.5005
R40967 VCC.n13045 VCC.n13044 4.5005
R40968 VCC.n12949 VCC.n12948 4.5005
R40969 VCC.n12945 VCC.n12942 4.5005
R40970 VCC.n12981 VCC.n12920 4.5005
R40971 VCC.n12991 VCC.n12990 4.5005
R40972 VCC.n12992 VCC.n12991 4.5005
R40973 VCC.n12944 VCC.n12943 4.5005
R40974 VCC.n12966 VCC.n12919 4.5005
R40975 VCC.n12966 VCC.n12929 4.5005
R40976 VCC.n12951 VCC.n12950 4.5005
R40977 VCC.n12952 VCC.n12951 4.5005
R40978 VCC.n12996 VCC.n12911 4.5005
R40979 VCC.n12996 VCC.n12900 4.5005
R40980 VCC.n13057 VCC.n13056 4.5005
R40981 VCC.n13021 VCC.n13020 4.5005
R40982 VCC.n13019 VCC.n12891 4.5005
R40983 VCC.n12999 VCC.n12912 4.5005
R40984 VCC.n13007 VCC.n13006 4.5005
R40985 VCC.n13008 VCC.n13007 4.5005
R40986 VCC.n12903 VCC.n12893 4.5005
R40987 VCC.n12904 VCC.n12903 4.5005
R40988 VCC.n13029 VCC.n13028 4.5005
R40989 VCC.n13030 VCC.n13029 4.5005
R40990 VCC.n13048 VCC.n13047 4.5005
R40991 VCC.n12883 VCC.n12881 4.5005
R40992 VCC.n13041 VCC.n12883 4.5005
R40993 VCC.n12984 VCC.n12983 4.5005
R40994 VCC.n13181 VCC.n12819 4.5005
R40995 VCC.n13180 VCC.n13179 4.5005
R40996 VCC.n13074 VCC.n13073 4.5005
R40997 VCC.n13069 VCC.n13066 4.5005
R40998 VCC.n13098 VCC.n13097 4.5005
R40999 VCC.n13068 VCC.n13067 4.5005
R41000 VCC.n13192 VCC.n13191 4.5005
R41001 VCC.n13148 VCC.n13147 4.5005
R41002 VCC.n13146 VCC.n12831 4.5005
R41003 VCC.n13183 VCC.n13182 4.5005
R41004 VCC.n13100 VCC.n13099 4.5005
R41005 VCC.n13113 VCC.n13112 4.5005
R41006 VCC.n13112 VCC.n13111 4.5005
R41007 VCC.n12862 VCC.n12858 4.5005
R41008 VCC.n13085 VCC.n12862 4.5005
R41009 VCC.n13076 VCC.n13075 4.5005
R41010 VCC.n13076 VCC.n12869 4.5005
R41011 VCC.n13128 VCC.n13127 4.5005
R41012 VCC.n13129 VCC.n13128 4.5005
R41013 VCC.n13120 VCC.n12841 4.5005
R41014 VCC.n13131 VCC.n12841 4.5005
R41015 VCC.n13135 VCC.n12833 4.5005
R41016 VCC.n13136 VCC.n13135 4.5005
R41017 VCC.n13156 VCC.n13155 4.5005
R41018 VCC.n13157 VCC.n13156 4.5005
R41019 VCC.n12822 VCC.n12820 4.5005
R41020 VCC.n13176 VCC.n12822 4.5005
R41021 VCC.n12762 VCC.n12757 4.5005
R41022 VCC.n13289 VCC.n13288 4.5005
R41023 VCC.n13199 VCC.n13198 4.5005
R41024 VCC.n12805 VCC.n12803 4.5005
R41025 VCC.n13224 VCC.n13223 4.5005
R41026 VCC.n12791 VCC.n12789 4.5005
R41027 VCC.n12789 VCC.n12788 4.5005
R41028 VCC.n12793 VCC.n12792 4.5005
R41029 VCC.n13207 VCC.n12795 4.5005
R41030 VCC.n13212 VCC.n13211 4.5005
R41031 VCC.n13196 VCC.n13195 4.5005
R41032 VCC.n13201 VCC.n13200 4.5005
R41033 VCC.n12764 VCC.n12763 4.5005
R41034 VCC.n13275 VCC.n12764 4.5005
R41035 VCC.n13263 VCC.n13262 4.5005
R41036 VCC.n12774 VCC.n12761 4.5005
R41037 VCC.n13253 VCC.n13252 4.5005
R41038 VCC.n12783 VCC.n12781 4.5005
R41039 VCC.n13254 VCC.n12776 4.5005
R41040 VCC.n13264 VCC.n12772 4.5005
R41041 VCC.n13266 VCC.n13265 4.5005
R41042 VCC.n13266 VCC.n12770 4.5005
R41043 VCC.n13287 VCC.n12756 4.5005
R41044 VCC.n13298 VCC.n13297 4.5005
R41045 VCC.n12798 VCC.n12796 4.5005
R41046 VCC.n13756 VCC.n13358 4.5005
R41047 VCC.n13759 VCC.n13758 4.5005
R41048 VCC.n13833 VCC.n13313 4.5005
R41049 VCC.n13835 VCC.n13834 4.5005
R41050 VCC.n13330 VCC.n13329 4.5005
R41051 VCC.n13350 VCC.n13348 4.5005
R41052 VCC.n13360 VCC.n13347 4.5005
R41053 VCC.n13789 VCC.n13788 4.5005
R41054 VCC.n13798 VCC.n13797 4.5005
R41055 VCC.n13341 VCC.n13340 4.5005
R41056 VCC.n13321 VCC.n13320 4.5005
R41057 VCC.n13824 VCC.n13823 4.5005
R41058 VCC.n13836 VCC.n13311 4.5005
R41059 VCC.n13325 VCC.n13323 4.5005
R41060 VCC.n13796 VCC.n13795 4.5005
R41061 VCC.n13757 VCC.n13755 4.5005
R41062 VCC.n13753 VCC.n13752 4.5005
R41063 VCC.n13768 VCC.n13359 4.5005
R41064 VCC.n13838 VCC.n13837 4.5005
R41065 VCC.n13838 VCC.n13309 4.5005
R41066 VCC.n13328 VCC.n13326 4.5005
R41067 VCC.n13333 VCC.n13326 4.5005
R41068 VCC.n13784 VCC.n13783 4.5005
R41069 VCC.n13785 VCC.n13784 4.5005
R41070 VCC.n13851 VCC.n13850 4.5005
R41071 VCC.n13738 VCC.n13375 4.5005
R41072 VCC.n13737 VCC.n13736 4.5005
R41073 VCC.n13702 VCC.n13387 4.5005
R41074 VCC.n13656 VCC.n13655 4.5005
R41075 VCC.n13630 VCC.n13629 4.5005
R41076 VCC.n13625 VCC.n13621 4.5005
R41077 VCC.n13631 VCC.n13427 4.5005
R41078 VCC.n13427 VCC.n13425 4.5005
R41079 VCC.n13749 VCC.n13748 4.5005
R41080 VCC.n13704 VCC.n13703 4.5005
R41081 VCC.n13624 VCC.n13623 4.5005
R41082 VCC.n13418 VCC.n13414 4.5005
R41083 VCC.n13641 VCC.n13418 4.5005
R41084 VCC.n13654 VCC.n13653 4.5005
R41085 VCC.n13669 VCC.n13668 4.5005
R41086 VCC.n13668 VCC.n13667 4.5005
R41087 VCC.n13684 VCC.n13683 4.5005
R41088 VCC.n13685 VCC.n13684 4.5005
R41089 VCC.n13676 VCC.n13397 4.5005
R41090 VCC.n13687 VCC.n13397 4.5005
R41091 VCC.n13691 VCC.n13389 4.5005
R41092 VCC.n13692 VCC.n13691 4.5005
R41093 VCC.n13712 VCC.n13711 4.5005
R41094 VCC.n13713 VCC.n13712 4.5005
R41095 VCC.n13740 VCC.n13739 4.5005
R41096 VCC.n13378 VCC.n13376 4.5005
R41097 VCC.n13733 VCC.n13378 4.5005
R41098 VCC.n13603 VCC.n13437 4.5005
R41099 VCC.n13602 VCC.n13601 4.5005
R41100 VCC.n13576 VCC.n13448 4.5005
R41101 VCC.n13541 VCC.n13540 4.5005
R41102 VCC.n13506 VCC.n13505 4.5005
R41103 VCC.n13502 VCC.n13499 4.5005
R41104 VCC.n13508 VCC.n13507 4.5005
R41105 VCC.n13509 VCC.n13508 4.5005
R41106 VCC.n13614 VCC.n13613 4.5005
R41107 VCC.n13578 VCC.n13577 4.5005
R41108 VCC.n13501 VCC.n13500 4.5005
R41109 VCC.n13523 VCC.n13476 4.5005
R41110 VCC.n13523 VCC.n13486 4.5005
R41111 VCC.n13538 VCC.n13477 4.5005
R41112 VCC.n13548 VCC.n13547 4.5005
R41113 VCC.n13549 VCC.n13548 4.5005
R41114 VCC.n13553 VCC.n13468 4.5005
R41115 VCC.n13553 VCC.n13457 4.5005
R41116 VCC.n13556 VCC.n13469 4.5005
R41117 VCC.n13564 VCC.n13563 4.5005
R41118 VCC.n13565 VCC.n13564 4.5005
R41119 VCC.n13460 VCC.n13450 4.5005
R41120 VCC.n13461 VCC.n13460 4.5005
R41121 VCC.n13586 VCC.n13585 4.5005
R41122 VCC.n13587 VCC.n13586 4.5005
R41123 VCC.n13605 VCC.n13604 4.5005
R41124 VCC.n13440 VCC.n13438 4.5005
R41125 VCC.n13598 VCC.n13440 4.5005
R41126 VCC.n14153 VCC.n13987 4.5005
R41127 VCC.n14152 VCC.n14151 4.5005
R41128 VCC.n14056 VCC.n14055 4.5005
R41129 VCC.n14052 VCC.n14049 4.5005
R41130 VCC.n14088 VCC.n14027 4.5005
R41131 VCC.n14098 VCC.n14097 4.5005
R41132 VCC.n14099 VCC.n14098 4.5005
R41133 VCC.n14051 VCC.n14050 4.5005
R41134 VCC.n14073 VCC.n14026 4.5005
R41135 VCC.n14073 VCC.n14036 4.5005
R41136 VCC.n14058 VCC.n14057 4.5005
R41137 VCC.n14059 VCC.n14058 4.5005
R41138 VCC.n14103 VCC.n14018 4.5005
R41139 VCC.n14103 VCC.n14007 4.5005
R41140 VCC.n14164 VCC.n14163 4.5005
R41141 VCC.n14128 VCC.n14127 4.5005
R41142 VCC.n14126 VCC.n13998 4.5005
R41143 VCC.n14106 VCC.n14019 4.5005
R41144 VCC.n14114 VCC.n14113 4.5005
R41145 VCC.n14115 VCC.n14114 4.5005
R41146 VCC.n14010 VCC.n14000 4.5005
R41147 VCC.n14011 VCC.n14010 4.5005
R41148 VCC.n14136 VCC.n14135 4.5005
R41149 VCC.n14137 VCC.n14136 4.5005
R41150 VCC.n14155 VCC.n14154 4.5005
R41151 VCC.n13990 VCC.n13988 4.5005
R41152 VCC.n14148 VCC.n13990 4.5005
R41153 VCC.n14091 VCC.n14090 4.5005
R41154 VCC.n14288 VCC.n13926 4.5005
R41155 VCC.n14287 VCC.n14286 4.5005
R41156 VCC.n14181 VCC.n14180 4.5005
R41157 VCC.n14176 VCC.n14173 4.5005
R41158 VCC.n14205 VCC.n14204 4.5005
R41159 VCC.n14175 VCC.n14174 4.5005
R41160 VCC.n14299 VCC.n14298 4.5005
R41161 VCC.n14255 VCC.n14254 4.5005
R41162 VCC.n14253 VCC.n13938 4.5005
R41163 VCC.n14290 VCC.n14289 4.5005
R41164 VCC.n14207 VCC.n14206 4.5005
R41165 VCC.n14220 VCC.n14219 4.5005
R41166 VCC.n14219 VCC.n14218 4.5005
R41167 VCC.n13969 VCC.n13965 4.5005
R41168 VCC.n14192 VCC.n13969 4.5005
R41169 VCC.n14183 VCC.n14182 4.5005
R41170 VCC.n14183 VCC.n13976 4.5005
R41171 VCC.n14235 VCC.n14234 4.5005
R41172 VCC.n14236 VCC.n14235 4.5005
R41173 VCC.n14227 VCC.n13948 4.5005
R41174 VCC.n14238 VCC.n13948 4.5005
R41175 VCC.n14242 VCC.n13940 4.5005
R41176 VCC.n14243 VCC.n14242 4.5005
R41177 VCC.n14263 VCC.n14262 4.5005
R41178 VCC.n14264 VCC.n14263 4.5005
R41179 VCC.n13929 VCC.n13927 4.5005
R41180 VCC.n14283 VCC.n13929 4.5005
R41181 VCC.n13869 VCC.n13864 4.5005
R41182 VCC.n14396 VCC.n14395 4.5005
R41183 VCC.n14306 VCC.n14305 4.5005
R41184 VCC.n13912 VCC.n13910 4.5005
R41185 VCC.n14331 VCC.n14330 4.5005
R41186 VCC.n13898 VCC.n13896 4.5005
R41187 VCC.n13896 VCC.n13895 4.5005
R41188 VCC.n13900 VCC.n13899 4.5005
R41189 VCC.n14314 VCC.n13902 4.5005
R41190 VCC.n14319 VCC.n14318 4.5005
R41191 VCC.n14303 VCC.n14302 4.5005
R41192 VCC.n14308 VCC.n14307 4.5005
R41193 VCC.n13871 VCC.n13870 4.5005
R41194 VCC.n14382 VCC.n13871 4.5005
R41195 VCC.n14370 VCC.n14369 4.5005
R41196 VCC.n13881 VCC.n13868 4.5005
R41197 VCC.n14360 VCC.n14359 4.5005
R41198 VCC.n13890 VCC.n13888 4.5005
R41199 VCC.n14361 VCC.n13883 4.5005
R41200 VCC.n14371 VCC.n13879 4.5005
R41201 VCC.n14373 VCC.n14372 4.5005
R41202 VCC.n14373 VCC.n13877 4.5005
R41203 VCC.n14394 VCC.n13863 4.5005
R41204 VCC.n14405 VCC.n14404 4.5005
R41205 VCC.n13905 VCC.n13903 4.5005
R41206 VCC.n14863 VCC.n14465 4.5005
R41207 VCC.n14866 VCC.n14865 4.5005
R41208 VCC.n14940 VCC.n14420 4.5005
R41209 VCC.n14942 VCC.n14941 4.5005
R41210 VCC.n14437 VCC.n14436 4.5005
R41211 VCC.n14457 VCC.n14455 4.5005
R41212 VCC.n14467 VCC.n14454 4.5005
R41213 VCC.n14896 VCC.n14895 4.5005
R41214 VCC.n14905 VCC.n14904 4.5005
R41215 VCC.n14448 VCC.n14447 4.5005
R41216 VCC.n14428 VCC.n14427 4.5005
R41217 VCC.n14931 VCC.n14930 4.5005
R41218 VCC.n14943 VCC.n14418 4.5005
R41219 VCC.n14432 VCC.n14430 4.5005
R41220 VCC.n14903 VCC.n14902 4.5005
R41221 VCC.n14864 VCC.n14862 4.5005
R41222 VCC.n14860 VCC.n14859 4.5005
R41223 VCC.n14875 VCC.n14466 4.5005
R41224 VCC.n14945 VCC.n14944 4.5005
R41225 VCC.n14945 VCC.n14416 4.5005
R41226 VCC.n14435 VCC.n14433 4.5005
R41227 VCC.n14440 VCC.n14433 4.5005
R41228 VCC.n14891 VCC.n14890 4.5005
R41229 VCC.n14892 VCC.n14891 4.5005
R41230 VCC.n14958 VCC.n14957 4.5005
R41231 VCC.n14845 VCC.n14482 4.5005
R41232 VCC.n14844 VCC.n14843 4.5005
R41233 VCC.n14809 VCC.n14494 4.5005
R41234 VCC.n14763 VCC.n14762 4.5005
R41235 VCC.n14737 VCC.n14736 4.5005
R41236 VCC.n14732 VCC.n14728 4.5005
R41237 VCC.n14738 VCC.n14534 4.5005
R41238 VCC.n14534 VCC.n14532 4.5005
R41239 VCC.n14856 VCC.n14855 4.5005
R41240 VCC.n14811 VCC.n14810 4.5005
R41241 VCC.n14731 VCC.n14730 4.5005
R41242 VCC.n14525 VCC.n14521 4.5005
R41243 VCC.n14748 VCC.n14525 4.5005
R41244 VCC.n14761 VCC.n14760 4.5005
R41245 VCC.n14776 VCC.n14775 4.5005
R41246 VCC.n14775 VCC.n14774 4.5005
R41247 VCC.n14791 VCC.n14790 4.5005
R41248 VCC.n14792 VCC.n14791 4.5005
R41249 VCC.n14783 VCC.n14504 4.5005
R41250 VCC.n14794 VCC.n14504 4.5005
R41251 VCC.n14798 VCC.n14496 4.5005
R41252 VCC.n14799 VCC.n14798 4.5005
R41253 VCC.n14819 VCC.n14818 4.5005
R41254 VCC.n14820 VCC.n14819 4.5005
R41255 VCC.n14847 VCC.n14846 4.5005
R41256 VCC.n14485 VCC.n14483 4.5005
R41257 VCC.n14840 VCC.n14485 4.5005
R41258 VCC.n14710 VCC.n14544 4.5005
R41259 VCC.n14709 VCC.n14708 4.5005
R41260 VCC.n14683 VCC.n14555 4.5005
R41261 VCC.n14648 VCC.n14647 4.5005
R41262 VCC.n14613 VCC.n14612 4.5005
R41263 VCC.n14609 VCC.n14606 4.5005
R41264 VCC.n14615 VCC.n14614 4.5005
R41265 VCC.n14616 VCC.n14615 4.5005
R41266 VCC.n14721 VCC.n14720 4.5005
R41267 VCC.n14685 VCC.n14684 4.5005
R41268 VCC.n14608 VCC.n14607 4.5005
R41269 VCC.n14630 VCC.n14583 4.5005
R41270 VCC.n14630 VCC.n14593 4.5005
R41271 VCC.n14645 VCC.n14584 4.5005
R41272 VCC.n14655 VCC.n14654 4.5005
R41273 VCC.n14656 VCC.n14655 4.5005
R41274 VCC.n14660 VCC.n14575 4.5005
R41275 VCC.n14660 VCC.n14564 4.5005
R41276 VCC.n14663 VCC.n14576 4.5005
R41277 VCC.n14671 VCC.n14670 4.5005
R41278 VCC.n14672 VCC.n14671 4.5005
R41279 VCC.n14567 VCC.n14557 4.5005
R41280 VCC.n14568 VCC.n14567 4.5005
R41281 VCC.n14693 VCC.n14692 4.5005
R41282 VCC.n14694 VCC.n14693 4.5005
R41283 VCC.n14712 VCC.n14711 4.5005
R41284 VCC.n14547 VCC.n14545 4.5005
R41285 VCC.n14705 VCC.n14547 4.5005
R41286 VCC.n15260 VCC.n15094 4.5005
R41287 VCC.n15259 VCC.n15258 4.5005
R41288 VCC.n15163 VCC.n15162 4.5005
R41289 VCC.n15159 VCC.n15156 4.5005
R41290 VCC.n15195 VCC.n15134 4.5005
R41291 VCC.n15205 VCC.n15204 4.5005
R41292 VCC.n15206 VCC.n15205 4.5005
R41293 VCC.n15158 VCC.n15157 4.5005
R41294 VCC.n15180 VCC.n15133 4.5005
R41295 VCC.n15180 VCC.n15143 4.5005
R41296 VCC.n15165 VCC.n15164 4.5005
R41297 VCC.n15166 VCC.n15165 4.5005
R41298 VCC.n15210 VCC.n15125 4.5005
R41299 VCC.n15210 VCC.n15114 4.5005
R41300 VCC.n15271 VCC.n15270 4.5005
R41301 VCC.n15235 VCC.n15234 4.5005
R41302 VCC.n15233 VCC.n15105 4.5005
R41303 VCC.n15213 VCC.n15126 4.5005
R41304 VCC.n15221 VCC.n15220 4.5005
R41305 VCC.n15222 VCC.n15221 4.5005
R41306 VCC.n15117 VCC.n15107 4.5005
R41307 VCC.n15118 VCC.n15117 4.5005
R41308 VCC.n15243 VCC.n15242 4.5005
R41309 VCC.n15244 VCC.n15243 4.5005
R41310 VCC.n15262 VCC.n15261 4.5005
R41311 VCC.n15097 VCC.n15095 4.5005
R41312 VCC.n15255 VCC.n15097 4.5005
R41313 VCC.n15198 VCC.n15197 4.5005
R41314 VCC.n15395 VCC.n15033 4.5005
R41315 VCC.n15394 VCC.n15393 4.5005
R41316 VCC.n15288 VCC.n15287 4.5005
R41317 VCC.n15283 VCC.n15280 4.5005
R41318 VCC.n15312 VCC.n15311 4.5005
R41319 VCC.n15282 VCC.n15281 4.5005
R41320 VCC.n15406 VCC.n15405 4.5005
R41321 VCC.n15362 VCC.n15361 4.5005
R41322 VCC.n15360 VCC.n15045 4.5005
R41323 VCC.n15397 VCC.n15396 4.5005
R41324 VCC.n15314 VCC.n15313 4.5005
R41325 VCC.n15327 VCC.n15326 4.5005
R41326 VCC.n15326 VCC.n15325 4.5005
R41327 VCC.n15076 VCC.n15072 4.5005
R41328 VCC.n15299 VCC.n15076 4.5005
R41329 VCC.n15290 VCC.n15289 4.5005
R41330 VCC.n15290 VCC.n15083 4.5005
R41331 VCC.n15342 VCC.n15341 4.5005
R41332 VCC.n15343 VCC.n15342 4.5005
R41333 VCC.n15334 VCC.n15055 4.5005
R41334 VCC.n15345 VCC.n15055 4.5005
R41335 VCC.n15349 VCC.n15047 4.5005
R41336 VCC.n15350 VCC.n15349 4.5005
R41337 VCC.n15370 VCC.n15369 4.5005
R41338 VCC.n15371 VCC.n15370 4.5005
R41339 VCC.n15036 VCC.n15034 4.5005
R41340 VCC.n15390 VCC.n15036 4.5005
R41341 VCC.n14976 VCC.n14971 4.5005
R41342 VCC.n15503 VCC.n15502 4.5005
R41343 VCC.n15413 VCC.n15412 4.5005
R41344 VCC.n15019 VCC.n15017 4.5005
R41345 VCC.n15438 VCC.n15437 4.5005
R41346 VCC.n15005 VCC.n15003 4.5005
R41347 VCC.n15003 VCC.n15002 4.5005
R41348 VCC.n15007 VCC.n15006 4.5005
R41349 VCC.n15421 VCC.n15009 4.5005
R41350 VCC.n15426 VCC.n15425 4.5005
R41351 VCC.n15410 VCC.n15409 4.5005
R41352 VCC.n15415 VCC.n15414 4.5005
R41353 VCC.n14978 VCC.n14977 4.5005
R41354 VCC.n15489 VCC.n14978 4.5005
R41355 VCC.n15477 VCC.n15476 4.5005
R41356 VCC.n14988 VCC.n14975 4.5005
R41357 VCC.n15467 VCC.n15466 4.5005
R41358 VCC.n14997 VCC.n14995 4.5005
R41359 VCC.n15468 VCC.n14990 4.5005
R41360 VCC.n15478 VCC.n14986 4.5005
R41361 VCC.n15480 VCC.n15479 4.5005
R41362 VCC.n15480 VCC.n14984 4.5005
R41363 VCC.n15501 VCC.n14970 4.5005
R41364 VCC.n15512 VCC.n15511 4.5005
R41365 VCC.n15012 VCC.n15010 4.5005
R41366 VCC.n15970 VCC.n15572 4.5005
R41367 VCC.n15973 VCC.n15972 4.5005
R41368 VCC.n16047 VCC.n15527 4.5005
R41369 VCC.n16049 VCC.n16048 4.5005
R41370 VCC.n15544 VCC.n15543 4.5005
R41371 VCC.n15564 VCC.n15562 4.5005
R41372 VCC.n15574 VCC.n15561 4.5005
R41373 VCC.n16003 VCC.n16002 4.5005
R41374 VCC.n16012 VCC.n16011 4.5005
R41375 VCC.n15555 VCC.n15554 4.5005
R41376 VCC.n15535 VCC.n15534 4.5005
R41377 VCC.n16038 VCC.n16037 4.5005
R41378 VCC.n16050 VCC.n15525 4.5005
R41379 VCC.n15539 VCC.n15537 4.5005
R41380 VCC.n16010 VCC.n16009 4.5005
R41381 VCC.n15971 VCC.n15969 4.5005
R41382 VCC.n15967 VCC.n15966 4.5005
R41383 VCC.n15982 VCC.n15573 4.5005
R41384 VCC.n16052 VCC.n16051 4.5005
R41385 VCC.n16052 VCC.n15523 4.5005
R41386 VCC.n15542 VCC.n15540 4.5005
R41387 VCC.n15547 VCC.n15540 4.5005
R41388 VCC.n15998 VCC.n15997 4.5005
R41389 VCC.n15999 VCC.n15998 4.5005
R41390 VCC.n16065 VCC.n16064 4.5005
R41391 VCC.n15952 VCC.n15589 4.5005
R41392 VCC.n15951 VCC.n15950 4.5005
R41393 VCC.n15916 VCC.n15601 4.5005
R41394 VCC.n15870 VCC.n15869 4.5005
R41395 VCC.n15844 VCC.n15843 4.5005
R41396 VCC.n15839 VCC.n15835 4.5005
R41397 VCC.n15845 VCC.n15641 4.5005
R41398 VCC.n15641 VCC.n15639 4.5005
R41399 VCC.n15963 VCC.n15962 4.5005
R41400 VCC.n15918 VCC.n15917 4.5005
R41401 VCC.n15838 VCC.n15837 4.5005
R41402 VCC.n15632 VCC.n15628 4.5005
R41403 VCC.n15855 VCC.n15632 4.5005
R41404 VCC.n15868 VCC.n15867 4.5005
R41405 VCC.n15883 VCC.n15882 4.5005
R41406 VCC.n15882 VCC.n15881 4.5005
R41407 VCC.n15898 VCC.n15897 4.5005
R41408 VCC.n15899 VCC.n15898 4.5005
R41409 VCC.n15890 VCC.n15611 4.5005
R41410 VCC.n15901 VCC.n15611 4.5005
R41411 VCC.n15905 VCC.n15603 4.5005
R41412 VCC.n15906 VCC.n15905 4.5005
R41413 VCC.n15926 VCC.n15925 4.5005
R41414 VCC.n15927 VCC.n15926 4.5005
R41415 VCC.n15954 VCC.n15953 4.5005
R41416 VCC.n15592 VCC.n15590 4.5005
R41417 VCC.n15947 VCC.n15592 4.5005
R41418 VCC.n15817 VCC.n15651 4.5005
R41419 VCC.n15816 VCC.n15815 4.5005
R41420 VCC.n15790 VCC.n15662 4.5005
R41421 VCC.n15755 VCC.n15754 4.5005
R41422 VCC.n15720 VCC.n15719 4.5005
R41423 VCC.n15716 VCC.n15713 4.5005
R41424 VCC.n15722 VCC.n15721 4.5005
R41425 VCC.n15723 VCC.n15722 4.5005
R41426 VCC.n15828 VCC.n15827 4.5005
R41427 VCC.n15792 VCC.n15791 4.5005
R41428 VCC.n15715 VCC.n15714 4.5005
R41429 VCC.n15737 VCC.n15690 4.5005
R41430 VCC.n15737 VCC.n15700 4.5005
R41431 VCC.n15752 VCC.n15691 4.5005
R41432 VCC.n15762 VCC.n15761 4.5005
R41433 VCC.n15763 VCC.n15762 4.5005
R41434 VCC.n15767 VCC.n15682 4.5005
R41435 VCC.n15767 VCC.n15671 4.5005
R41436 VCC.n15770 VCC.n15683 4.5005
R41437 VCC.n15778 VCC.n15777 4.5005
R41438 VCC.n15779 VCC.n15778 4.5005
R41439 VCC.n15674 VCC.n15664 4.5005
R41440 VCC.n15675 VCC.n15674 4.5005
R41441 VCC.n15800 VCC.n15799 4.5005
R41442 VCC.n15801 VCC.n15800 4.5005
R41443 VCC.n15819 VCC.n15818 4.5005
R41444 VCC.n15654 VCC.n15652 4.5005
R41445 VCC.n15812 VCC.n15654 4.5005
R41446 VCC.n16367 VCC.n16201 4.5005
R41447 VCC.n16366 VCC.n16365 4.5005
R41448 VCC.n16270 VCC.n16269 4.5005
R41449 VCC.n16266 VCC.n16263 4.5005
R41450 VCC.n16302 VCC.n16241 4.5005
R41451 VCC.n16312 VCC.n16311 4.5005
R41452 VCC.n16313 VCC.n16312 4.5005
R41453 VCC.n16265 VCC.n16264 4.5005
R41454 VCC.n16287 VCC.n16240 4.5005
R41455 VCC.n16287 VCC.n16250 4.5005
R41456 VCC.n16272 VCC.n16271 4.5005
R41457 VCC.n16273 VCC.n16272 4.5005
R41458 VCC.n16317 VCC.n16232 4.5005
R41459 VCC.n16317 VCC.n16221 4.5005
R41460 VCC.n16378 VCC.n16377 4.5005
R41461 VCC.n16342 VCC.n16341 4.5005
R41462 VCC.n16340 VCC.n16212 4.5005
R41463 VCC.n16320 VCC.n16233 4.5005
R41464 VCC.n16328 VCC.n16327 4.5005
R41465 VCC.n16329 VCC.n16328 4.5005
R41466 VCC.n16224 VCC.n16214 4.5005
R41467 VCC.n16225 VCC.n16224 4.5005
R41468 VCC.n16350 VCC.n16349 4.5005
R41469 VCC.n16351 VCC.n16350 4.5005
R41470 VCC.n16369 VCC.n16368 4.5005
R41471 VCC.n16204 VCC.n16202 4.5005
R41472 VCC.n16362 VCC.n16204 4.5005
R41473 VCC.n16305 VCC.n16304 4.5005
R41474 VCC.n16502 VCC.n16140 4.5005
R41475 VCC.n16501 VCC.n16500 4.5005
R41476 VCC.n16395 VCC.n16394 4.5005
R41477 VCC.n16390 VCC.n16387 4.5005
R41478 VCC.n16419 VCC.n16418 4.5005
R41479 VCC.n16389 VCC.n16388 4.5005
R41480 VCC.n16513 VCC.n16512 4.5005
R41481 VCC.n16469 VCC.n16468 4.5005
R41482 VCC.n16467 VCC.n16152 4.5005
R41483 VCC.n16504 VCC.n16503 4.5005
R41484 VCC.n16421 VCC.n16420 4.5005
R41485 VCC.n16434 VCC.n16433 4.5005
R41486 VCC.n16433 VCC.n16432 4.5005
R41487 VCC.n16183 VCC.n16179 4.5005
R41488 VCC.n16406 VCC.n16183 4.5005
R41489 VCC.n16397 VCC.n16396 4.5005
R41490 VCC.n16397 VCC.n16190 4.5005
R41491 VCC.n16449 VCC.n16448 4.5005
R41492 VCC.n16450 VCC.n16449 4.5005
R41493 VCC.n16441 VCC.n16162 4.5005
R41494 VCC.n16452 VCC.n16162 4.5005
R41495 VCC.n16456 VCC.n16154 4.5005
R41496 VCC.n16457 VCC.n16456 4.5005
R41497 VCC.n16477 VCC.n16476 4.5005
R41498 VCC.n16478 VCC.n16477 4.5005
R41499 VCC.n16143 VCC.n16141 4.5005
R41500 VCC.n16497 VCC.n16143 4.5005
R41501 VCC.n16083 VCC.n16078 4.5005
R41502 VCC.n16610 VCC.n16609 4.5005
R41503 VCC.n16520 VCC.n16519 4.5005
R41504 VCC.n16126 VCC.n16124 4.5005
R41505 VCC.n16545 VCC.n16544 4.5005
R41506 VCC.n16112 VCC.n16110 4.5005
R41507 VCC.n16110 VCC.n16109 4.5005
R41508 VCC.n16114 VCC.n16113 4.5005
R41509 VCC.n16528 VCC.n16116 4.5005
R41510 VCC.n16533 VCC.n16532 4.5005
R41511 VCC.n16517 VCC.n16516 4.5005
R41512 VCC.n16522 VCC.n16521 4.5005
R41513 VCC.n16085 VCC.n16084 4.5005
R41514 VCC.n16596 VCC.n16085 4.5005
R41515 VCC.n16584 VCC.n16583 4.5005
R41516 VCC.n16095 VCC.n16082 4.5005
R41517 VCC.n16574 VCC.n16573 4.5005
R41518 VCC.n16104 VCC.n16102 4.5005
R41519 VCC.n16575 VCC.n16097 4.5005
R41520 VCC.n16585 VCC.n16093 4.5005
R41521 VCC.n16587 VCC.n16586 4.5005
R41522 VCC.n16587 VCC.n16091 4.5005
R41523 VCC.n16608 VCC.n16077 4.5005
R41524 VCC.n16619 VCC.n16618 4.5005
R41525 VCC.n16119 VCC.n16117 4.5005
R41526 VCC.n17077 VCC.n16679 4.5005
R41527 VCC.n17080 VCC.n17079 4.5005
R41528 VCC.n17154 VCC.n16634 4.5005
R41529 VCC.n17156 VCC.n17155 4.5005
R41530 VCC.n16651 VCC.n16650 4.5005
R41531 VCC.n16671 VCC.n16669 4.5005
R41532 VCC.n16681 VCC.n16668 4.5005
R41533 VCC.n17110 VCC.n17109 4.5005
R41534 VCC.n17119 VCC.n17118 4.5005
R41535 VCC.n16662 VCC.n16661 4.5005
R41536 VCC.n16642 VCC.n16641 4.5005
R41537 VCC.n17145 VCC.n17144 4.5005
R41538 VCC.n17157 VCC.n16632 4.5005
R41539 VCC.n16646 VCC.n16644 4.5005
R41540 VCC.n17117 VCC.n17116 4.5005
R41541 VCC.n17078 VCC.n17076 4.5005
R41542 VCC.n17074 VCC.n17073 4.5005
R41543 VCC.n17089 VCC.n16680 4.5005
R41544 VCC.n17159 VCC.n17158 4.5005
R41545 VCC.n17159 VCC.n16630 4.5005
R41546 VCC.n16649 VCC.n16647 4.5005
R41547 VCC.n16654 VCC.n16647 4.5005
R41548 VCC.n17105 VCC.n17104 4.5005
R41549 VCC.n17106 VCC.n17105 4.5005
R41550 VCC.n17172 VCC.n17171 4.5005
R41551 VCC.n17059 VCC.n16696 4.5005
R41552 VCC.n17058 VCC.n17057 4.5005
R41553 VCC.n17023 VCC.n16708 4.5005
R41554 VCC.n16977 VCC.n16976 4.5005
R41555 VCC.n16951 VCC.n16950 4.5005
R41556 VCC.n16946 VCC.n16942 4.5005
R41557 VCC.n16952 VCC.n16748 4.5005
R41558 VCC.n16748 VCC.n16746 4.5005
R41559 VCC.n17070 VCC.n17069 4.5005
R41560 VCC.n17025 VCC.n17024 4.5005
R41561 VCC.n16945 VCC.n16944 4.5005
R41562 VCC.n16739 VCC.n16735 4.5005
R41563 VCC.n16962 VCC.n16739 4.5005
R41564 VCC.n16975 VCC.n16974 4.5005
R41565 VCC.n16990 VCC.n16989 4.5005
R41566 VCC.n16989 VCC.n16988 4.5005
R41567 VCC.n17005 VCC.n17004 4.5005
R41568 VCC.n17006 VCC.n17005 4.5005
R41569 VCC.n16997 VCC.n16718 4.5005
R41570 VCC.n17008 VCC.n16718 4.5005
R41571 VCC.n17012 VCC.n16710 4.5005
R41572 VCC.n17013 VCC.n17012 4.5005
R41573 VCC.n17033 VCC.n17032 4.5005
R41574 VCC.n17034 VCC.n17033 4.5005
R41575 VCC.n17061 VCC.n17060 4.5005
R41576 VCC.n16699 VCC.n16697 4.5005
R41577 VCC.n17054 VCC.n16699 4.5005
R41578 VCC.n16924 VCC.n16758 4.5005
R41579 VCC.n16923 VCC.n16922 4.5005
R41580 VCC.n16897 VCC.n16769 4.5005
R41581 VCC.n16862 VCC.n16861 4.5005
R41582 VCC.n16827 VCC.n16826 4.5005
R41583 VCC.n16823 VCC.n16820 4.5005
R41584 VCC.n16829 VCC.n16828 4.5005
R41585 VCC.n16830 VCC.n16829 4.5005
R41586 VCC.n16935 VCC.n16934 4.5005
R41587 VCC.n16899 VCC.n16898 4.5005
R41588 VCC.n16822 VCC.n16821 4.5005
R41589 VCC.n16844 VCC.n16797 4.5005
R41590 VCC.n16844 VCC.n16807 4.5005
R41591 VCC.n16859 VCC.n16798 4.5005
R41592 VCC.n16869 VCC.n16868 4.5005
R41593 VCC.n16870 VCC.n16869 4.5005
R41594 VCC.n16874 VCC.n16789 4.5005
R41595 VCC.n16874 VCC.n16778 4.5005
R41596 VCC.n16877 VCC.n16790 4.5005
R41597 VCC.n16885 VCC.n16884 4.5005
R41598 VCC.n16886 VCC.n16885 4.5005
R41599 VCC.n16781 VCC.n16771 4.5005
R41600 VCC.n16782 VCC.n16781 4.5005
R41601 VCC.n16907 VCC.n16906 4.5005
R41602 VCC.n16908 VCC.n16907 4.5005
R41603 VCC.n16926 VCC.n16925 4.5005
R41604 VCC.n16761 VCC.n16759 4.5005
R41605 VCC.n16919 VCC.n16761 4.5005
R41606 VCC.n17422 VCC.n17247 4.5005
R41607 VCC.n17421 VCC.n17420 4.5005
R41608 VCC.n17315 VCC.n17314 4.5005
R41609 VCC.n17310 VCC.n17307 4.5005
R41610 VCC.n17339 VCC.n17338 4.5005
R41611 VCC.n17309 VCC.n17308 4.5005
R41612 VCC.n17433 VCC.n17432 4.5005
R41613 VCC.n17389 VCC.n17388 4.5005
R41614 VCC.n17387 VCC.n17259 4.5005
R41615 VCC.n17424 VCC.n17423 4.5005
R41616 VCC.n17341 VCC.n17340 4.5005
R41617 VCC.n17354 VCC.n17353 4.5005
R41618 VCC.n17353 VCC.n17352 4.5005
R41619 VCC.n17290 VCC.n17286 4.5005
R41620 VCC.n17326 VCC.n17290 4.5005
R41621 VCC.n17317 VCC.n17316 4.5005
R41622 VCC.n17317 VCC.n17297 4.5005
R41623 VCC.n17369 VCC.n17368 4.5005
R41624 VCC.n17370 VCC.n17369 4.5005
R41625 VCC.n17361 VCC.n17269 4.5005
R41626 VCC.n17372 VCC.n17269 4.5005
R41627 VCC.n17376 VCC.n17261 4.5005
R41628 VCC.n17377 VCC.n17376 4.5005
R41629 VCC.n17397 VCC.n17396 4.5005
R41630 VCC.n17398 VCC.n17397 4.5005
R41631 VCC.n17250 VCC.n17248 4.5005
R41632 VCC.n17417 VCC.n17250 4.5005
R41633 VCC.n17190 VCC.n17185 4.5005
R41634 VCC.n17530 VCC.n17529 4.5005
R41635 VCC.n17440 VCC.n17439 4.5005
R41636 VCC.n17233 VCC.n17231 4.5005
R41637 VCC.n17465 VCC.n17464 4.5005
R41638 VCC.n17219 VCC.n17217 4.5005
R41639 VCC.n17217 VCC.n17216 4.5005
R41640 VCC.n17221 VCC.n17220 4.5005
R41641 VCC.n17448 VCC.n17223 4.5005
R41642 VCC.n17453 VCC.n17452 4.5005
R41643 VCC.n17437 VCC.n17436 4.5005
R41644 VCC.n17442 VCC.n17441 4.5005
R41645 VCC.n17192 VCC.n17191 4.5005
R41646 VCC.n17516 VCC.n17192 4.5005
R41647 VCC.n17504 VCC.n17503 4.5005
R41648 VCC.n17202 VCC.n17189 4.5005
R41649 VCC.n17494 VCC.n17493 4.5005
R41650 VCC.n17211 VCC.n17209 4.5005
R41651 VCC.n17495 VCC.n17204 4.5005
R41652 VCC.n17505 VCC.n17200 4.5005
R41653 VCC.n17507 VCC.n17506 4.5005
R41654 VCC.n17507 VCC.n17198 4.5005
R41655 VCC.n17528 VCC.n17184 4.5005
R41656 VCC.n17539 VCC.n17538 4.5005
R41657 VCC.n17226 VCC.n17224 4.5005
R41658 VCC.n548 VCC.n4 4.31039
R41659 VCC.n1102 VCC.n558 4.31039
R41660 VCC.n1655 VCC.n1111 4.31039
R41661 VCC.n2211 VCC.n1667 4.31039
R41662 VCC.n2764 VCC.n2220 4.31039
R41663 VCC.n3320 VCC.n2776 4.31039
R41664 VCC.n3873 VCC.n3329 4.31039
R41665 VCC.n4429 VCC.n3885 4.31039
R41666 VCC.n4982 VCC.n4438 4.31039
R41667 VCC.n5538 VCC.n4994 4.31039
R41668 VCC.n6091 VCC.n5547 4.31039
R41669 VCC.n6647 VCC.n6103 4.31039
R41670 VCC.n7200 VCC.n6656 4.31039
R41671 VCC.n7756 VCC.n7212 4.31039
R41672 VCC.n8309 VCC.n7765 4.31039
R41673 VCC.n8865 VCC.n8321 4.31039
R41674 VCC.n9418 VCC.n8874 4.31039
R41675 VCC.n9974 VCC.n9430 4.31039
R41676 VCC.n10526 VCC.n9982 4.31039
R41677 VCC.n11081 VCC.n10537 4.31039
R41678 VCC.n11633 VCC.n11089 4.31039
R41679 VCC.n12188 VCC.n11644 4.31039
R41680 VCC.n12740 VCC.n12196 4.31039
R41681 VCC.n13295 VCC.n12751 4.31039
R41682 VCC.n13847 VCC.n13303 4.31039
R41683 VCC.n14402 VCC.n13858 4.31039
R41684 VCC.n14954 VCC.n14410 4.31039
R41685 VCC.n15509 VCC.n14965 4.31039
R41686 VCC.n16061 VCC.n15517 4.31039
R41687 VCC.n16616 VCC.n16072 4.31039
R41688 VCC.n17168 VCC.n16624 4.31039
R41689 VCC.n17536 VCC.n17179 4.31039
R41690 VCC.n472 VCC.n41 3.51902
R41691 VCC.n525 VCC.n22 3.51902
R41692 VCC.n1024 VCC.n593 3.51902
R41693 VCC.n1077 VCC.n574 3.51902
R41694 VCC.n1585 VCC.n1584 3.51902
R41695 VCC.n1621 VCC.n1620 3.51902
R41696 VCC.n2133 VCC.n1702 3.51902
R41697 VCC.n2186 VCC.n1683 3.51902
R41698 VCC.n2694 VCC.n2693 3.51902
R41699 VCC.n2730 VCC.n2729 3.51902
R41700 VCC.n3242 VCC.n2811 3.51902
R41701 VCC.n3295 VCC.n2792 3.51902
R41702 VCC.n3803 VCC.n3802 3.51902
R41703 VCC.n3839 VCC.n3838 3.51902
R41704 VCC.n4351 VCC.n3920 3.51902
R41705 VCC.n4404 VCC.n3901 3.51902
R41706 VCC.n4912 VCC.n4911 3.51902
R41707 VCC.n4948 VCC.n4947 3.51902
R41708 VCC.n5460 VCC.n5029 3.51902
R41709 VCC.n5513 VCC.n5010 3.51902
R41710 VCC.n6021 VCC.n6020 3.51902
R41711 VCC.n6057 VCC.n6056 3.51902
R41712 VCC.n6569 VCC.n6138 3.51902
R41713 VCC.n6622 VCC.n6119 3.51902
R41714 VCC.n7130 VCC.n7129 3.51902
R41715 VCC.n7166 VCC.n7165 3.51902
R41716 VCC.n7678 VCC.n7247 3.51902
R41717 VCC.n7731 VCC.n7228 3.51902
R41718 VCC.n8239 VCC.n8238 3.51902
R41719 VCC.n8275 VCC.n8274 3.51902
R41720 VCC.n8787 VCC.n8356 3.51902
R41721 VCC.n8840 VCC.n8337 3.51902
R41722 VCC.n9348 VCC.n9347 3.51902
R41723 VCC.n9384 VCC.n9383 3.51902
R41724 VCC.n9896 VCC.n9465 3.51902
R41725 VCC.n9949 VCC.n9446 3.51902
R41726 VCC.n10456 VCC.n10455 3.51902
R41727 VCC.n10492 VCC.n10491 3.51902
R41728 VCC.n11003 VCC.n10572 3.51902
R41729 VCC.n11056 VCC.n10553 3.51902
R41730 VCC.n11563 VCC.n11562 3.51902
R41731 VCC.n11599 VCC.n11598 3.51902
R41732 VCC.n12110 VCC.n11679 3.51902
R41733 VCC.n12163 VCC.n11660 3.51902
R41734 VCC.n12670 VCC.n12669 3.51902
R41735 VCC.n12706 VCC.n12705 3.51902
R41736 VCC.n13217 VCC.n12786 3.51902
R41737 VCC.n13270 VCC.n12767 3.51902
R41738 VCC.n13777 VCC.n13776 3.51902
R41739 VCC.n13813 VCC.n13812 3.51902
R41740 VCC.n14324 VCC.n13893 3.51902
R41741 VCC.n14377 VCC.n13874 3.51902
R41742 VCC.n14884 VCC.n14883 3.51902
R41743 VCC.n14920 VCC.n14919 3.51902
R41744 VCC.n15431 VCC.n15000 3.51902
R41745 VCC.n15484 VCC.n14981 3.51902
R41746 VCC.n15991 VCC.n15990 3.51902
R41747 VCC.n16027 VCC.n16026 3.51902
R41748 VCC.n16538 VCC.n16107 3.51902
R41749 VCC.n16591 VCC.n16088 3.51902
R41750 VCC.n17098 VCC.n17097 3.51902
R41751 VCC.n17134 VCC.n17133 3.51902
R41752 VCC.n17458 VCC.n17214 3.51902
R41753 VCC.n17511 VCC.n17195 3.51902
R41754 VCC.n313 VCC.n312 3.42479
R41755 VCC.n315 VCC.n314 3.42479
R41756 VCC.n865 VCC.n864 3.42479
R41757 VCC.n867 VCC.n866 3.42479
R41758 VCC.n1425 VCC.n1424 3.42479
R41759 VCC.n1423 VCC.n1422 3.42479
R41760 VCC.n1974 VCC.n1973 3.42479
R41761 VCC.n1976 VCC.n1975 3.42479
R41762 VCC.n2534 VCC.n2533 3.42479
R41763 VCC.n2532 VCC.n2531 3.42479
R41764 VCC.n3083 VCC.n3082 3.42479
R41765 VCC.n3085 VCC.n3084 3.42479
R41766 VCC.n3643 VCC.n3642 3.42479
R41767 VCC.n3641 VCC.n3640 3.42479
R41768 VCC.n4192 VCC.n4191 3.42479
R41769 VCC.n4194 VCC.n4193 3.42479
R41770 VCC.n4752 VCC.n4751 3.42479
R41771 VCC.n4750 VCC.n4749 3.42479
R41772 VCC.n5301 VCC.n5300 3.42479
R41773 VCC.n5303 VCC.n5302 3.42479
R41774 VCC.n5861 VCC.n5860 3.42479
R41775 VCC.n5859 VCC.n5858 3.42479
R41776 VCC.n6410 VCC.n6409 3.42479
R41777 VCC.n6412 VCC.n6411 3.42479
R41778 VCC.n6970 VCC.n6969 3.42479
R41779 VCC.n6968 VCC.n6967 3.42479
R41780 VCC.n7519 VCC.n7518 3.42479
R41781 VCC.n7521 VCC.n7520 3.42479
R41782 VCC.n8079 VCC.n8078 3.42479
R41783 VCC.n8077 VCC.n8076 3.42479
R41784 VCC.n8630 VCC.n8629 3.42479
R41785 VCC.n8628 VCC.n8627 3.42479
R41786 VCC.n9188 VCC.n9187 3.42479
R41787 VCC.n9186 VCC.n9185 3.42479
R41788 VCC.n9737 VCC.n9736 3.42479
R41789 VCC.n9739 VCC.n9738 3.42479
R41790 VCC.n10296 VCC.n10295 3.42479
R41791 VCC.n10294 VCC.n10293 3.42479
R41792 VCC.n10844 VCC.n10843 3.42479
R41793 VCC.n10846 VCC.n10845 3.42479
R41794 VCC.n11403 VCC.n11402 3.42479
R41795 VCC.n11401 VCC.n11400 3.42479
R41796 VCC.n11951 VCC.n11950 3.42479
R41797 VCC.n11953 VCC.n11952 3.42479
R41798 VCC.n12510 VCC.n12509 3.42479
R41799 VCC.n12508 VCC.n12507 3.42479
R41800 VCC.n13058 VCC.n13057 3.42479
R41801 VCC.n13060 VCC.n13059 3.42479
R41802 VCC.n13617 VCC.n13616 3.42479
R41803 VCC.n13615 VCC.n13614 3.42479
R41804 VCC.n14165 VCC.n14164 3.42479
R41805 VCC.n14167 VCC.n14166 3.42479
R41806 VCC.n14724 VCC.n14723 3.42479
R41807 VCC.n14722 VCC.n14721 3.42479
R41808 VCC.n15272 VCC.n15271 3.42479
R41809 VCC.n15274 VCC.n15273 3.42479
R41810 VCC.n15831 VCC.n15830 3.42479
R41811 VCC.n15829 VCC.n15828 3.42479
R41812 VCC.n16379 VCC.n16378 3.42479
R41813 VCC.n16381 VCC.n16380 3.42479
R41814 VCC.n16938 VCC.n16937 3.42479
R41815 VCC.n16936 VCC.n16935 3.42479
R41816 VCC.n17301 VCC.n17300 3.42479
R41817 VCC.n192 VCC.n191 3.42389
R41818 VCC.n448 VCC.n447 3.42389
R41819 VCC.n450 VCC.n449 3.42389
R41820 VCC.n744 VCC.n743 3.42389
R41821 VCC.n1000 VCC.n999 3.42389
R41822 VCC.n1002 VCC.n1001 3.42389
R41823 VCC.n1560 VCC.n1559 3.42389
R41824 VCC.n1558 VCC.n1557 3.42389
R41825 VCC.n1302 VCC.n1301 3.42389
R41826 VCC.n1853 VCC.n1852 3.42389
R41827 VCC.n2109 VCC.n2108 3.42389
R41828 VCC.n2111 VCC.n2110 3.42389
R41829 VCC.n2669 VCC.n2668 3.42389
R41830 VCC.n2667 VCC.n2666 3.42389
R41831 VCC.n2411 VCC.n2410 3.42389
R41832 VCC.n2962 VCC.n2961 3.42389
R41833 VCC.n3218 VCC.n3217 3.42389
R41834 VCC.n3220 VCC.n3219 3.42389
R41835 VCC.n3778 VCC.n3777 3.42389
R41836 VCC.n3776 VCC.n3775 3.42389
R41837 VCC.n3520 VCC.n3519 3.42389
R41838 VCC.n4071 VCC.n4070 3.42389
R41839 VCC.n4327 VCC.n4326 3.42389
R41840 VCC.n4329 VCC.n4328 3.42389
R41841 VCC.n4887 VCC.n4886 3.42389
R41842 VCC.n4885 VCC.n4884 3.42389
R41843 VCC.n4629 VCC.n4628 3.42389
R41844 VCC.n5180 VCC.n5179 3.42389
R41845 VCC.n5436 VCC.n5435 3.42389
R41846 VCC.n5438 VCC.n5437 3.42389
R41847 VCC.n5996 VCC.n5995 3.42389
R41848 VCC.n5994 VCC.n5993 3.42389
R41849 VCC.n5738 VCC.n5737 3.42389
R41850 VCC.n6289 VCC.n6288 3.42389
R41851 VCC.n6545 VCC.n6544 3.42389
R41852 VCC.n6547 VCC.n6546 3.42389
R41853 VCC.n7105 VCC.n7104 3.42389
R41854 VCC.n7103 VCC.n7102 3.42389
R41855 VCC.n6847 VCC.n6846 3.42389
R41856 VCC.n7398 VCC.n7397 3.42389
R41857 VCC.n7654 VCC.n7653 3.42389
R41858 VCC.n7656 VCC.n7655 3.42389
R41859 VCC.n8214 VCC.n8213 3.42389
R41860 VCC.n8212 VCC.n8211 3.42389
R41861 VCC.n7956 VCC.n7955 3.42389
R41862 VCC.n8763 VCC.n8762 3.42389
R41863 VCC.n8765 VCC.n8764 3.42389
R41864 VCC.n8507 VCC.n8506 3.42389
R41865 VCC.n9323 VCC.n9322 3.42389
R41866 VCC.n9321 VCC.n9320 3.42389
R41867 VCC.n9065 VCC.n9064 3.42389
R41868 VCC.n9616 VCC.n9615 3.42389
R41869 VCC.n9872 VCC.n9871 3.42389
R41870 VCC.n9874 VCC.n9873 3.42389
R41871 VCC.n10431 VCC.n10430 3.42389
R41872 VCC.n10429 VCC.n10428 3.42389
R41873 VCC.n10173 VCC.n10172 3.42389
R41874 VCC.n10723 VCC.n10722 3.42389
R41875 VCC.n10979 VCC.n10978 3.42389
R41876 VCC.n10981 VCC.n10980 3.42389
R41877 VCC.n11538 VCC.n11537 3.42389
R41878 VCC.n11536 VCC.n11535 3.42389
R41879 VCC.n11280 VCC.n11279 3.42389
R41880 VCC.n11830 VCC.n11829 3.42389
R41881 VCC.n12086 VCC.n12085 3.42389
R41882 VCC.n12088 VCC.n12087 3.42389
R41883 VCC.n12645 VCC.n12644 3.42389
R41884 VCC.n12643 VCC.n12642 3.42389
R41885 VCC.n12387 VCC.n12386 3.42389
R41886 VCC.n12937 VCC.n12936 3.42389
R41887 VCC.n13193 VCC.n13192 3.42389
R41888 VCC.n13195 VCC.n13194 3.42389
R41889 VCC.n13752 VCC.n13751 3.42389
R41890 VCC.n13750 VCC.n13749 3.42389
R41891 VCC.n13494 VCC.n13493 3.42389
R41892 VCC.n14044 VCC.n14043 3.42389
R41893 VCC.n14300 VCC.n14299 3.42389
R41894 VCC.n14302 VCC.n14301 3.42389
R41895 VCC.n14859 VCC.n14858 3.42389
R41896 VCC.n14857 VCC.n14856 3.42389
R41897 VCC.n14601 VCC.n14600 3.42389
R41898 VCC.n15151 VCC.n15150 3.42389
R41899 VCC.n15407 VCC.n15406 3.42389
R41900 VCC.n15409 VCC.n15408 3.42389
R41901 VCC.n15966 VCC.n15965 3.42389
R41902 VCC.n15964 VCC.n15963 3.42389
R41903 VCC.n15708 VCC.n15707 3.42389
R41904 VCC.n16258 VCC.n16257 3.42389
R41905 VCC.n16514 VCC.n16513 3.42389
R41906 VCC.n16516 VCC.n16515 3.42389
R41907 VCC.n17073 VCC.n17072 3.42389
R41908 VCC.n17071 VCC.n17070 3.42389
R41909 VCC.n16815 VCC.n16814 3.42389
R41910 VCC.n17434 VCC.n17433 3.42389
R41911 VCC.n17436 VCC.n17435 3.42389
R41912 VCC.n552 VCC.n551 3.423
R41913 VCC.n1106 VCC.n1105 3.423
R41914 VCC.n1660 VCC.n1659 3.423
R41915 VCC.n2215 VCC.n2214 3.423
R41916 VCC.n2769 VCC.n2768 3.423
R41917 VCC.n3324 VCC.n3323 3.423
R41918 VCC.n3878 VCC.n3877 3.423
R41919 VCC.n4433 VCC.n4432 3.423
R41920 VCC.n4987 VCC.n4986 3.423
R41921 VCC.n5542 VCC.n5541 3.423
R41922 VCC.n6096 VCC.n6095 3.423
R41923 VCC.n6651 VCC.n6650 3.423
R41924 VCC.n7205 VCC.n7204 3.423
R41925 VCC.n7760 VCC.n7759 3.423
R41926 VCC.n8314 VCC.n8313 3.423
R41927 VCC.n8869 VCC.n8868 3.423
R41928 VCC.n9423 VCC.n9422 3.423
R41929 VCC.n9978 VCC.n9977 3.423
R41930 VCC.n10531 VCC.n10530 3.423
R41931 VCC.n11085 VCC.n11084 3.423
R41932 VCC.n11638 VCC.n11637 3.423
R41933 VCC.n12192 VCC.n12191 3.423
R41934 VCC.n12745 VCC.n12744 3.423
R41935 VCC.n13299 VCC.n13298 3.423
R41936 VCC.n13852 VCC.n13851 3.423
R41937 VCC.n14406 VCC.n14405 3.423
R41938 VCC.n14959 VCC.n14958 3.423
R41939 VCC.n15513 VCC.n15512 3.423
R41940 VCC.n16066 VCC.n16065 3.423
R41941 VCC.n16620 VCC.n16619 3.423
R41942 VCC.n17173 VCC.n17172 3.423
R41943 VCC.n17540 VCC.n17539 3.423
R41944 VCC.n514 VCC.n513 3.4105
R41945 VCC.n536 VCC.n535 3.4105
R41946 VCC.n535 VCC.n534 3.4105
R41947 VCC.n504 VCC.n33 3.4105
R41948 VCC.n33 VCC.n32 3.4105
R41949 VCC.n506 VCC.n505 3.4105
R41950 VCC.n512 VCC.n511 3.4105
R41951 VCC.n511 VCC.n510 3.4105
R41952 VCC.n486 VCC.n485 3.4105
R41953 VCC.n486 VCC.n45 3.4105
R41954 VCC.n482 VCC.n35 3.4105
R41955 VCC.n503 VCC.n502 3.4105
R41956 VCC.n502 VCC.n501 3.4105
R41957 VCC.n464 VCC.n461 3.4105
R41958 VCC.n464 VCC.n463 3.4105
R41959 VCC.n481 VCC.n480 3.4105
R41960 VCC.n444 VCC.n443 3.4105
R41961 VCC.n445 VCC.n444 3.4105
R41962 VCC.n409 VCC.n408 3.4105
R41963 VCC.n442 VCC.n441 3.4105
R41964 VCC.n441 VCC.n440 3.4105
R41965 VCC.n379 VCC.n378 3.4105
R41966 VCC.n378 VCC.n377 3.4105
R41967 VCC.n374 VCC.n372 3.4105
R41968 VCC.n407 VCC.n406 3.4105
R41969 VCC.n406 VCC.n405 3.4105
R41970 VCC.n103 VCC.n102 3.4105
R41971 VCC.n350 VCC.n103 3.4105
R41972 VCC.n371 VCC.n100 3.4105
R41973 VCC.n381 VCC.n380 3.4105
R41974 VCC.n381 VCC.n99 3.4105
R41975 VCC.n344 VCC.n114 3.4105
R41976 VCC.n344 VCC.n343 3.4105
R41977 VCC.n348 VCC.n347 3.4105
R41978 VCC.n318 VCC.n317 3.4105
R41979 VCC.n318 VCC.n125 3.4105
R41980 VCC.n309 VCC.n308 3.4105
R41981 VCC.n310 VCC.n309 3.4105
R41982 VCC.n282 VCC.n281 3.4105
R41983 VCC.n307 VCC.n306 3.4105
R41984 VCC.n306 VCC.n305 3.4105
R41985 VCC.n258 VCC.n163 3.4105
R41986 VCC.n163 VCC.n157 3.4105
R41987 VCC.n260 VCC.n259 3.4105
R41988 VCC.n280 VCC.n279 3.4105
R41989 VCC.n279 VCC.n278 3.4105
R41990 VCC.n242 VCC.n171 3.4105
R41991 VCC.n171 VCC.n170 3.4105
R41992 VCC.n172 VCC.n165 3.4105
R41993 VCC.n257 VCC.n256 3.4105
R41994 VCC.n256 VCC.n255 3.4105
R41995 VCC.n219 VCC.n218 3.4105
R41996 VCC.n220 VCC.n219 3.4105
R41997 VCC.n241 VCC.n240 3.4105
R41998 VCC.n217 VCC.n216 3.4105
R41999 VCC.n216 VCC.n215 3.4105
R42000 VCC.n460 VCC.n459 3.4105
R42001 VCC.n459 VCC.n458 3.4105
R42002 VCC.n538 VCC.n537 3.4105
R42003 VCC.n538 VCC.n2 3.4105
R42004 VCC.n1090 VCC.n1089 3.4105
R42005 VCC.n1090 VCC.n556 3.4105
R42006 VCC.n1066 VCC.n1065 3.4105
R42007 VCC.n1088 VCC.n1087 3.4105
R42008 VCC.n1087 VCC.n1086 3.4105
R42009 VCC.n1056 VCC.n585 3.4105
R42010 VCC.n585 VCC.n584 3.4105
R42011 VCC.n1058 VCC.n1057 3.4105
R42012 VCC.n1064 VCC.n1063 3.4105
R42013 VCC.n1063 VCC.n1062 3.4105
R42014 VCC.n1038 VCC.n1037 3.4105
R42015 VCC.n1038 VCC.n597 3.4105
R42016 VCC.n1034 VCC.n587 3.4105
R42017 VCC.n1055 VCC.n1054 3.4105
R42018 VCC.n1054 VCC.n1053 3.4105
R42019 VCC.n1016 VCC.n1013 3.4105
R42020 VCC.n1016 VCC.n1015 3.4105
R42021 VCC.n1033 VCC.n1032 3.4105
R42022 VCC.n1012 VCC.n1011 3.4105
R42023 VCC.n1011 VCC.n1010 3.4105
R42024 VCC.n996 VCC.n995 3.4105
R42025 VCC.n997 VCC.n996 3.4105
R42026 VCC.n961 VCC.n960 3.4105
R42027 VCC.n994 VCC.n993 3.4105
R42028 VCC.n993 VCC.n992 3.4105
R42029 VCC.n931 VCC.n930 3.4105
R42030 VCC.n930 VCC.n929 3.4105
R42031 VCC.n926 VCC.n924 3.4105
R42032 VCC.n959 VCC.n958 3.4105
R42033 VCC.n958 VCC.n957 3.4105
R42034 VCC.n655 VCC.n654 3.4105
R42035 VCC.n902 VCC.n655 3.4105
R42036 VCC.n923 VCC.n652 3.4105
R42037 VCC.n933 VCC.n932 3.4105
R42038 VCC.n933 VCC.n651 3.4105
R42039 VCC.n896 VCC.n666 3.4105
R42040 VCC.n896 VCC.n895 3.4105
R42041 VCC.n900 VCC.n899 3.4105
R42042 VCC.n870 VCC.n869 3.4105
R42043 VCC.n870 VCC.n677 3.4105
R42044 VCC.n861 VCC.n860 3.4105
R42045 VCC.n862 VCC.n861 3.4105
R42046 VCC.n834 VCC.n833 3.4105
R42047 VCC.n859 VCC.n858 3.4105
R42048 VCC.n858 VCC.n857 3.4105
R42049 VCC.n810 VCC.n715 3.4105
R42050 VCC.n715 VCC.n709 3.4105
R42051 VCC.n812 VCC.n811 3.4105
R42052 VCC.n832 VCC.n831 3.4105
R42053 VCC.n831 VCC.n830 3.4105
R42054 VCC.n794 VCC.n723 3.4105
R42055 VCC.n723 VCC.n722 3.4105
R42056 VCC.n724 VCC.n717 3.4105
R42057 VCC.n809 VCC.n808 3.4105
R42058 VCC.n808 VCC.n807 3.4105
R42059 VCC.n771 VCC.n770 3.4105
R42060 VCC.n772 VCC.n771 3.4105
R42061 VCC.n793 VCC.n792 3.4105
R42062 VCC.n769 VCC.n768 3.4105
R42063 VCC.n768 VCC.n767 3.4105
R42064 VCC.n1419 VCC.n1418 3.4105
R42065 VCC.n1420 VCC.n1419 3.4105
R42066 VCC.n1392 VCC.n1391 3.4105
R42067 VCC.n1417 VCC.n1416 3.4105
R42068 VCC.n1416 VCC.n1415 3.4105
R42069 VCC.n1368 VCC.n1273 3.4105
R42070 VCC.n1273 VCC.n1267 3.4105
R42071 VCC.n1370 VCC.n1369 3.4105
R42072 VCC.n1390 VCC.n1389 3.4105
R42073 VCC.n1389 VCC.n1388 3.4105
R42074 VCC.n1352 VCC.n1281 3.4105
R42075 VCC.n1281 VCC.n1280 3.4105
R42076 VCC.n1282 VCC.n1275 3.4105
R42077 VCC.n1367 VCC.n1366 3.4105
R42078 VCC.n1366 VCC.n1365 3.4105
R42079 VCC.n1329 VCC.n1328 3.4105
R42080 VCC.n1330 VCC.n1329 3.4105
R42081 VCC.n1351 VCC.n1350 3.4105
R42082 VCC.n1327 VCC.n1326 3.4105
R42083 VCC.n1326 VCC.n1325 3.4105
R42084 VCC.n1571 VCC.n1570 3.4105
R42085 VCC.n1570 VCC.n1569 3.4105
R42086 VCC.n1630 VCC.n1629 3.4105
R42087 VCC.n1635 VCC.n1634 3.4105
R42088 VCC.n1634 VCC.n1633 3.4105
R42089 VCC.n1613 VCC.n1612 3.4105
R42090 VCC.n1614 VCC.n1613 3.4105
R42091 VCC.n1611 VCC.n1610 3.4105
R42092 VCC.n1628 VCC.n1627 3.4105
R42093 VCC.n1627 VCC.n1626 3.4105
R42094 VCC.n1600 VCC.n1153 3.4105
R42095 VCC.n1153 VCC.n1152 3.4105
R42096 VCC.n1151 VCC.n1150 3.4105
R42097 VCC.n1608 VCC.n1607 3.4105
R42098 VCC.n1607 VCC.n1146 3.4105
R42099 VCC.n1573 VCC.n1572 3.4105
R42100 VCC.n1573 VCC.n1169 3.4105
R42101 VCC.n1599 VCC.n1598 3.4105
R42102 VCC.n1637 VCC.n1636 3.4105
R42103 VCC.n1637 VCC.n1110 3.4105
R42104 VCC.n1554 VCC.n1553 3.4105
R42105 VCC.n1555 VCC.n1554 3.4105
R42106 VCC.n1518 VCC.n1517 3.4105
R42107 VCC.n1552 VCC.n1551 3.4105
R42108 VCC.n1551 VCC.n1550 3.4105
R42109 VCC.n1488 VCC.n1487 3.4105
R42110 VCC.n1487 VCC.n1486 3.4105
R42111 VCC.n1483 VCC.n1481 3.4105
R42112 VCC.n1516 VCC.n1515 3.4105
R42113 VCC.n1515 VCC.n1514 3.4105
R42114 VCC.n1212 VCC.n1211 3.4105
R42115 VCC.n1459 VCC.n1212 3.4105
R42116 VCC.n1480 VCC.n1209 3.4105
R42117 VCC.n1490 VCC.n1489 3.4105
R42118 VCC.n1490 VCC.n1208 3.4105
R42119 VCC.n1453 VCC.n1223 3.4105
R42120 VCC.n1453 VCC.n1452 3.4105
R42121 VCC.n1457 VCC.n1456 3.4105
R42122 VCC.n1428 VCC.n1427 3.4105
R42123 VCC.n1428 VCC.n1234 3.4105
R42124 VCC.n2199 VCC.n2198 3.4105
R42125 VCC.n2199 VCC.n1665 3.4105
R42126 VCC.n2175 VCC.n2174 3.4105
R42127 VCC.n2197 VCC.n2196 3.4105
R42128 VCC.n2196 VCC.n2195 3.4105
R42129 VCC.n2165 VCC.n1694 3.4105
R42130 VCC.n1694 VCC.n1693 3.4105
R42131 VCC.n2167 VCC.n2166 3.4105
R42132 VCC.n2173 VCC.n2172 3.4105
R42133 VCC.n2172 VCC.n2171 3.4105
R42134 VCC.n2147 VCC.n2146 3.4105
R42135 VCC.n2147 VCC.n1706 3.4105
R42136 VCC.n2143 VCC.n1696 3.4105
R42137 VCC.n2164 VCC.n2163 3.4105
R42138 VCC.n2163 VCC.n2162 3.4105
R42139 VCC.n2125 VCC.n2122 3.4105
R42140 VCC.n2125 VCC.n2124 3.4105
R42141 VCC.n2142 VCC.n2141 3.4105
R42142 VCC.n2121 VCC.n2120 3.4105
R42143 VCC.n2120 VCC.n2119 3.4105
R42144 VCC.n2105 VCC.n2104 3.4105
R42145 VCC.n2106 VCC.n2105 3.4105
R42146 VCC.n2070 VCC.n2069 3.4105
R42147 VCC.n2103 VCC.n2102 3.4105
R42148 VCC.n2102 VCC.n2101 3.4105
R42149 VCC.n2040 VCC.n2039 3.4105
R42150 VCC.n2039 VCC.n2038 3.4105
R42151 VCC.n2035 VCC.n2033 3.4105
R42152 VCC.n2068 VCC.n2067 3.4105
R42153 VCC.n2067 VCC.n2066 3.4105
R42154 VCC.n1764 VCC.n1763 3.4105
R42155 VCC.n2011 VCC.n1764 3.4105
R42156 VCC.n2032 VCC.n1761 3.4105
R42157 VCC.n2042 VCC.n2041 3.4105
R42158 VCC.n2042 VCC.n1760 3.4105
R42159 VCC.n2005 VCC.n1775 3.4105
R42160 VCC.n2005 VCC.n2004 3.4105
R42161 VCC.n2009 VCC.n2008 3.4105
R42162 VCC.n1979 VCC.n1978 3.4105
R42163 VCC.n1979 VCC.n1786 3.4105
R42164 VCC.n1970 VCC.n1969 3.4105
R42165 VCC.n1971 VCC.n1970 3.4105
R42166 VCC.n1943 VCC.n1942 3.4105
R42167 VCC.n1968 VCC.n1967 3.4105
R42168 VCC.n1967 VCC.n1966 3.4105
R42169 VCC.n1919 VCC.n1824 3.4105
R42170 VCC.n1824 VCC.n1818 3.4105
R42171 VCC.n1921 VCC.n1920 3.4105
R42172 VCC.n1941 VCC.n1940 3.4105
R42173 VCC.n1940 VCC.n1939 3.4105
R42174 VCC.n1903 VCC.n1832 3.4105
R42175 VCC.n1832 VCC.n1831 3.4105
R42176 VCC.n1833 VCC.n1826 3.4105
R42177 VCC.n1918 VCC.n1917 3.4105
R42178 VCC.n1917 VCC.n1916 3.4105
R42179 VCC.n1880 VCC.n1879 3.4105
R42180 VCC.n1881 VCC.n1880 3.4105
R42181 VCC.n1902 VCC.n1901 3.4105
R42182 VCC.n1878 VCC.n1877 3.4105
R42183 VCC.n1877 VCC.n1876 3.4105
R42184 VCC.n2528 VCC.n2527 3.4105
R42185 VCC.n2529 VCC.n2528 3.4105
R42186 VCC.n2501 VCC.n2500 3.4105
R42187 VCC.n2526 VCC.n2525 3.4105
R42188 VCC.n2525 VCC.n2524 3.4105
R42189 VCC.n2477 VCC.n2382 3.4105
R42190 VCC.n2382 VCC.n2376 3.4105
R42191 VCC.n2479 VCC.n2478 3.4105
R42192 VCC.n2499 VCC.n2498 3.4105
R42193 VCC.n2498 VCC.n2497 3.4105
R42194 VCC.n2461 VCC.n2390 3.4105
R42195 VCC.n2390 VCC.n2389 3.4105
R42196 VCC.n2391 VCC.n2384 3.4105
R42197 VCC.n2476 VCC.n2475 3.4105
R42198 VCC.n2475 VCC.n2474 3.4105
R42199 VCC.n2438 VCC.n2437 3.4105
R42200 VCC.n2439 VCC.n2438 3.4105
R42201 VCC.n2460 VCC.n2459 3.4105
R42202 VCC.n2436 VCC.n2435 3.4105
R42203 VCC.n2435 VCC.n2434 3.4105
R42204 VCC.n2680 VCC.n2679 3.4105
R42205 VCC.n2679 VCC.n2678 3.4105
R42206 VCC.n2739 VCC.n2738 3.4105
R42207 VCC.n2744 VCC.n2743 3.4105
R42208 VCC.n2743 VCC.n2742 3.4105
R42209 VCC.n2722 VCC.n2721 3.4105
R42210 VCC.n2723 VCC.n2722 3.4105
R42211 VCC.n2720 VCC.n2719 3.4105
R42212 VCC.n2737 VCC.n2736 3.4105
R42213 VCC.n2736 VCC.n2735 3.4105
R42214 VCC.n2709 VCC.n2262 3.4105
R42215 VCC.n2262 VCC.n2261 3.4105
R42216 VCC.n2260 VCC.n2259 3.4105
R42217 VCC.n2717 VCC.n2716 3.4105
R42218 VCC.n2716 VCC.n2255 3.4105
R42219 VCC.n2682 VCC.n2681 3.4105
R42220 VCC.n2682 VCC.n2278 3.4105
R42221 VCC.n2708 VCC.n2707 3.4105
R42222 VCC.n2746 VCC.n2745 3.4105
R42223 VCC.n2746 VCC.n2219 3.4105
R42224 VCC.n2663 VCC.n2662 3.4105
R42225 VCC.n2664 VCC.n2663 3.4105
R42226 VCC.n2627 VCC.n2626 3.4105
R42227 VCC.n2661 VCC.n2660 3.4105
R42228 VCC.n2660 VCC.n2659 3.4105
R42229 VCC.n2597 VCC.n2596 3.4105
R42230 VCC.n2596 VCC.n2595 3.4105
R42231 VCC.n2592 VCC.n2590 3.4105
R42232 VCC.n2625 VCC.n2624 3.4105
R42233 VCC.n2624 VCC.n2623 3.4105
R42234 VCC.n2321 VCC.n2320 3.4105
R42235 VCC.n2568 VCC.n2321 3.4105
R42236 VCC.n2589 VCC.n2318 3.4105
R42237 VCC.n2599 VCC.n2598 3.4105
R42238 VCC.n2599 VCC.n2317 3.4105
R42239 VCC.n2562 VCC.n2332 3.4105
R42240 VCC.n2562 VCC.n2561 3.4105
R42241 VCC.n2566 VCC.n2565 3.4105
R42242 VCC.n2537 VCC.n2536 3.4105
R42243 VCC.n2537 VCC.n2343 3.4105
R42244 VCC.n3308 VCC.n3307 3.4105
R42245 VCC.n3308 VCC.n2774 3.4105
R42246 VCC.n3284 VCC.n3283 3.4105
R42247 VCC.n3306 VCC.n3305 3.4105
R42248 VCC.n3305 VCC.n3304 3.4105
R42249 VCC.n3274 VCC.n2803 3.4105
R42250 VCC.n2803 VCC.n2802 3.4105
R42251 VCC.n3276 VCC.n3275 3.4105
R42252 VCC.n3282 VCC.n3281 3.4105
R42253 VCC.n3281 VCC.n3280 3.4105
R42254 VCC.n3256 VCC.n3255 3.4105
R42255 VCC.n3256 VCC.n2815 3.4105
R42256 VCC.n3252 VCC.n2805 3.4105
R42257 VCC.n3273 VCC.n3272 3.4105
R42258 VCC.n3272 VCC.n3271 3.4105
R42259 VCC.n3234 VCC.n3231 3.4105
R42260 VCC.n3234 VCC.n3233 3.4105
R42261 VCC.n3251 VCC.n3250 3.4105
R42262 VCC.n3230 VCC.n3229 3.4105
R42263 VCC.n3229 VCC.n3228 3.4105
R42264 VCC.n3214 VCC.n3213 3.4105
R42265 VCC.n3215 VCC.n3214 3.4105
R42266 VCC.n3179 VCC.n3178 3.4105
R42267 VCC.n3212 VCC.n3211 3.4105
R42268 VCC.n3211 VCC.n3210 3.4105
R42269 VCC.n3149 VCC.n3148 3.4105
R42270 VCC.n3148 VCC.n3147 3.4105
R42271 VCC.n3144 VCC.n3142 3.4105
R42272 VCC.n3177 VCC.n3176 3.4105
R42273 VCC.n3176 VCC.n3175 3.4105
R42274 VCC.n2873 VCC.n2872 3.4105
R42275 VCC.n3120 VCC.n2873 3.4105
R42276 VCC.n3141 VCC.n2870 3.4105
R42277 VCC.n3151 VCC.n3150 3.4105
R42278 VCC.n3151 VCC.n2869 3.4105
R42279 VCC.n3114 VCC.n2884 3.4105
R42280 VCC.n3114 VCC.n3113 3.4105
R42281 VCC.n3118 VCC.n3117 3.4105
R42282 VCC.n3088 VCC.n3087 3.4105
R42283 VCC.n3088 VCC.n2895 3.4105
R42284 VCC.n3079 VCC.n3078 3.4105
R42285 VCC.n3080 VCC.n3079 3.4105
R42286 VCC.n3052 VCC.n3051 3.4105
R42287 VCC.n3077 VCC.n3076 3.4105
R42288 VCC.n3076 VCC.n3075 3.4105
R42289 VCC.n3028 VCC.n2933 3.4105
R42290 VCC.n2933 VCC.n2927 3.4105
R42291 VCC.n3030 VCC.n3029 3.4105
R42292 VCC.n3050 VCC.n3049 3.4105
R42293 VCC.n3049 VCC.n3048 3.4105
R42294 VCC.n3012 VCC.n2941 3.4105
R42295 VCC.n2941 VCC.n2940 3.4105
R42296 VCC.n2942 VCC.n2935 3.4105
R42297 VCC.n3027 VCC.n3026 3.4105
R42298 VCC.n3026 VCC.n3025 3.4105
R42299 VCC.n2989 VCC.n2988 3.4105
R42300 VCC.n2990 VCC.n2989 3.4105
R42301 VCC.n3011 VCC.n3010 3.4105
R42302 VCC.n2987 VCC.n2986 3.4105
R42303 VCC.n2986 VCC.n2985 3.4105
R42304 VCC.n3637 VCC.n3636 3.4105
R42305 VCC.n3638 VCC.n3637 3.4105
R42306 VCC.n3610 VCC.n3609 3.4105
R42307 VCC.n3635 VCC.n3634 3.4105
R42308 VCC.n3634 VCC.n3633 3.4105
R42309 VCC.n3586 VCC.n3491 3.4105
R42310 VCC.n3491 VCC.n3485 3.4105
R42311 VCC.n3588 VCC.n3587 3.4105
R42312 VCC.n3608 VCC.n3607 3.4105
R42313 VCC.n3607 VCC.n3606 3.4105
R42314 VCC.n3570 VCC.n3499 3.4105
R42315 VCC.n3499 VCC.n3498 3.4105
R42316 VCC.n3500 VCC.n3493 3.4105
R42317 VCC.n3585 VCC.n3584 3.4105
R42318 VCC.n3584 VCC.n3583 3.4105
R42319 VCC.n3547 VCC.n3546 3.4105
R42320 VCC.n3548 VCC.n3547 3.4105
R42321 VCC.n3569 VCC.n3568 3.4105
R42322 VCC.n3545 VCC.n3544 3.4105
R42323 VCC.n3544 VCC.n3543 3.4105
R42324 VCC.n3789 VCC.n3788 3.4105
R42325 VCC.n3788 VCC.n3787 3.4105
R42326 VCC.n3848 VCC.n3847 3.4105
R42327 VCC.n3853 VCC.n3852 3.4105
R42328 VCC.n3852 VCC.n3851 3.4105
R42329 VCC.n3831 VCC.n3830 3.4105
R42330 VCC.n3832 VCC.n3831 3.4105
R42331 VCC.n3829 VCC.n3828 3.4105
R42332 VCC.n3846 VCC.n3845 3.4105
R42333 VCC.n3845 VCC.n3844 3.4105
R42334 VCC.n3818 VCC.n3371 3.4105
R42335 VCC.n3371 VCC.n3370 3.4105
R42336 VCC.n3369 VCC.n3368 3.4105
R42337 VCC.n3826 VCC.n3825 3.4105
R42338 VCC.n3825 VCC.n3364 3.4105
R42339 VCC.n3791 VCC.n3790 3.4105
R42340 VCC.n3791 VCC.n3387 3.4105
R42341 VCC.n3817 VCC.n3816 3.4105
R42342 VCC.n3855 VCC.n3854 3.4105
R42343 VCC.n3855 VCC.n3328 3.4105
R42344 VCC.n3772 VCC.n3771 3.4105
R42345 VCC.n3773 VCC.n3772 3.4105
R42346 VCC.n3736 VCC.n3735 3.4105
R42347 VCC.n3770 VCC.n3769 3.4105
R42348 VCC.n3769 VCC.n3768 3.4105
R42349 VCC.n3706 VCC.n3705 3.4105
R42350 VCC.n3705 VCC.n3704 3.4105
R42351 VCC.n3701 VCC.n3699 3.4105
R42352 VCC.n3734 VCC.n3733 3.4105
R42353 VCC.n3733 VCC.n3732 3.4105
R42354 VCC.n3430 VCC.n3429 3.4105
R42355 VCC.n3677 VCC.n3430 3.4105
R42356 VCC.n3698 VCC.n3427 3.4105
R42357 VCC.n3708 VCC.n3707 3.4105
R42358 VCC.n3708 VCC.n3426 3.4105
R42359 VCC.n3671 VCC.n3441 3.4105
R42360 VCC.n3671 VCC.n3670 3.4105
R42361 VCC.n3675 VCC.n3674 3.4105
R42362 VCC.n3646 VCC.n3645 3.4105
R42363 VCC.n3646 VCC.n3452 3.4105
R42364 VCC.n4417 VCC.n4416 3.4105
R42365 VCC.n4417 VCC.n3883 3.4105
R42366 VCC.n4393 VCC.n4392 3.4105
R42367 VCC.n4415 VCC.n4414 3.4105
R42368 VCC.n4414 VCC.n4413 3.4105
R42369 VCC.n4383 VCC.n3912 3.4105
R42370 VCC.n3912 VCC.n3911 3.4105
R42371 VCC.n4385 VCC.n4384 3.4105
R42372 VCC.n4391 VCC.n4390 3.4105
R42373 VCC.n4390 VCC.n4389 3.4105
R42374 VCC.n4365 VCC.n4364 3.4105
R42375 VCC.n4365 VCC.n3924 3.4105
R42376 VCC.n4361 VCC.n3914 3.4105
R42377 VCC.n4382 VCC.n4381 3.4105
R42378 VCC.n4381 VCC.n4380 3.4105
R42379 VCC.n4343 VCC.n4340 3.4105
R42380 VCC.n4343 VCC.n4342 3.4105
R42381 VCC.n4360 VCC.n4359 3.4105
R42382 VCC.n4339 VCC.n4338 3.4105
R42383 VCC.n4338 VCC.n4337 3.4105
R42384 VCC.n4323 VCC.n4322 3.4105
R42385 VCC.n4324 VCC.n4323 3.4105
R42386 VCC.n4288 VCC.n4287 3.4105
R42387 VCC.n4321 VCC.n4320 3.4105
R42388 VCC.n4320 VCC.n4319 3.4105
R42389 VCC.n4258 VCC.n4257 3.4105
R42390 VCC.n4257 VCC.n4256 3.4105
R42391 VCC.n4253 VCC.n4251 3.4105
R42392 VCC.n4286 VCC.n4285 3.4105
R42393 VCC.n4285 VCC.n4284 3.4105
R42394 VCC.n3982 VCC.n3981 3.4105
R42395 VCC.n4229 VCC.n3982 3.4105
R42396 VCC.n4250 VCC.n3979 3.4105
R42397 VCC.n4260 VCC.n4259 3.4105
R42398 VCC.n4260 VCC.n3978 3.4105
R42399 VCC.n4223 VCC.n3993 3.4105
R42400 VCC.n4223 VCC.n4222 3.4105
R42401 VCC.n4227 VCC.n4226 3.4105
R42402 VCC.n4197 VCC.n4196 3.4105
R42403 VCC.n4197 VCC.n4004 3.4105
R42404 VCC.n4188 VCC.n4187 3.4105
R42405 VCC.n4189 VCC.n4188 3.4105
R42406 VCC.n4161 VCC.n4160 3.4105
R42407 VCC.n4186 VCC.n4185 3.4105
R42408 VCC.n4185 VCC.n4184 3.4105
R42409 VCC.n4137 VCC.n4042 3.4105
R42410 VCC.n4042 VCC.n4036 3.4105
R42411 VCC.n4139 VCC.n4138 3.4105
R42412 VCC.n4159 VCC.n4158 3.4105
R42413 VCC.n4158 VCC.n4157 3.4105
R42414 VCC.n4121 VCC.n4050 3.4105
R42415 VCC.n4050 VCC.n4049 3.4105
R42416 VCC.n4051 VCC.n4044 3.4105
R42417 VCC.n4136 VCC.n4135 3.4105
R42418 VCC.n4135 VCC.n4134 3.4105
R42419 VCC.n4098 VCC.n4097 3.4105
R42420 VCC.n4099 VCC.n4098 3.4105
R42421 VCC.n4120 VCC.n4119 3.4105
R42422 VCC.n4096 VCC.n4095 3.4105
R42423 VCC.n4095 VCC.n4094 3.4105
R42424 VCC.n4746 VCC.n4745 3.4105
R42425 VCC.n4747 VCC.n4746 3.4105
R42426 VCC.n4719 VCC.n4718 3.4105
R42427 VCC.n4744 VCC.n4743 3.4105
R42428 VCC.n4743 VCC.n4742 3.4105
R42429 VCC.n4695 VCC.n4600 3.4105
R42430 VCC.n4600 VCC.n4594 3.4105
R42431 VCC.n4697 VCC.n4696 3.4105
R42432 VCC.n4717 VCC.n4716 3.4105
R42433 VCC.n4716 VCC.n4715 3.4105
R42434 VCC.n4679 VCC.n4608 3.4105
R42435 VCC.n4608 VCC.n4607 3.4105
R42436 VCC.n4609 VCC.n4602 3.4105
R42437 VCC.n4694 VCC.n4693 3.4105
R42438 VCC.n4693 VCC.n4692 3.4105
R42439 VCC.n4656 VCC.n4655 3.4105
R42440 VCC.n4657 VCC.n4656 3.4105
R42441 VCC.n4678 VCC.n4677 3.4105
R42442 VCC.n4654 VCC.n4653 3.4105
R42443 VCC.n4653 VCC.n4652 3.4105
R42444 VCC.n4898 VCC.n4897 3.4105
R42445 VCC.n4897 VCC.n4896 3.4105
R42446 VCC.n4957 VCC.n4956 3.4105
R42447 VCC.n4962 VCC.n4961 3.4105
R42448 VCC.n4961 VCC.n4960 3.4105
R42449 VCC.n4940 VCC.n4939 3.4105
R42450 VCC.n4941 VCC.n4940 3.4105
R42451 VCC.n4938 VCC.n4937 3.4105
R42452 VCC.n4955 VCC.n4954 3.4105
R42453 VCC.n4954 VCC.n4953 3.4105
R42454 VCC.n4927 VCC.n4480 3.4105
R42455 VCC.n4480 VCC.n4479 3.4105
R42456 VCC.n4478 VCC.n4477 3.4105
R42457 VCC.n4935 VCC.n4934 3.4105
R42458 VCC.n4934 VCC.n4473 3.4105
R42459 VCC.n4900 VCC.n4899 3.4105
R42460 VCC.n4900 VCC.n4496 3.4105
R42461 VCC.n4926 VCC.n4925 3.4105
R42462 VCC.n4964 VCC.n4963 3.4105
R42463 VCC.n4964 VCC.n4437 3.4105
R42464 VCC.n4881 VCC.n4880 3.4105
R42465 VCC.n4882 VCC.n4881 3.4105
R42466 VCC.n4845 VCC.n4844 3.4105
R42467 VCC.n4879 VCC.n4878 3.4105
R42468 VCC.n4878 VCC.n4877 3.4105
R42469 VCC.n4815 VCC.n4814 3.4105
R42470 VCC.n4814 VCC.n4813 3.4105
R42471 VCC.n4810 VCC.n4808 3.4105
R42472 VCC.n4843 VCC.n4842 3.4105
R42473 VCC.n4842 VCC.n4841 3.4105
R42474 VCC.n4539 VCC.n4538 3.4105
R42475 VCC.n4786 VCC.n4539 3.4105
R42476 VCC.n4807 VCC.n4536 3.4105
R42477 VCC.n4817 VCC.n4816 3.4105
R42478 VCC.n4817 VCC.n4535 3.4105
R42479 VCC.n4780 VCC.n4550 3.4105
R42480 VCC.n4780 VCC.n4779 3.4105
R42481 VCC.n4784 VCC.n4783 3.4105
R42482 VCC.n4755 VCC.n4754 3.4105
R42483 VCC.n4755 VCC.n4561 3.4105
R42484 VCC.n5526 VCC.n5525 3.4105
R42485 VCC.n5526 VCC.n4992 3.4105
R42486 VCC.n5502 VCC.n5501 3.4105
R42487 VCC.n5524 VCC.n5523 3.4105
R42488 VCC.n5523 VCC.n5522 3.4105
R42489 VCC.n5492 VCC.n5021 3.4105
R42490 VCC.n5021 VCC.n5020 3.4105
R42491 VCC.n5494 VCC.n5493 3.4105
R42492 VCC.n5500 VCC.n5499 3.4105
R42493 VCC.n5499 VCC.n5498 3.4105
R42494 VCC.n5474 VCC.n5473 3.4105
R42495 VCC.n5474 VCC.n5033 3.4105
R42496 VCC.n5470 VCC.n5023 3.4105
R42497 VCC.n5491 VCC.n5490 3.4105
R42498 VCC.n5490 VCC.n5489 3.4105
R42499 VCC.n5452 VCC.n5449 3.4105
R42500 VCC.n5452 VCC.n5451 3.4105
R42501 VCC.n5469 VCC.n5468 3.4105
R42502 VCC.n5448 VCC.n5447 3.4105
R42503 VCC.n5447 VCC.n5446 3.4105
R42504 VCC.n5432 VCC.n5431 3.4105
R42505 VCC.n5433 VCC.n5432 3.4105
R42506 VCC.n5397 VCC.n5396 3.4105
R42507 VCC.n5430 VCC.n5429 3.4105
R42508 VCC.n5429 VCC.n5428 3.4105
R42509 VCC.n5367 VCC.n5366 3.4105
R42510 VCC.n5366 VCC.n5365 3.4105
R42511 VCC.n5362 VCC.n5360 3.4105
R42512 VCC.n5395 VCC.n5394 3.4105
R42513 VCC.n5394 VCC.n5393 3.4105
R42514 VCC.n5091 VCC.n5090 3.4105
R42515 VCC.n5338 VCC.n5091 3.4105
R42516 VCC.n5359 VCC.n5088 3.4105
R42517 VCC.n5369 VCC.n5368 3.4105
R42518 VCC.n5369 VCC.n5087 3.4105
R42519 VCC.n5332 VCC.n5102 3.4105
R42520 VCC.n5332 VCC.n5331 3.4105
R42521 VCC.n5336 VCC.n5335 3.4105
R42522 VCC.n5306 VCC.n5305 3.4105
R42523 VCC.n5306 VCC.n5113 3.4105
R42524 VCC.n5297 VCC.n5296 3.4105
R42525 VCC.n5298 VCC.n5297 3.4105
R42526 VCC.n5270 VCC.n5269 3.4105
R42527 VCC.n5295 VCC.n5294 3.4105
R42528 VCC.n5294 VCC.n5293 3.4105
R42529 VCC.n5246 VCC.n5151 3.4105
R42530 VCC.n5151 VCC.n5145 3.4105
R42531 VCC.n5248 VCC.n5247 3.4105
R42532 VCC.n5268 VCC.n5267 3.4105
R42533 VCC.n5267 VCC.n5266 3.4105
R42534 VCC.n5230 VCC.n5159 3.4105
R42535 VCC.n5159 VCC.n5158 3.4105
R42536 VCC.n5160 VCC.n5153 3.4105
R42537 VCC.n5245 VCC.n5244 3.4105
R42538 VCC.n5244 VCC.n5243 3.4105
R42539 VCC.n5207 VCC.n5206 3.4105
R42540 VCC.n5208 VCC.n5207 3.4105
R42541 VCC.n5229 VCC.n5228 3.4105
R42542 VCC.n5205 VCC.n5204 3.4105
R42543 VCC.n5204 VCC.n5203 3.4105
R42544 VCC.n5855 VCC.n5854 3.4105
R42545 VCC.n5856 VCC.n5855 3.4105
R42546 VCC.n5828 VCC.n5827 3.4105
R42547 VCC.n5853 VCC.n5852 3.4105
R42548 VCC.n5852 VCC.n5851 3.4105
R42549 VCC.n5804 VCC.n5709 3.4105
R42550 VCC.n5709 VCC.n5703 3.4105
R42551 VCC.n5806 VCC.n5805 3.4105
R42552 VCC.n5826 VCC.n5825 3.4105
R42553 VCC.n5825 VCC.n5824 3.4105
R42554 VCC.n5788 VCC.n5717 3.4105
R42555 VCC.n5717 VCC.n5716 3.4105
R42556 VCC.n5718 VCC.n5711 3.4105
R42557 VCC.n5803 VCC.n5802 3.4105
R42558 VCC.n5802 VCC.n5801 3.4105
R42559 VCC.n5765 VCC.n5764 3.4105
R42560 VCC.n5766 VCC.n5765 3.4105
R42561 VCC.n5787 VCC.n5786 3.4105
R42562 VCC.n5763 VCC.n5762 3.4105
R42563 VCC.n5762 VCC.n5761 3.4105
R42564 VCC.n6007 VCC.n6006 3.4105
R42565 VCC.n6006 VCC.n6005 3.4105
R42566 VCC.n6066 VCC.n6065 3.4105
R42567 VCC.n6071 VCC.n6070 3.4105
R42568 VCC.n6070 VCC.n6069 3.4105
R42569 VCC.n6049 VCC.n6048 3.4105
R42570 VCC.n6050 VCC.n6049 3.4105
R42571 VCC.n6047 VCC.n6046 3.4105
R42572 VCC.n6064 VCC.n6063 3.4105
R42573 VCC.n6063 VCC.n6062 3.4105
R42574 VCC.n6036 VCC.n5589 3.4105
R42575 VCC.n5589 VCC.n5588 3.4105
R42576 VCC.n5587 VCC.n5586 3.4105
R42577 VCC.n6044 VCC.n6043 3.4105
R42578 VCC.n6043 VCC.n5582 3.4105
R42579 VCC.n6009 VCC.n6008 3.4105
R42580 VCC.n6009 VCC.n5605 3.4105
R42581 VCC.n6035 VCC.n6034 3.4105
R42582 VCC.n6073 VCC.n6072 3.4105
R42583 VCC.n6073 VCC.n5546 3.4105
R42584 VCC.n5990 VCC.n5989 3.4105
R42585 VCC.n5991 VCC.n5990 3.4105
R42586 VCC.n5954 VCC.n5953 3.4105
R42587 VCC.n5988 VCC.n5987 3.4105
R42588 VCC.n5987 VCC.n5986 3.4105
R42589 VCC.n5924 VCC.n5923 3.4105
R42590 VCC.n5923 VCC.n5922 3.4105
R42591 VCC.n5919 VCC.n5917 3.4105
R42592 VCC.n5952 VCC.n5951 3.4105
R42593 VCC.n5951 VCC.n5950 3.4105
R42594 VCC.n5648 VCC.n5647 3.4105
R42595 VCC.n5895 VCC.n5648 3.4105
R42596 VCC.n5916 VCC.n5645 3.4105
R42597 VCC.n5926 VCC.n5925 3.4105
R42598 VCC.n5926 VCC.n5644 3.4105
R42599 VCC.n5889 VCC.n5659 3.4105
R42600 VCC.n5889 VCC.n5888 3.4105
R42601 VCC.n5893 VCC.n5892 3.4105
R42602 VCC.n5864 VCC.n5863 3.4105
R42603 VCC.n5864 VCC.n5670 3.4105
R42604 VCC.n6635 VCC.n6634 3.4105
R42605 VCC.n6635 VCC.n6101 3.4105
R42606 VCC.n6611 VCC.n6610 3.4105
R42607 VCC.n6633 VCC.n6632 3.4105
R42608 VCC.n6632 VCC.n6631 3.4105
R42609 VCC.n6601 VCC.n6130 3.4105
R42610 VCC.n6130 VCC.n6129 3.4105
R42611 VCC.n6603 VCC.n6602 3.4105
R42612 VCC.n6609 VCC.n6608 3.4105
R42613 VCC.n6608 VCC.n6607 3.4105
R42614 VCC.n6583 VCC.n6582 3.4105
R42615 VCC.n6583 VCC.n6142 3.4105
R42616 VCC.n6579 VCC.n6132 3.4105
R42617 VCC.n6600 VCC.n6599 3.4105
R42618 VCC.n6599 VCC.n6598 3.4105
R42619 VCC.n6561 VCC.n6558 3.4105
R42620 VCC.n6561 VCC.n6560 3.4105
R42621 VCC.n6578 VCC.n6577 3.4105
R42622 VCC.n6557 VCC.n6556 3.4105
R42623 VCC.n6556 VCC.n6555 3.4105
R42624 VCC.n6541 VCC.n6540 3.4105
R42625 VCC.n6542 VCC.n6541 3.4105
R42626 VCC.n6506 VCC.n6505 3.4105
R42627 VCC.n6539 VCC.n6538 3.4105
R42628 VCC.n6538 VCC.n6537 3.4105
R42629 VCC.n6476 VCC.n6475 3.4105
R42630 VCC.n6475 VCC.n6474 3.4105
R42631 VCC.n6471 VCC.n6469 3.4105
R42632 VCC.n6504 VCC.n6503 3.4105
R42633 VCC.n6503 VCC.n6502 3.4105
R42634 VCC.n6200 VCC.n6199 3.4105
R42635 VCC.n6447 VCC.n6200 3.4105
R42636 VCC.n6468 VCC.n6197 3.4105
R42637 VCC.n6478 VCC.n6477 3.4105
R42638 VCC.n6478 VCC.n6196 3.4105
R42639 VCC.n6441 VCC.n6211 3.4105
R42640 VCC.n6441 VCC.n6440 3.4105
R42641 VCC.n6445 VCC.n6444 3.4105
R42642 VCC.n6415 VCC.n6414 3.4105
R42643 VCC.n6415 VCC.n6222 3.4105
R42644 VCC.n6406 VCC.n6405 3.4105
R42645 VCC.n6407 VCC.n6406 3.4105
R42646 VCC.n6379 VCC.n6378 3.4105
R42647 VCC.n6404 VCC.n6403 3.4105
R42648 VCC.n6403 VCC.n6402 3.4105
R42649 VCC.n6355 VCC.n6260 3.4105
R42650 VCC.n6260 VCC.n6254 3.4105
R42651 VCC.n6357 VCC.n6356 3.4105
R42652 VCC.n6377 VCC.n6376 3.4105
R42653 VCC.n6376 VCC.n6375 3.4105
R42654 VCC.n6339 VCC.n6268 3.4105
R42655 VCC.n6268 VCC.n6267 3.4105
R42656 VCC.n6269 VCC.n6262 3.4105
R42657 VCC.n6354 VCC.n6353 3.4105
R42658 VCC.n6353 VCC.n6352 3.4105
R42659 VCC.n6316 VCC.n6315 3.4105
R42660 VCC.n6317 VCC.n6316 3.4105
R42661 VCC.n6338 VCC.n6337 3.4105
R42662 VCC.n6314 VCC.n6313 3.4105
R42663 VCC.n6313 VCC.n6312 3.4105
R42664 VCC.n6964 VCC.n6963 3.4105
R42665 VCC.n6965 VCC.n6964 3.4105
R42666 VCC.n6937 VCC.n6936 3.4105
R42667 VCC.n6962 VCC.n6961 3.4105
R42668 VCC.n6961 VCC.n6960 3.4105
R42669 VCC.n6913 VCC.n6818 3.4105
R42670 VCC.n6818 VCC.n6812 3.4105
R42671 VCC.n6915 VCC.n6914 3.4105
R42672 VCC.n6935 VCC.n6934 3.4105
R42673 VCC.n6934 VCC.n6933 3.4105
R42674 VCC.n6897 VCC.n6826 3.4105
R42675 VCC.n6826 VCC.n6825 3.4105
R42676 VCC.n6827 VCC.n6820 3.4105
R42677 VCC.n6912 VCC.n6911 3.4105
R42678 VCC.n6911 VCC.n6910 3.4105
R42679 VCC.n6874 VCC.n6873 3.4105
R42680 VCC.n6875 VCC.n6874 3.4105
R42681 VCC.n6896 VCC.n6895 3.4105
R42682 VCC.n6872 VCC.n6871 3.4105
R42683 VCC.n6871 VCC.n6870 3.4105
R42684 VCC.n7116 VCC.n7115 3.4105
R42685 VCC.n7115 VCC.n7114 3.4105
R42686 VCC.n7175 VCC.n7174 3.4105
R42687 VCC.n7180 VCC.n7179 3.4105
R42688 VCC.n7179 VCC.n7178 3.4105
R42689 VCC.n7158 VCC.n7157 3.4105
R42690 VCC.n7159 VCC.n7158 3.4105
R42691 VCC.n7156 VCC.n7155 3.4105
R42692 VCC.n7173 VCC.n7172 3.4105
R42693 VCC.n7172 VCC.n7171 3.4105
R42694 VCC.n7145 VCC.n6698 3.4105
R42695 VCC.n6698 VCC.n6697 3.4105
R42696 VCC.n6696 VCC.n6695 3.4105
R42697 VCC.n7153 VCC.n7152 3.4105
R42698 VCC.n7152 VCC.n6691 3.4105
R42699 VCC.n7118 VCC.n7117 3.4105
R42700 VCC.n7118 VCC.n6714 3.4105
R42701 VCC.n7144 VCC.n7143 3.4105
R42702 VCC.n7182 VCC.n7181 3.4105
R42703 VCC.n7182 VCC.n6655 3.4105
R42704 VCC.n7099 VCC.n7098 3.4105
R42705 VCC.n7100 VCC.n7099 3.4105
R42706 VCC.n7063 VCC.n7062 3.4105
R42707 VCC.n7097 VCC.n7096 3.4105
R42708 VCC.n7096 VCC.n7095 3.4105
R42709 VCC.n7033 VCC.n7032 3.4105
R42710 VCC.n7032 VCC.n7031 3.4105
R42711 VCC.n7028 VCC.n7026 3.4105
R42712 VCC.n7061 VCC.n7060 3.4105
R42713 VCC.n7060 VCC.n7059 3.4105
R42714 VCC.n6757 VCC.n6756 3.4105
R42715 VCC.n7004 VCC.n6757 3.4105
R42716 VCC.n7025 VCC.n6754 3.4105
R42717 VCC.n7035 VCC.n7034 3.4105
R42718 VCC.n7035 VCC.n6753 3.4105
R42719 VCC.n6998 VCC.n6768 3.4105
R42720 VCC.n6998 VCC.n6997 3.4105
R42721 VCC.n7002 VCC.n7001 3.4105
R42722 VCC.n6973 VCC.n6972 3.4105
R42723 VCC.n6973 VCC.n6779 3.4105
R42724 VCC.n7744 VCC.n7743 3.4105
R42725 VCC.n7744 VCC.n7210 3.4105
R42726 VCC.n7720 VCC.n7719 3.4105
R42727 VCC.n7742 VCC.n7741 3.4105
R42728 VCC.n7741 VCC.n7740 3.4105
R42729 VCC.n7710 VCC.n7239 3.4105
R42730 VCC.n7239 VCC.n7238 3.4105
R42731 VCC.n7712 VCC.n7711 3.4105
R42732 VCC.n7718 VCC.n7717 3.4105
R42733 VCC.n7717 VCC.n7716 3.4105
R42734 VCC.n7692 VCC.n7691 3.4105
R42735 VCC.n7692 VCC.n7251 3.4105
R42736 VCC.n7688 VCC.n7241 3.4105
R42737 VCC.n7709 VCC.n7708 3.4105
R42738 VCC.n7708 VCC.n7707 3.4105
R42739 VCC.n7670 VCC.n7667 3.4105
R42740 VCC.n7670 VCC.n7669 3.4105
R42741 VCC.n7687 VCC.n7686 3.4105
R42742 VCC.n7666 VCC.n7665 3.4105
R42743 VCC.n7665 VCC.n7664 3.4105
R42744 VCC.n7650 VCC.n7649 3.4105
R42745 VCC.n7651 VCC.n7650 3.4105
R42746 VCC.n7615 VCC.n7614 3.4105
R42747 VCC.n7648 VCC.n7647 3.4105
R42748 VCC.n7647 VCC.n7646 3.4105
R42749 VCC.n7585 VCC.n7584 3.4105
R42750 VCC.n7584 VCC.n7583 3.4105
R42751 VCC.n7580 VCC.n7578 3.4105
R42752 VCC.n7613 VCC.n7612 3.4105
R42753 VCC.n7612 VCC.n7611 3.4105
R42754 VCC.n7309 VCC.n7308 3.4105
R42755 VCC.n7556 VCC.n7309 3.4105
R42756 VCC.n7577 VCC.n7306 3.4105
R42757 VCC.n7587 VCC.n7586 3.4105
R42758 VCC.n7587 VCC.n7305 3.4105
R42759 VCC.n7550 VCC.n7320 3.4105
R42760 VCC.n7550 VCC.n7549 3.4105
R42761 VCC.n7554 VCC.n7553 3.4105
R42762 VCC.n7524 VCC.n7523 3.4105
R42763 VCC.n7524 VCC.n7331 3.4105
R42764 VCC.n7515 VCC.n7514 3.4105
R42765 VCC.n7516 VCC.n7515 3.4105
R42766 VCC.n7488 VCC.n7487 3.4105
R42767 VCC.n7513 VCC.n7512 3.4105
R42768 VCC.n7512 VCC.n7511 3.4105
R42769 VCC.n7464 VCC.n7369 3.4105
R42770 VCC.n7369 VCC.n7363 3.4105
R42771 VCC.n7466 VCC.n7465 3.4105
R42772 VCC.n7486 VCC.n7485 3.4105
R42773 VCC.n7485 VCC.n7484 3.4105
R42774 VCC.n7448 VCC.n7377 3.4105
R42775 VCC.n7377 VCC.n7376 3.4105
R42776 VCC.n7378 VCC.n7371 3.4105
R42777 VCC.n7463 VCC.n7462 3.4105
R42778 VCC.n7462 VCC.n7461 3.4105
R42779 VCC.n7425 VCC.n7424 3.4105
R42780 VCC.n7426 VCC.n7425 3.4105
R42781 VCC.n7447 VCC.n7446 3.4105
R42782 VCC.n7423 VCC.n7422 3.4105
R42783 VCC.n7422 VCC.n7421 3.4105
R42784 VCC.n8073 VCC.n8072 3.4105
R42785 VCC.n8074 VCC.n8073 3.4105
R42786 VCC.n8046 VCC.n8045 3.4105
R42787 VCC.n8071 VCC.n8070 3.4105
R42788 VCC.n8070 VCC.n8069 3.4105
R42789 VCC.n8022 VCC.n7927 3.4105
R42790 VCC.n7927 VCC.n7921 3.4105
R42791 VCC.n8024 VCC.n8023 3.4105
R42792 VCC.n8044 VCC.n8043 3.4105
R42793 VCC.n8043 VCC.n8042 3.4105
R42794 VCC.n8006 VCC.n7935 3.4105
R42795 VCC.n7935 VCC.n7934 3.4105
R42796 VCC.n7936 VCC.n7929 3.4105
R42797 VCC.n8021 VCC.n8020 3.4105
R42798 VCC.n8020 VCC.n8019 3.4105
R42799 VCC.n7983 VCC.n7982 3.4105
R42800 VCC.n7984 VCC.n7983 3.4105
R42801 VCC.n8005 VCC.n8004 3.4105
R42802 VCC.n7981 VCC.n7980 3.4105
R42803 VCC.n7980 VCC.n7979 3.4105
R42804 VCC.n8225 VCC.n8224 3.4105
R42805 VCC.n8224 VCC.n8223 3.4105
R42806 VCC.n8284 VCC.n8283 3.4105
R42807 VCC.n8289 VCC.n8288 3.4105
R42808 VCC.n8288 VCC.n8287 3.4105
R42809 VCC.n8267 VCC.n8266 3.4105
R42810 VCC.n8268 VCC.n8267 3.4105
R42811 VCC.n8265 VCC.n8264 3.4105
R42812 VCC.n8282 VCC.n8281 3.4105
R42813 VCC.n8281 VCC.n8280 3.4105
R42814 VCC.n8254 VCC.n7807 3.4105
R42815 VCC.n7807 VCC.n7806 3.4105
R42816 VCC.n7805 VCC.n7804 3.4105
R42817 VCC.n8262 VCC.n8261 3.4105
R42818 VCC.n8261 VCC.n7800 3.4105
R42819 VCC.n8227 VCC.n8226 3.4105
R42820 VCC.n8227 VCC.n7823 3.4105
R42821 VCC.n8253 VCC.n8252 3.4105
R42822 VCC.n8291 VCC.n8290 3.4105
R42823 VCC.n8291 VCC.n7764 3.4105
R42824 VCC.n8208 VCC.n8207 3.4105
R42825 VCC.n8209 VCC.n8208 3.4105
R42826 VCC.n8172 VCC.n8171 3.4105
R42827 VCC.n8206 VCC.n8205 3.4105
R42828 VCC.n8205 VCC.n8204 3.4105
R42829 VCC.n8142 VCC.n8141 3.4105
R42830 VCC.n8141 VCC.n8140 3.4105
R42831 VCC.n8137 VCC.n8135 3.4105
R42832 VCC.n8170 VCC.n8169 3.4105
R42833 VCC.n8169 VCC.n8168 3.4105
R42834 VCC.n7866 VCC.n7865 3.4105
R42835 VCC.n8113 VCC.n7866 3.4105
R42836 VCC.n8134 VCC.n7863 3.4105
R42837 VCC.n8144 VCC.n8143 3.4105
R42838 VCC.n8144 VCC.n7862 3.4105
R42839 VCC.n8107 VCC.n7877 3.4105
R42840 VCC.n8107 VCC.n8106 3.4105
R42841 VCC.n8111 VCC.n8110 3.4105
R42842 VCC.n8082 VCC.n8081 3.4105
R42843 VCC.n8082 VCC.n7888 3.4105
R42844 VCC.n8624 VCC.n8623 3.4105
R42845 VCC.n8625 VCC.n8624 3.4105
R42846 VCC.n8597 VCC.n8596 3.4105
R42847 VCC.n8622 VCC.n8621 3.4105
R42848 VCC.n8621 VCC.n8620 3.4105
R42849 VCC.n8573 VCC.n8478 3.4105
R42850 VCC.n8478 VCC.n8472 3.4105
R42851 VCC.n8575 VCC.n8574 3.4105
R42852 VCC.n8595 VCC.n8594 3.4105
R42853 VCC.n8594 VCC.n8593 3.4105
R42854 VCC.n8557 VCC.n8486 3.4105
R42855 VCC.n8486 VCC.n8485 3.4105
R42856 VCC.n8487 VCC.n8480 3.4105
R42857 VCC.n8572 VCC.n8571 3.4105
R42858 VCC.n8571 VCC.n8570 3.4105
R42859 VCC.n8534 VCC.n8533 3.4105
R42860 VCC.n8535 VCC.n8534 3.4105
R42861 VCC.n8556 VCC.n8555 3.4105
R42862 VCC.n8532 VCC.n8531 3.4105
R42863 VCC.n8531 VCC.n8530 3.4105
R42864 VCC.n8853 VCC.n8852 3.4105
R42865 VCC.n8853 VCC.n8319 3.4105
R42866 VCC.n8829 VCC.n8828 3.4105
R42867 VCC.n8851 VCC.n8850 3.4105
R42868 VCC.n8850 VCC.n8849 3.4105
R42869 VCC.n8819 VCC.n8348 3.4105
R42870 VCC.n8348 VCC.n8347 3.4105
R42871 VCC.n8821 VCC.n8820 3.4105
R42872 VCC.n8827 VCC.n8826 3.4105
R42873 VCC.n8826 VCC.n8825 3.4105
R42874 VCC.n8801 VCC.n8800 3.4105
R42875 VCC.n8801 VCC.n8360 3.4105
R42876 VCC.n8797 VCC.n8350 3.4105
R42877 VCC.n8818 VCC.n8817 3.4105
R42878 VCC.n8817 VCC.n8816 3.4105
R42879 VCC.n8779 VCC.n8776 3.4105
R42880 VCC.n8779 VCC.n8778 3.4105
R42881 VCC.n8796 VCC.n8795 3.4105
R42882 VCC.n8775 VCC.n8774 3.4105
R42883 VCC.n8774 VCC.n8773 3.4105
R42884 VCC.n8759 VCC.n8758 3.4105
R42885 VCC.n8760 VCC.n8759 3.4105
R42886 VCC.n8724 VCC.n8723 3.4105
R42887 VCC.n8757 VCC.n8756 3.4105
R42888 VCC.n8756 VCC.n8755 3.4105
R42889 VCC.n8694 VCC.n8693 3.4105
R42890 VCC.n8693 VCC.n8692 3.4105
R42891 VCC.n8689 VCC.n8687 3.4105
R42892 VCC.n8722 VCC.n8721 3.4105
R42893 VCC.n8721 VCC.n8720 3.4105
R42894 VCC.n8418 VCC.n8417 3.4105
R42895 VCC.n8665 VCC.n8418 3.4105
R42896 VCC.n8686 VCC.n8415 3.4105
R42897 VCC.n8696 VCC.n8695 3.4105
R42898 VCC.n8696 VCC.n8414 3.4105
R42899 VCC.n8659 VCC.n8429 3.4105
R42900 VCC.n8659 VCC.n8658 3.4105
R42901 VCC.n8663 VCC.n8662 3.4105
R42902 VCC.n8633 VCC.n8632 3.4105
R42903 VCC.n8633 VCC.n8440 3.4105
R42904 VCC.n9182 VCC.n9181 3.4105
R42905 VCC.n9183 VCC.n9182 3.4105
R42906 VCC.n9155 VCC.n9154 3.4105
R42907 VCC.n9180 VCC.n9179 3.4105
R42908 VCC.n9179 VCC.n9178 3.4105
R42909 VCC.n9131 VCC.n9036 3.4105
R42910 VCC.n9036 VCC.n9030 3.4105
R42911 VCC.n9133 VCC.n9132 3.4105
R42912 VCC.n9153 VCC.n9152 3.4105
R42913 VCC.n9152 VCC.n9151 3.4105
R42914 VCC.n9115 VCC.n9044 3.4105
R42915 VCC.n9044 VCC.n9043 3.4105
R42916 VCC.n9045 VCC.n9038 3.4105
R42917 VCC.n9130 VCC.n9129 3.4105
R42918 VCC.n9129 VCC.n9128 3.4105
R42919 VCC.n9092 VCC.n9091 3.4105
R42920 VCC.n9093 VCC.n9092 3.4105
R42921 VCC.n9114 VCC.n9113 3.4105
R42922 VCC.n9090 VCC.n9089 3.4105
R42923 VCC.n9089 VCC.n9088 3.4105
R42924 VCC.n9334 VCC.n9333 3.4105
R42925 VCC.n9333 VCC.n9332 3.4105
R42926 VCC.n9393 VCC.n9392 3.4105
R42927 VCC.n9398 VCC.n9397 3.4105
R42928 VCC.n9397 VCC.n9396 3.4105
R42929 VCC.n9376 VCC.n9375 3.4105
R42930 VCC.n9377 VCC.n9376 3.4105
R42931 VCC.n9374 VCC.n9373 3.4105
R42932 VCC.n9391 VCC.n9390 3.4105
R42933 VCC.n9390 VCC.n9389 3.4105
R42934 VCC.n9363 VCC.n8916 3.4105
R42935 VCC.n8916 VCC.n8915 3.4105
R42936 VCC.n8914 VCC.n8913 3.4105
R42937 VCC.n9371 VCC.n9370 3.4105
R42938 VCC.n9370 VCC.n8909 3.4105
R42939 VCC.n9336 VCC.n9335 3.4105
R42940 VCC.n9336 VCC.n8932 3.4105
R42941 VCC.n9362 VCC.n9361 3.4105
R42942 VCC.n9400 VCC.n9399 3.4105
R42943 VCC.n9400 VCC.n8873 3.4105
R42944 VCC.n9317 VCC.n9316 3.4105
R42945 VCC.n9318 VCC.n9317 3.4105
R42946 VCC.n9281 VCC.n9280 3.4105
R42947 VCC.n9315 VCC.n9314 3.4105
R42948 VCC.n9314 VCC.n9313 3.4105
R42949 VCC.n9251 VCC.n9250 3.4105
R42950 VCC.n9250 VCC.n9249 3.4105
R42951 VCC.n9246 VCC.n9244 3.4105
R42952 VCC.n9279 VCC.n9278 3.4105
R42953 VCC.n9278 VCC.n9277 3.4105
R42954 VCC.n8975 VCC.n8974 3.4105
R42955 VCC.n9222 VCC.n8975 3.4105
R42956 VCC.n9243 VCC.n8972 3.4105
R42957 VCC.n9253 VCC.n9252 3.4105
R42958 VCC.n9253 VCC.n8971 3.4105
R42959 VCC.n9216 VCC.n8986 3.4105
R42960 VCC.n9216 VCC.n9215 3.4105
R42961 VCC.n9220 VCC.n9219 3.4105
R42962 VCC.n9191 VCC.n9190 3.4105
R42963 VCC.n9191 VCC.n8997 3.4105
R42964 VCC.n9962 VCC.n9961 3.4105
R42965 VCC.n9962 VCC.n9428 3.4105
R42966 VCC.n9938 VCC.n9937 3.4105
R42967 VCC.n9960 VCC.n9959 3.4105
R42968 VCC.n9959 VCC.n9958 3.4105
R42969 VCC.n9928 VCC.n9457 3.4105
R42970 VCC.n9457 VCC.n9456 3.4105
R42971 VCC.n9930 VCC.n9929 3.4105
R42972 VCC.n9936 VCC.n9935 3.4105
R42973 VCC.n9935 VCC.n9934 3.4105
R42974 VCC.n9910 VCC.n9909 3.4105
R42975 VCC.n9910 VCC.n9469 3.4105
R42976 VCC.n9906 VCC.n9459 3.4105
R42977 VCC.n9927 VCC.n9926 3.4105
R42978 VCC.n9926 VCC.n9925 3.4105
R42979 VCC.n9888 VCC.n9885 3.4105
R42980 VCC.n9888 VCC.n9887 3.4105
R42981 VCC.n9905 VCC.n9904 3.4105
R42982 VCC.n9884 VCC.n9883 3.4105
R42983 VCC.n9883 VCC.n9882 3.4105
R42984 VCC.n9868 VCC.n9867 3.4105
R42985 VCC.n9869 VCC.n9868 3.4105
R42986 VCC.n9833 VCC.n9832 3.4105
R42987 VCC.n9866 VCC.n9865 3.4105
R42988 VCC.n9865 VCC.n9864 3.4105
R42989 VCC.n9803 VCC.n9802 3.4105
R42990 VCC.n9802 VCC.n9801 3.4105
R42991 VCC.n9798 VCC.n9796 3.4105
R42992 VCC.n9831 VCC.n9830 3.4105
R42993 VCC.n9830 VCC.n9829 3.4105
R42994 VCC.n9527 VCC.n9526 3.4105
R42995 VCC.n9774 VCC.n9527 3.4105
R42996 VCC.n9795 VCC.n9524 3.4105
R42997 VCC.n9805 VCC.n9804 3.4105
R42998 VCC.n9805 VCC.n9523 3.4105
R42999 VCC.n9768 VCC.n9538 3.4105
R43000 VCC.n9768 VCC.n9767 3.4105
R43001 VCC.n9772 VCC.n9771 3.4105
R43002 VCC.n9742 VCC.n9741 3.4105
R43003 VCC.n9742 VCC.n9549 3.4105
R43004 VCC.n9733 VCC.n9732 3.4105
R43005 VCC.n9734 VCC.n9733 3.4105
R43006 VCC.n9706 VCC.n9705 3.4105
R43007 VCC.n9731 VCC.n9730 3.4105
R43008 VCC.n9730 VCC.n9729 3.4105
R43009 VCC.n9682 VCC.n9587 3.4105
R43010 VCC.n9587 VCC.n9581 3.4105
R43011 VCC.n9684 VCC.n9683 3.4105
R43012 VCC.n9704 VCC.n9703 3.4105
R43013 VCC.n9703 VCC.n9702 3.4105
R43014 VCC.n9666 VCC.n9595 3.4105
R43015 VCC.n9595 VCC.n9594 3.4105
R43016 VCC.n9596 VCC.n9589 3.4105
R43017 VCC.n9681 VCC.n9680 3.4105
R43018 VCC.n9680 VCC.n9679 3.4105
R43019 VCC.n9643 VCC.n9642 3.4105
R43020 VCC.n9644 VCC.n9643 3.4105
R43021 VCC.n9665 VCC.n9664 3.4105
R43022 VCC.n9641 VCC.n9640 3.4105
R43023 VCC.n9640 VCC.n9639 3.4105
R43024 VCC.n10290 VCC.n10289 3.4105
R43025 VCC.n10291 VCC.n10290 3.4105
R43026 VCC.n10263 VCC.n10262 3.4105
R43027 VCC.n10288 VCC.n10287 3.4105
R43028 VCC.n10287 VCC.n10286 3.4105
R43029 VCC.n10239 VCC.n10144 3.4105
R43030 VCC.n10144 VCC.n10138 3.4105
R43031 VCC.n10241 VCC.n10240 3.4105
R43032 VCC.n10261 VCC.n10260 3.4105
R43033 VCC.n10260 VCC.n10259 3.4105
R43034 VCC.n10223 VCC.n10152 3.4105
R43035 VCC.n10152 VCC.n10151 3.4105
R43036 VCC.n10153 VCC.n10146 3.4105
R43037 VCC.n10238 VCC.n10237 3.4105
R43038 VCC.n10237 VCC.n10236 3.4105
R43039 VCC.n10200 VCC.n10199 3.4105
R43040 VCC.n10201 VCC.n10200 3.4105
R43041 VCC.n10222 VCC.n10221 3.4105
R43042 VCC.n10198 VCC.n10197 3.4105
R43043 VCC.n10197 VCC.n10196 3.4105
R43044 VCC.n10442 VCC.n10441 3.4105
R43045 VCC.n10441 VCC.n10440 3.4105
R43046 VCC.n10501 VCC.n10500 3.4105
R43047 VCC.n10506 VCC.n10505 3.4105
R43048 VCC.n10505 VCC.n10504 3.4105
R43049 VCC.n10484 VCC.n10483 3.4105
R43050 VCC.n10485 VCC.n10484 3.4105
R43051 VCC.n10482 VCC.n10481 3.4105
R43052 VCC.n10499 VCC.n10498 3.4105
R43053 VCC.n10498 VCC.n10497 3.4105
R43054 VCC.n10471 VCC.n10024 3.4105
R43055 VCC.n10024 VCC.n10023 3.4105
R43056 VCC.n10022 VCC.n10021 3.4105
R43057 VCC.n10479 VCC.n10478 3.4105
R43058 VCC.n10478 VCC.n10017 3.4105
R43059 VCC.n10444 VCC.n10443 3.4105
R43060 VCC.n10444 VCC.n10040 3.4105
R43061 VCC.n10470 VCC.n10469 3.4105
R43062 VCC.n10508 VCC.n10507 3.4105
R43063 VCC.n10508 VCC.n9981 3.4105
R43064 VCC.n10425 VCC.n10424 3.4105
R43065 VCC.n10426 VCC.n10425 3.4105
R43066 VCC.n10389 VCC.n10388 3.4105
R43067 VCC.n10423 VCC.n10422 3.4105
R43068 VCC.n10422 VCC.n10421 3.4105
R43069 VCC.n10359 VCC.n10358 3.4105
R43070 VCC.n10358 VCC.n10357 3.4105
R43071 VCC.n10354 VCC.n10352 3.4105
R43072 VCC.n10387 VCC.n10386 3.4105
R43073 VCC.n10386 VCC.n10385 3.4105
R43074 VCC.n10083 VCC.n10082 3.4105
R43075 VCC.n10330 VCC.n10083 3.4105
R43076 VCC.n10351 VCC.n10080 3.4105
R43077 VCC.n10361 VCC.n10360 3.4105
R43078 VCC.n10361 VCC.n10079 3.4105
R43079 VCC.n10324 VCC.n10094 3.4105
R43080 VCC.n10324 VCC.n10323 3.4105
R43081 VCC.n10328 VCC.n10327 3.4105
R43082 VCC.n10299 VCC.n10298 3.4105
R43083 VCC.n10299 VCC.n10105 3.4105
R43084 VCC.n11069 VCC.n11068 3.4105
R43085 VCC.n11069 VCC.n10535 3.4105
R43086 VCC.n11045 VCC.n11044 3.4105
R43087 VCC.n11067 VCC.n11066 3.4105
R43088 VCC.n11066 VCC.n11065 3.4105
R43089 VCC.n11035 VCC.n10564 3.4105
R43090 VCC.n10564 VCC.n10563 3.4105
R43091 VCC.n11037 VCC.n11036 3.4105
R43092 VCC.n11043 VCC.n11042 3.4105
R43093 VCC.n11042 VCC.n11041 3.4105
R43094 VCC.n11017 VCC.n11016 3.4105
R43095 VCC.n11017 VCC.n10576 3.4105
R43096 VCC.n11013 VCC.n10566 3.4105
R43097 VCC.n11034 VCC.n11033 3.4105
R43098 VCC.n11033 VCC.n11032 3.4105
R43099 VCC.n10995 VCC.n10992 3.4105
R43100 VCC.n10995 VCC.n10994 3.4105
R43101 VCC.n11012 VCC.n11011 3.4105
R43102 VCC.n10991 VCC.n10990 3.4105
R43103 VCC.n10990 VCC.n10989 3.4105
R43104 VCC.n10975 VCC.n10974 3.4105
R43105 VCC.n10976 VCC.n10975 3.4105
R43106 VCC.n10940 VCC.n10939 3.4105
R43107 VCC.n10973 VCC.n10972 3.4105
R43108 VCC.n10972 VCC.n10971 3.4105
R43109 VCC.n10910 VCC.n10909 3.4105
R43110 VCC.n10909 VCC.n10908 3.4105
R43111 VCC.n10905 VCC.n10903 3.4105
R43112 VCC.n10938 VCC.n10937 3.4105
R43113 VCC.n10937 VCC.n10936 3.4105
R43114 VCC.n10634 VCC.n10633 3.4105
R43115 VCC.n10881 VCC.n10634 3.4105
R43116 VCC.n10902 VCC.n10631 3.4105
R43117 VCC.n10912 VCC.n10911 3.4105
R43118 VCC.n10912 VCC.n10630 3.4105
R43119 VCC.n10875 VCC.n10645 3.4105
R43120 VCC.n10875 VCC.n10874 3.4105
R43121 VCC.n10879 VCC.n10878 3.4105
R43122 VCC.n10849 VCC.n10848 3.4105
R43123 VCC.n10849 VCC.n10656 3.4105
R43124 VCC.n10840 VCC.n10839 3.4105
R43125 VCC.n10841 VCC.n10840 3.4105
R43126 VCC.n10813 VCC.n10812 3.4105
R43127 VCC.n10838 VCC.n10837 3.4105
R43128 VCC.n10837 VCC.n10836 3.4105
R43129 VCC.n10789 VCC.n10694 3.4105
R43130 VCC.n10694 VCC.n10688 3.4105
R43131 VCC.n10791 VCC.n10790 3.4105
R43132 VCC.n10811 VCC.n10810 3.4105
R43133 VCC.n10810 VCC.n10809 3.4105
R43134 VCC.n10773 VCC.n10702 3.4105
R43135 VCC.n10702 VCC.n10701 3.4105
R43136 VCC.n10703 VCC.n10696 3.4105
R43137 VCC.n10788 VCC.n10787 3.4105
R43138 VCC.n10787 VCC.n10786 3.4105
R43139 VCC.n10750 VCC.n10749 3.4105
R43140 VCC.n10751 VCC.n10750 3.4105
R43141 VCC.n10772 VCC.n10771 3.4105
R43142 VCC.n10748 VCC.n10747 3.4105
R43143 VCC.n10747 VCC.n10746 3.4105
R43144 VCC.n11397 VCC.n11396 3.4105
R43145 VCC.n11398 VCC.n11397 3.4105
R43146 VCC.n11370 VCC.n11369 3.4105
R43147 VCC.n11395 VCC.n11394 3.4105
R43148 VCC.n11394 VCC.n11393 3.4105
R43149 VCC.n11346 VCC.n11251 3.4105
R43150 VCC.n11251 VCC.n11245 3.4105
R43151 VCC.n11348 VCC.n11347 3.4105
R43152 VCC.n11368 VCC.n11367 3.4105
R43153 VCC.n11367 VCC.n11366 3.4105
R43154 VCC.n11330 VCC.n11259 3.4105
R43155 VCC.n11259 VCC.n11258 3.4105
R43156 VCC.n11260 VCC.n11253 3.4105
R43157 VCC.n11345 VCC.n11344 3.4105
R43158 VCC.n11344 VCC.n11343 3.4105
R43159 VCC.n11307 VCC.n11306 3.4105
R43160 VCC.n11308 VCC.n11307 3.4105
R43161 VCC.n11329 VCC.n11328 3.4105
R43162 VCC.n11305 VCC.n11304 3.4105
R43163 VCC.n11304 VCC.n11303 3.4105
R43164 VCC.n11549 VCC.n11548 3.4105
R43165 VCC.n11548 VCC.n11547 3.4105
R43166 VCC.n11608 VCC.n11607 3.4105
R43167 VCC.n11613 VCC.n11612 3.4105
R43168 VCC.n11612 VCC.n11611 3.4105
R43169 VCC.n11591 VCC.n11590 3.4105
R43170 VCC.n11592 VCC.n11591 3.4105
R43171 VCC.n11589 VCC.n11588 3.4105
R43172 VCC.n11606 VCC.n11605 3.4105
R43173 VCC.n11605 VCC.n11604 3.4105
R43174 VCC.n11578 VCC.n11131 3.4105
R43175 VCC.n11131 VCC.n11130 3.4105
R43176 VCC.n11129 VCC.n11128 3.4105
R43177 VCC.n11586 VCC.n11585 3.4105
R43178 VCC.n11585 VCC.n11124 3.4105
R43179 VCC.n11551 VCC.n11550 3.4105
R43180 VCC.n11551 VCC.n11147 3.4105
R43181 VCC.n11577 VCC.n11576 3.4105
R43182 VCC.n11615 VCC.n11614 3.4105
R43183 VCC.n11615 VCC.n11088 3.4105
R43184 VCC.n11532 VCC.n11531 3.4105
R43185 VCC.n11533 VCC.n11532 3.4105
R43186 VCC.n11496 VCC.n11495 3.4105
R43187 VCC.n11530 VCC.n11529 3.4105
R43188 VCC.n11529 VCC.n11528 3.4105
R43189 VCC.n11466 VCC.n11465 3.4105
R43190 VCC.n11465 VCC.n11464 3.4105
R43191 VCC.n11461 VCC.n11459 3.4105
R43192 VCC.n11494 VCC.n11493 3.4105
R43193 VCC.n11493 VCC.n11492 3.4105
R43194 VCC.n11190 VCC.n11189 3.4105
R43195 VCC.n11437 VCC.n11190 3.4105
R43196 VCC.n11458 VCC.n11187 3.4105
R43197 VCC.n11468 VCC.n11467 3.4105
R43198 VCC.n11468 VCC.n11186 3.4105
R43199 VCC.n11431 VCC.n11201 3.4105
R43200 VCC.n11431 VCC.n11430 3.4105
R43201 VCC.n11435 VCC.n11434 3.4105
R43202 VCC.n11406 VCC.n11405 3.4105
R43203 VCC.n11406 VCC.n11212 3.4105
R43204 VCC.n12176 VCC.n12175 3.4105
R43205 VCC.n12176 VCC.n11642 3.4105
R43206 VCC.n12152 VCC.n12151 3.4105
R43207 VCC.n12174 VCC.n12173 3.4105
R43208 VCC.n12173 VCC.n12172 3.4105
R43209 VCC.n12142 VCC.n11671 3.4105
R43210 VCC.n11671 VCC.n11670 3.4105
R43211 VCC.n12144 VCC.n12143 3.4105
R43212 VCC.n12150 VCC.n12149 3.4105
R43213 VCC.n12149 VCC.n12148 3.4105
R43214 VCC.n12124 VCC.n12123 3.4105
R43215 VCC.n12124 VCC.n11683 3.4105
R43216 VCC.n12120 VCC.n11673 3.4105
R43217 VCC.n12141 VCC.n12140 3.4105
R43218 VCC.n12140 VCC.n12139 3.4105
R43219 VCC.n12102 VCC.n12099 3.4105
R43220 VCC.n12102 VCC.n12101 3.4105
R43221 VCC.n12119 VCC.n12118 3.4105
R43222 VCC.n12098 VCC.n12097 3.4105
R43223 VCC.n12097 VCC.n12096 3.4105
R43224 VCC.n12082 VCC.n12081 3.4105
R43225 VCC.n12083 VCC.n12082 3.4105
R43226 VCC.n12047 VCC.n12046 3.4105
R43227 VCC.n12080 VCC.n12079 3.4105
R43228 VCC.n12079 VCC.n12078 3.4105
R43229 VCC.n12017 VCC.n12016 3.4105
R43230 VCC.n12016 VCC.n12015 3.4105
R43231 VCC.n12012 VCC.n12010 3.4105
R43232 VCC.n12045 VCC.n12044 3.4105
R43233 VCC.n12044 VCC.n12043 3.4105
R43234 VCC.n11741 VCC.n11740 3.4105
R43235 VCC.n11988 VCC.n11741 3.4105
R43236 VCC.n12009 VCC.n11738 3.4105
R43237 VCC.n12019 VCC.n12018 3.4105
R43238 VCC.n12019 VCC.n11737 3.4105
R43239 VCC.n11982 VCC.n11752 3.4105
R43240 VCC.n11982 VCC.n11981 3.4105
R43241 VCC.n11986 VCC.n11985 3.4105
R43242 VCC.n11956 VCC.n11955 3.4105
R43243 VCC.n11956 VCC.n11763 3.4105
R43244 VCC.n11947 VCC.n11946 3.4105
R43245 VCC.n11948 VCC.n11947 3.4105
R43246 VCC.n11920 VCC.n11919 3.4105
R43247 VCC.n11945 VCC.n11944 3.4105
R43248 VCC.n11944 VCC.n11943 3.4105
R43249 VCC.n11896 VCC.n11801 3.4105
R43250 VCC.n11801 VCC.n11795 3.4105
R43251 VCC.n11898 VCC.n11897 3.4105
R43252 VCC.n11918 VCC.n11917 3.4105
R43253 VCC.n11917 VCC.n11916 3.4105
R43254 VCC.n11880 VCC.n11809 3.4105
R43255 VCC.n11809 VCC.n11808 3.4105
R43256 VCC.n11810 VCC.n11803 3.4105
R43257 VCC.n11895 VCC.n11894 3.4105
R43258 VCC.n11894 VCC.n11893 3.4105
R43259 VCC.n11857 VCC.n11856 3.4105
R43260 VCC.n11858 VCC.n11857 3.4105
R43261 VCC.n11879 VCC.n11878 3.4105
R43262 VCC.n11855 VCC.n11854 3.4105
R43263 VCC.n11854 VCC.n11853 3.4105
R43264 VCC.n12504 VCC.n12503 3.4105
R43265 VCC.n12505 VCC.n12504 3.4105
R43266 VCC.n12477 VCC.n12476 3.4105
R43267 VCC.n12502 VCC.n12501 3.4105
R43268 VCC.n12501 VCC.n12500 3.4105
R43269 VCC.n12453 VCC.n12358 3.4105
R43270 VCC.n12358 VCC.n12352 3.4105
R43271 VCC.n12455 VCC.n12454 3.4105
R43272 VCC.n12475 VCC.n12474 3.4105
R43273 VCC.n12474 VCC.n12473 3.4105
R43274 VCC.n12437 VCC.n12366 3.4105
R43275 VCC.n12366 VCC.n12365 3.4105
R43276 VCC.n12367 VCC.n12360 3.4105
R43277 VCC.n12452 VCC.n12451 3.4105
R43278 VCC.n12451 VCC.n12450 3.4105
R43279 VCC.n12414 VCC.n12413 3.4105
R43280 VCC.n12415 VCC.n12414 3.4105
R43281 VCC.n12436 VCC.n12435 3.4105
R43282 VCC.n12412 VCC.n12411 3.4105
R43283 VCC.n12411 VCC.n12410 3.4105
R43284 VCC.n12656 VCC.n12655 3.4105
R43285 VCC.n12655 VCC.n12654 3.4105
R43286 VCC.n12715 VCC.n12714 3.4105
R43287 VCC.n12720 VCC.n12719 3.4105
R43288 VCC.n12719 VCC.n12718 3.4105
R43289 VCC.n12698 VCC.n12697 3.4105
R43290 VCC.n12699 VCC.n12698 3.4105
R43291 VCC.n12696 VCC.n12695 3.4105
R43292 VCC.n12713 VCC.n12712 3.4105
R43293 VCC.n12712 VCC.n12711 3.4105
R43294 VCC.n12685 VCC.n12238 3.4105
R43295 VCC.n12238 VCC.n12237 3.4105
R43296 VCC.n12236 VCC.n12235 3.4105
R43297 VCC.n12693 VCC.n12692 3.4105
R43298 VCC.n12692 VCC.n12231 3.4105
R43299 VCC.n12658 VCC.n12657 3.4105
R43300 VCC.n12658 VCC.n12254 3.4105
R43301 VCC.n12684 VCC.n12683 3.4105
R43302 VCC.n12722 VCC.n12721 3.4105
R43303 VCC.n12722 VCC.n12195 3.4105
R43304 VCC.n12639 VCC.n12638 3.4105
R43305 VCC.n12640 VCC.n12639 3.4105
R43306 VCC.n12603 VCC.n12602 3.4105
R43307 VCC.n12637 VCC.n12636 3.4105
R43308 VCC.n12636 VCC.n12635 3.4105
R43309 VCC.n12573 VCC.n12572 3.4105
R43310 VCC.n12572 VCC.n12571 3.4105
R43311 VCC.n12568 VCC.n12566 3.4105
R43312 VCC.n12601 VCC.n12600 3.4105
R43313 VCC.n12600 VCC.n12599 3.4105
R43314 VCC.n12297 VCC.n12296 3.4105
R43315 VCC.n12544 VCC.n12297 3.4105
R43316 VCC.n12565 VCC.n12294 3.4105
R43317 VCC.n12575 VCC.n12574 3.4105
R43318 VCC.n12575 VCC.n12293 3.4105
R43319 VCC.n12538 VCC.n12308 3.4105
R43320 VCC.n12538 VCC.n12537 3.4105
R43321 VCC.n12542 VCC.n12541 3.4105
R43322 VCC.n12513 VCC.n12512 3.4105
R43323 VCC.n12513 VCC.n12319 3.4105
R43324 VCC.n13283 VCC.n13282 3.4105
R43325 VCC.n13283 VCC.n12749 3.4105
R43326 VCC.n13259 VCC.n13258 3.4105
R43327 VCC.n13281 VCC.n13280 3.4105
R43328 VCC.n13280 VCC.n13279 3.4105
R43329 VCC.n13249 VCC.n12778 3.4105
R43330 VCC.n12778 VCC.n12777 3.4105
R43331 VCC.n13251 VCC.n13250 3.4105
R43332 VCC.n13257 VCC.n13256 3.4105
R43333 VCC.n13256 VCC.n13255 3.4105
R43334 VCC.n13231 VCC.n13230 3.4105
R43335 VCC.n13231 VCC.n12790 3.4105
R43336 VCC.n13227 VCC.n12780 3.4105
R43337 VCC.n13248 VCC.n13247 3.4105
R43338 VCC.n13247 VCC.n13246 3.4105
R43339 VCC.n13209 VCC.n13206 3.4105
R43340 VCC.n13209 VCC.n13208 3.4105
R43341 VCC.n13226 VCC.n13225 3.4105
R43342 VCC.n13205 VCC.n13204 3.4105
R43343 VCC.n13204 VCC.n13203 3.4105
R43344 VCC.n13189 VCC.n13188 3.4105
R43345 VCC.n13190 VCC.n13189 3.4105
R43346 VCC.n13154 VCC.n13153 3.4105
R43347 VCC.n13187 VCC.n13186 3.4105
R43348 VCC.n13186 VCC.n13185 3.4105
R43349 VCC.n13124 VCC.n13123 3.4105
R43350 VCC.n13123 VCC.n13122 3.4105
R43351 VCC.n13119 VCC.n13117 3.4105
R43352 VCC.n13152 VCC.n13151 3.4105
R43353 VCC.n13151 VCC.n13150 3.4105
R43354 VCC.n12848 VCC.n12847 3.4105
R43355 VCC.n13095 VCC.n12848 3.4105
R43356 VCC.n13116 VCC.n12845 3.4105
R43357 VCC.n13126 VCC.n13125 3.4105
R43358 VCC.n13126 VCC.n12844 3.4105
R43359 VCC.n13089 VCC.n12859 3.4105
R43360 VCC.n13089 VCC.n13088 3.4105
R43361 VCC.n13093 VCC.n13092 3.4105
R43362 VCC.n13063 VCC.n13062 3.4105
R43363 VCC.n13063 VCC.n12870 3.4105
R43364 VCC.n13054 VCC.n13053 3.4105
R43365 VCC.n13055 VCC.n13054 3.4105
R43366 VCC.n13027 VCC.n13026 3.4105
R43367 VCC.n13052 VCC.n13051 3.4105
R43368 VCC.n13051 VCC.n13050 3.4105
R43369 VCC.n13003 VCC.n12908 3.4105
R43370 VCC.n12908 VCC.n12902 3.4105
R43371 VCC.n13005 VCC.n13004 3.4105
R43372 VCC.n13025 VCC.n13024 3.4105
R43373 VCC.n13024 VCC.n13023 3.4105
R43374 VCC.n12987 VCC.n12916 3.4105
R43375 VCC.n12916 VCC.n12915 3.4105
R43376 VCC.n12917 VCC.n12910 3.4105
R43377 VCC.n13002 VCC.n13001 3.4105
R43378 VCC.n13001 VCC.n13000 3.4105
R43379 VCC.n12964 VCC.n12963 3.4105
R43380 VCC.n12965 VCC.n12964 3.4105
R43381 VCC.n12986 VCC.n12985 3.4105
R43382 VCC.n12962 VCC.n12961 3.4105
R43383 VCC.n12961 VCC.n12960 3.4105
R43384 VCC.n13611 VCC.n13610 3.4105
R43385 VCC.n13612 VCC.n13611 3.4105
R43386 VCC.n13584 VCC.n13583 3.4105
R43387 VCC.n13609 VCC.n13608 3.4105
R43388 VCC.n13608 VCC.n13607 3.4105
R43389 VCC.n13560 VCC.n13465 3.4105
R43390 VCC.n13465 VCC.n13459 3.4105
R43391 VCC.n13562 VCC.n13561 3.4105
R43392 VCC.n13582 VCC.n13581 3.4105
R43393 VCC.n13581 VCC.n13580 3.4105
R43394 VCC.n13544 VCC.n13473 3.4105
R43395 VCC.n13473 VCC.n13472 3.4105
R43396 VCC.n13474 VCC.n13467 3.4105
R43397 VCC.n13559 VCC.n13558 3.4105
R43398 VCC.n13558 VCC.n13557 3.4105
R43399 VCC.n13521 VCC.n13520 3.4105
R43400 VCC.n13522 VCC.n13521 3.4105
R43401 VCC.n13543 VCC.n13542 3.4105
R43402 VCC.n13519 VCC.n13518 3.4105
R43403 VCC.n13518 VCC.n13517 3.4105
R43404 VCC.n13763 VCC.n13762 3.4105
R43405 VCC.n13762 VCC.n13761 3.4105
R43406 VCC.n13822 VCC.n13821 3.4105
R43407 VCC.n13827 VCC.n13826 3.4105
R43408 VCC.n13826 VCC.n13825 3.4105
R43409 VCC.n13805 VCC.n13804 3.4105
R43410 VCC.n13806 VCC.n13805 3.4105
R43411 VCC.n13803 VCC.n13802 3.4105
R43412 VCC.n13820 VCC.n13819 3.4105
R43413 VCC.n13819 VCC.n13818 3.4105
R43414 VCC.n13792 VCC.n13345 3.4105
R43415 VCC.n13345 VCC.n13344 3.4105
R43416 VCC.n13343 VCC.n13342 3.4105
R43417 VCC.n13800 VCC.n13799 3.4105
R43418 VCC.n13799 VCC.n13338 3.4105
R43419 VCC.n13765 VCC.n13764 3.4105
R43420 VCC.n13765 VCC.n13361 3.4105
R43421 VCC.n13791 VCC.n13790 3.4105
R43422 VCC.n13829 VCC.n13828 3.4105
R43423 VCC.n13829 VCC.n13302 3.4105
R43424 VCC.n13746 VCC.n13745 3.4105
R43425 VCC.n13747 VCC.n13746 3.4105
R43426 VCC.n13710 VCC.n13709 3.4105
R43427 VCC.n13744 VCC.n13743 3.4105
R43428 VCC.n13743 VCC.n13742 3.4105
R43429 VCC.n13680 VCC.n13679 3.4105
R43430 VCC.n13679 VCC.n13678 3.4105
R43431 VCC.n13675 VCC.n13673 3.4105
R43432 VCC.n13708 VCC.n13707 3.4105
R43433 VCC.n13707 VCC.n13706 3.4105
R43434 VCC.n13404 VCC.n13403 3.4105
R43435 VCC.n13651 VCC.n13404 3.4105
R43436 VCC.n13672 VCC.n13401 3.4105
R43437 VCC.n13682 VCC.n13681 3.4105
R43438 VCC.n13682 VCC.n13400 3.4105
R43439 VCC.n13645 VCC.n13415 3.4105
R43440 VCC.n13645 VCC.n13644 3.4105
R43441 VCC.n13649 VCC.n13648 3.4105
R43442 VCC.n13620 VCC.n13619 3.4105
R43443 VCC.n13620 VCC.n13426 3.4105
R43444 VCC.n14390 VCC.n14389 3.4105
R43445 VCC.n14390 VCC.n13856 3.4105
R43446 VCC.n14366 VCC.n14365 3.4105
R43447 VCC.n14388 VCC.n14387 3.4105
R43448 VCC.n14387 VCC.n14386 3.4105
R43449 VCC.n14356 VCC.n13885 3.4105
R43450 VCC.n13885 VCC.n13884 3.4105
R43451 VCC.n14358 VCC.n14357 3.4105
R43452 VCC.n14364 VCC.n14363 3.4105
R43453 VCC.n14363 VCC.n14362 3.4105
R43454 VCC.n14338 VCC.n14337 3.4105
R43455 VCC.n14338 VCC.n13897 3.4105
R43456 VCC.n14334 VCC.n13887 3.4105
R43457 VCC.n14355 VCC.n14354 3.4105
R43458 VCC.n14354 VCC.n14353 3.4105
R43459 VCC.n14316 VCC.n14313 3.4105
R43460 VCC.n14316 VCC.n14315 3.4105
R43461 VCC.n14333 VCC.n14332 3.4105
R43462 VCC.n14312 VCC.n14311 3.4105
R43463 VCC.n14311 VCC.n14310 3.4105
R43464 VCC.n14296 VCC.n14295 3.4105
R43465 VCC.n14297 VCC.n14296 3.4105
R43466 VCC.n14261 VCC.n14260 3.4105
R43467 VCC.n14294 VCC.n14293 3.4105
R43468 VCC.n14293 VCC.n14292 3.4105
R43469 VCC.n14231 VCC.n14230 3.4105
R43470 VCC.n14230 VCC.n14229 3.4105
R43471 VCC.n14226 VCC.n14224 3.4105
R43472 VCC.n14259 VCC.n14258 3.4105
R43473 VCC.n14258 VCC.n14257 3.4105
R43474 VCC.n13955 VCC.n13954 3.4105
R43475 VCC.n14202 VCC.n13955 3.4105
R43476 VCC.n14223 VCC.n13952 3.4105
R43477 VCC.n14233 VCC.n14232 3.4105
R43478 VCC.n14233 VCC.n13951 3.4105
R43479 VCC.n14196 VCC.n13966 3.4105
R43480 VCC.n14196 VCC.n14195 3.4105
R43481 VCC.n14200 VCC.n14199 3.4105
R43482 VCC.n14170 VCC.n14169 3.4105
R43483 VCC.n14170 VCC.n13977 3.4105
R43484 VCC.n14161 VCC.n14160 3.4105
R43485 VCC.n14162 VCC.n14161 3.4105
R43486 VCC.n14134 VCC.n14133 3.4105
R43487 VCC.n14159 VCC.n14158 3.4105
R43488 VCC.n14158 VCC.n14157 3.4105
R43489 VCC.n14110 VCC.n14015 3.4105
R43490 VCC.n14015 VCC.n14009 3.4105
R43491 VCC.n14112 VCC.n14111 3.4105
R43492 VCC.n14132 VCC.n14131 3.4105
R43493 VCC.n14131 VCC.n14130 3.4105
R43494 VCC.n14094 VCC.n14023 3.4105
R43495 VCC.n14023 VCC.n14022 3.4105
R43496 VCC.n14024 VCC.n14017 3.4105
R43497 VCC.n14109 VCC.n14108 3.4105
R43498 VCC.n14108 VCC.n14107 3.4105
R43499 VCC.n14071 VCC.n14070 3.4105
R43500 VCC.n14072 VCC.n14071 3.4105
R43501 VCC.n14093 VCC.n14092 3.4105
R43502 VCC.n14069 VCC.n14068 3.4105
R43503 VCC.n14068 VCC.n14067 3.4105
R43504 VCC.n14718 VCC.n14717 3.4105
R43505 VCC.n14719 VCC.n14718 3.4105
R43506 VCC.n14691 VCC.n14690 3.4105
R43507 VCC.n14716 VCC.n14715 3.4105
R43508 VCC.n14715 VCC.n14714 3.4105
R43509 VCC.n14667 VCC.n14572 3.4105
R43510 VCC.n14572 VCC.n14566 3.4105
R43511 VCC.n14669 VCC.n14668 3.4105
R43512 VCC.n14689 VCC.n14688 3.4105
R43513 VCC.n14688 VCC.n14687 3.4105
R43514 VCC.n14651 VCC.n14580 3.4105
R43515 VCC.n14580 VCC.n14579 3.4105
R43516 VCC.n14581 VCC.n14574 3.4105
R43517 VCC.n14666 VCC.n14665 3.4105
R43518 VCC.n14665 VCC.n14664 3.4105
R43519 VCC.n14628 VCC.n14627 3.4105
R43520 VCC.n14629 VCC.n14628 3.4105
R43521 VCC.n14650 VCC.n14649 3.4105
R43522 VCC.n14626 VCC.n14625 3.4105
R43523 VCC.n14625 VCC.n14624 3.4105
R43524 VCC.n14870 VCC.n14869 3.4105
R43525 VCC.n14869 VCC.n14868 3.4105
R43526 VCC.n14929 VCC.n14928 3.4105
R43527 VCC.n14934 VCC.n14933 3.4105
R43528 VCC.n14933 VCC.n14932 3.4105
R43529 VCC.n14912 VCC.n14911 3.4105
R43530 VCC.n14913 VCC.n14912 3.4105
R43531 VCC.n14910 VCC.n14909 3.4105
R43532 VCC.n14927 VCC.n14926 3.4105
R43533 VCC.n14926 VCC.n14925 3.4105
R43534 VCC.n14899 VCC.n14452 3.4105
R43535 VCC.n14452 VCC.n14451 3.4105
R43536 VCC.n14450 VCC.n14449 3.4105
R43537 VCC.n14907 VCC.n14906 3.4105
R43538 VCC.n14906 VCC.n14445 3.4105
R43539 VCC.n14872 VCC.n14871 3.4105
R43540 VCC.n14872 VCC.n14468 3.4105
R43541 VCC.n14898 VCC.n14897 3.4105
R43542 VCC.n14936 VCC.n14935 3.4105
R43543 VCC.n14936 VCC.n14409 3.4105
R43544 VCC.n14853 VCC.n14852 3.4105
R43545 VCC.n14854 VCC.n14853 3.4105
R43546 VCC.n14817 VCC.n14816 3.4105
R43547 VCC.n14851 VCC.n14850 3.4105
R43548 VCC.n14850 VCC.n14849 3.4105
R43549 VCC.n14787 VCC.n14786 3.4105
R43550 VCC.n14786 VCC.n14785 3.4105
R43551 VCC.n14782 VCC.n14780 3.4105
R43552 VCC.n14815 VCC.n14814 3.4105
R43553 VCC.n14814 VCC.n14813 3.4105
R43554 VCC.n14511 VCC.n14510 3.4105
R43555 VCC.n14758 VCC.n14511 3.4105
R43556 VCC.n14779 VCC.n14508 3.4105
R43557 VCC.n14789 VCC.n14788 3.4105
R43558 VCC.n14789 VCC.n14507 3.4105
R43559 VCC.n14752 VCC.n14522 3.4105
R43560 VCC.n14752 VCC.n14751 3.4105
R43561 VCC.n14756 VCC.n14755 3.4105
R43562 VCC.n14727 VCC.n14726 3.4105
R43563 VCC.n14727 VCC.n14533 3.4105
R43564 VCC.n15497 VCC.n15496 3.4105
R43565 VCC.n15497 VCC.n14963 3.4105
R43566 VCC.n15473 VCC.n15472 3.4105
R43567 VCC.n15495 VCC.n15494 3.4105
R43568 VCC.n15494 VCC.n15493 3.4105
R43569 VCC.n15463 VCC.n14992 3.4105
R43570 VCC.n14992 VCC.n14991 3.4105
R43571 VCC.n15465 VCC.n15464 3.4105
R43572 VCC.n15471 VCC.n15470 3.4105
R43573 VCC.n15470 VCC.n15469 3.4105
R43574 VCC.n15445 VCC.n15444 3.4105
R43575 VCC.n15445 VCC.n15004 3.4105
R43576 VCC.n15441 VCC.n14994 3.4105
R43577 VCC.n15462 VCC.n15461 3.4105
R43578 VCC.n15461 VCC.n15460 3.4105
R43579 VCC.n15423 VCC.n15420 3.4105
R43580 VCC.n15423 VCC.n15422 3.4105
R43581 VCC.n15440 VCC.n15439 3.4105
R43582 VCC.n15419 VCC.n15418 3.4105
R43583 VCC.n15418 VCC.n15417 3.4105
R43584 VCC.n15403 VCC.n15402 3.4105
R43585 VCC.n15404 VCC.n15403 3.4105
R43586 VCC.n15368 VCC.n15367 3.4105
R43587 VCC.n15401 VCC.n15400 3.4105
R43588 VCC.n15400 VCC.n15399 3.4105
R43589 VCC.n15338 VCC.n15337 3.4105
R43590 VCC.n15337 VCC.n15336 3.4105
R43591 VCC.n15333 VCC.n15331 3.4105
R43592 VCC.n15366 VCC.n15365 3.4105
R43593 VCC.n15365 VCC.n15364 3.4105
R43594 VCC.n15062 VCC.n15061 3.4105
R43595 VCC.n15309 VCC.n15062 3.4105
R43596 VCC.n15330 VCC.n15059 3.4105
R43597 VCC.n15340 VCC.n15339 3.4105
R43598 VCC.n15340 VCC.n15058 3.4105
R43599 VCC.n15303 VCC.n15073 3.4105
R43600 VCC.n15303 VCC.n15302 3.4105
R43601 VCC.n15307 VCC.n15306 3.4105
R43602 VCC.n15277 VCC.n15276 3.4105
R43603 VCC.n15277 VCC.n15084 3.4105
R43604 VCC.n15268 VCC.n15267 3.4105
R43605 VCC.n15269 VCC.n15268 3.4105
R43606 VCC.n15241 VCC.n15240 3.4105
R43607 VCC.n15266 VCC.n15265 3.4105
R43608 VCC.n15265 VCC.n15264 3.4105
R43609 VCC.n15217 VCC.n15122 3.4105
R43610 VCC.n15122 VCC.n15116 3.4105
R43611 VCC.n15219 VCC.n15218 3.4105
R43612 VCC.n15239 VCC.n15238 3.4105
R43613 VCC.n15238 VCC.n15237 3.4105
R43614 VCC.n15201 VCC.n15130 3.4105
R43615 VCC.n15130 VCC.n15129 3.4105
R43616 VCC.n15131 VCC.n15124 3.4105
R43617 VCC.n15216 VCC.n15215 3.4105
R43618 VCC.n15215 VCC.n15214 3.4105
R43619 VCC.n15178 VCC.n15177 3.4105
R43620 VCC.n15179 VCC.n15178 3.4105
R43621 VCC.n15200 VCC.n15199 3.4105
R43622 VCC.n15176 VCC.n15175 3.4105
R43623 VCC.n15175 VCC.n15174 3.4105
R43624 VCC.n15825 VCC.n15824 3.4105
R43625 VCC.n15826 VCC.n15825 3.4105
R43626 VCC.n15798 VCC.n15797 3.4105
R43627 VCC.n15823 VCC.n15822 3.4105
R43628 VCC.n15822 VCC.n15821 3.4105
R43629 VCC.n15774 VCC.n15679 3.4105
R43630 VCC.n15679 VCC.n15673 3.4105
R43631 VCC.n15776 VCC.n15775 3.4105
R43632 VCC.n15796 VCC.n15795 3.4105
R43633 VCC.n15795 VCC.n15794 3.4105
R43634 VCC.n15758 VCC.n15687 3.4105
R43635 VCC.n15687 VCC.n15686 3.4105
R43636 VCC.n15688 VCC.n15681 3.4105
R43637 VCC.n15773 VCC.n15772 3.4105
R43638 VCC.n15772 VCC.n15771 3.4105
R43639 VCC.n15735 VCC.n15734 3.4105
R43640 VCC.n15736 VCC.n15735 3.4105
R43641 VCC.n15757 VCC.n15756 3.4105
R43642 VCC.n15733 VCC.n15732 3.4105
R43643 VCC.n15732 VCC.n15731 3.4105
R43644 VCC.n15977 VCC.n15976 3.4105
R43645 VCC.n15976 VCC.n15975 3.4105
R43646 VCC.n16036 VCC.n16035 3.4105
R43647 VCC.n16041 VCC.n16040 3.4105
R43648 VCC.n16040 VCC.n16039 3.4105
R43649 VCC.n16019 VCC.n16018 3.4105
R43650 VCC.n16020 VCC.n16019 3.4105
R43651 VCC.n16017 VCC.n16016 3.4105
R43652 VCC.n16034 VCC.n16033 3.4105
R43653 VCC.n16033 VCC.n16032 3.4105
R43654 VCC.n16006 VCC.n15559 3.4105
R43655 VCC.n15559 VCC.n15558 3.4105
R43656 VCC.n15557 VCC.n15556 3.4105
R43657 VCC.n16014 VCC.n16013 3.4105
R43658 VCC.n16013 VCC.n15552 3.4105
R43659 VCC.n15979 VCC.n15978 3.4105
R43660 VCC.n15979 VCC.n15575 3.4105
R43661 VCC.n16005 VCC.n16004 3.4105
R43662 VCC.n16043 VCC.n16042 3.4105
R43663 VCC.n16043 VCC.n15516 3.4105
R43664 VCC.n15960 VCC.n15959 3.4105
R43665 VCC.n15961 VCC.n15960 3.4105
R43666 VCC.n15924 VCC.n15923 3.4105
R43667 VCC.n15958 VCC.n15957 3.4105
R43668 VCC.n15957 VCC.n15956 3.4105
R43669 VCC.n15894 VCC.n15893 3.4105
R43670 VCC.n15893 VCC.n15892 3.4105
R43671 VCC.n15889 VCC.n15887 3.4105
R43672 VCC.n15922 VCC.n15921 3.4105
R43673 VCC.n15921 VCC.n15920 3.4105
R43674 VCC.n15618 VCC.n15617 3.4105
R43675 VCC.n15865 VCC.n15618 3.4105
R43676 VCC.n15886 VCC.n15615 3.4105
R43677 VCC.n15896 VCC.n15895 3.4105
R43678 VCC.n15896 VCC.n15614 3.4105
R43679 VCC.n15859 VCC.n15629 3.4105
R43680 VCC.n15859 VCC.n15858 3.4105
R43681 VCC.n15863 VCC.n15862 3.4105
R43682 VCC.n15834 VCC.n15833 3.4105
R43683 VCC.n15834 VCC.n15640 3.4105
R43684 VCC.n16604 VCC.n16603 3.4105
R43685 VCC.n16604 VCC.n16070 3.4105
R43686 VCC.n16580 VCC.n16579 3.4105
R43687 VCC.n16602 VCC.n16601 3.4105
R43688 VCC.n16601 VCC.n16600 3.4105
R43689 VCC.n16570 VCC.n16099 3.4105
R43690 VCC.n16099 VCC.n16098 3.4105
R43691 VCC.n16572 VCC.n16571 3.4105
R43692 VCC.n16578 VCC.n16577 3.4105
R43693 VCC.n16577 VCC.n16576 3.4105
R43694 VCC.n16552 VCC.n16551 3.4105
R43695 VCC.n16552 VCC.n16111 3.4105
R43696 VCC.n16548 VCC.n16101 3.4105
R43697 VCC.n16569 VCC.n16568 3.4105
R43698 VCC.n16568 VCC.n16567 3.4105
R43699 VCC.n16530 VCC.n16527 3.4105
R43700 VCC.n16530 VCC.n16529 3.4105
R43701 VCC.n16547 VCC.n16546 3.4105
R43702 VCC.n16526 VCC.n16525 3.4105
R43703 VCC.n16525 VCC.n16524 3.4105
R43704 VCC.n16510 VCC.n16509 3.4105
R43705 VCC.n16511 VCC.n16510 3.4105
R43706 VCC.n16475 VCC.n16474 3.4105
R43707 VCC.n16508 VCC.n16507 3.4105
R43708 VCC.n16507 VCC.n16506 3.4105
R43709 VCC.n16445 VCC.n16444 3.4105
R43710 VCC.n16444 VCC.n16443 3.4105
R43711 VCC.n16440 VCC.n16438 3.4105
R43712 VCC.n16473 VCC.n16472 3.4105
R43713 VCC.n16472 VCC.n16471 3.4105
R43714 VCC.n16169 VCC.n16168 3.4105
R43715 VCC.n16416 VCC.n16169 3.4105
R43716 VCC.n16437 VCC.n16166 3.4105
R43717 VCC.n16447 VCC.n16446 3.4105
R43718 VCC.n16447 VCC.n16165 3.4105
R43719 VCC.n16410 VCC.n16180 3.4105
R43720 VCC.n16410 VCC.n16409 3.4105
R43721 VCC.n16414 VCC.n16413 3.4105
R43722 VCC.n16384 VCC.n16383 3.4105
R43723 VCC.n16384 VCC.n16191 3.4105
R43724 VCC.n16375 VCC.n16374 3.4105
R43725 VCC.n16376 VCC.n16375 3.4105
R43726 VCC.n16348 VCC.n16347 3.4105
R43727 VCC.n16373 VCC.n16372 3.4105
R43728 VCC.n16372 VCC.n16371 3.4105
R43729 VCC.n16324 VCC.n16229 3.4105
R43730 VCC.n16229 VCC.n16223 3.4105
R43731 VCC.n16326 VCC.n16325 3.4105
R43732 VCC.n16346 VCC.n16345 3.4105
R43733 VCC.n16345 VCC.n16344 3.4105
R43734 VCC.n16308 VCC.n16237 3.4105
R43735 VCC.n16237 VCC.n16236 3.4105
R43736 VCC.n16238 VCC.n16231 3.4105
R43737 VCC.n16323 VCC.n16322 3.4105
R43738 VCC.n16322 VCC.n16321 3.4105
R43739 VCC.n16285 VCC.n16284 3.4105
R43740 VCC.n16286 VCC.n16285 3.4105
R43741 VCC.n16307 VCC.n16306 3.4105
R43742 VCC.n16283 VCC.n16282 3.4105
R43743 VCC.n16282 VCC.n16281 3.4105
R43744 VCC.n16932 VCC.n16931 3.4105
R43745 VCC.n16933 VCC.n16932 3.4105
R43746 VCC.n16905 VCC.n16904 3.4105
R43747 VCC.n16930 VCC.n16929 3.4105
R43748 VCC.n16929 VCC.n16928 3.4105
R43749 VCC.n16881 VCC.n16786 3.4105
R43750 VCC.n16786 VCC.n16780 3.4105
R43751 VCC.n16883 VCC.n16882 3.4105
R43752 VCC.n16903 VCC.n16902 3.4105
R43753 VCC.n16902 VCC.n16901 3.4105
R43754 VCC.n16865 VCC.n16794 3.4105
R43755 VCC.n16794 VCC.n16793 3.4105
R43756 VCC.n16795 VCC.n16788 3.4105
R43757 VCC.n16880 VCC.n16879 3.4105
R43758 VCC.n16879 VCC.n16878 3.4105
R43759 VCC.n16842 VCC.n16841 3.4105
R43760 VCC.n16843 VCC.n16842 3.4105
R43761 VCC.n16864 VCC.n16863 3.4105
R43762 VCC.n16840 VCC.n16839 3.4105
R43763 VCC.n16839 VCC.n16838 3.4105
R43764 VCC.n17084 VCC.n17083 3.4105
R43765 VCC.n17083 VCC.n17082 3.4105
R43766 VCC.n17143 VCC.n17142 3.4105
R43767 VCC.n17148 VCC.n17147 3.4105
R43768 VCC.n17147 VCC.n17146 3.4105
R43769 VCC.n17126 VCC.n17125 3.4105
R43770 VCC.n17127 VCC.n17126 3.4105
R43771 VCC.n17124 VCC.n17123 3.4105
R43772 VCC.n17141 VCC.n17140 3.4105
R43773 VCC.n17140 VCC.n17139 3.4105
R43774 VCC.n17113 VCC.n16666 3.4105
R43775 VCC.n16666 VCC.n16665 3.4105
R43776 VCC.n16664 VCC.n16663 3.4105
R43777 VCC.n17121 VCC.n17120 3.4105
R43778 VCC.n17120 VCC.n16659 3.4105
R43779 VCC.n17086 VCC.n17085 3.4105
R43780 VCC.n17086 VCC.n16682 3.4105
R43781 VCC.n17112 VCC.n17111 3.4105
R43782 VCC.n17150 VCC.n17149 3.4105
R43783 VCC.n17150 VCC.n16623 3.4105
R43784 VCC.n17067 VCC.n17066 3.4105
R43785 VCC.n17068 VCC.n17067 3.4105
R43786 VCC.n17031 VCC.n17030 3.4105
R43787 VCC.n17065 VCC.n17064 3.4105
R43788 VCC.n17064 VCC.n17063 3.4105
R43789 VCC.n17001 VCC.n17000 3.4105
R43790 VCC.n17000 VCC.n16999 3.4105
R43791 VCC.n16996 VCC.n16994 3.4105
R43792 VCC.n17029 VCC.n17028 3.4105
R43793 VCC.n17028 VCC.n17027 3.4105
R43794 VCC.n16725 VCC.n16724 3.4105
R43795 VCC.n16972 VCC.n16725 3.4105
R43796 VCC.n16993 VCC.n16722 3.4105
R43797 VCC.n17003 VCC.n17002 3.4105
R43798 VCC.n17003 VCC.n16721 3.4105
R43799 VCC.n16966 VCC.n16736 3.4105
R43800 VCC.n16966 VCC.n16965 3.4105
R43801 VCC.n16970 VCC.n16969 3.4105
R43802 VCC.n16941 VCC.n16940 3.4105
R43803 VCC.n16941 VCC.n16747 3.4105
R43804 VCC.n17524 VCC.n17523 3.4105
R43805 VCC.n17524 VCC.n17177 3.4105
R43806 VCC.n17500 VCC.n17499 3.4105
R43807 VCC.n17522 VCC.n17521 3.4105
R43808 VCC.n17521 VCC.n17520 3.4105
R43809 VCC.n17490 VCC.n17206 3.4105
R43810 VCC.n17206 VCC.n17205 3.4105
R43811 VCC.n17492 VCC.n17491 3.4105
R43812 VCC.n17498 VCC.n17497 3.4105
R43813 VCC.n17497 VCC.n17496 3.4105
R43814 VCC.n17472 VCC.n17471 3.4105
R43815 VCC.n17472 VCC.n17218 3.4105
R43816 VCC.n17468 VCC.n17208 3.4105
R43817 VCC.n17489 VCC.n17488 3.4105
R43818 VCC.n17488 VCC.n17487 3.4105
R43819 VCC.n17450 VCC.n17447 3.4105
R43820 VCC.n17450 VCC.n17449 3.4105
R43821 VCC.n17467 VCC.n17466 3.4105
R43822 VCC.n17446 VCC.n17445 3.4105
R43823 VCC.n17445 VCC.n17444 3.4105
R43824 VCC.n17430 VCC.n17429 3.4105
R43825 VCC.n17431 VCC.n17430 3.4105
R43826 VCC.n17395 VCC.n17394 3.4105
R43827 VCC.n17428 VCC.n17427 3.4105
R43828 VCC.n17427 VCC.n17426 3.4105
R43829 VCC.n17365 VCC.n17364 3.4105
R43830 VCC.n17364 VCC.n17363 3.4105
R43831 VCC.n17360 VCC.n17358 3.4105
R43832 VCC.n17393 VCC.n17392 3.4105
R43833 VCC.n17392 VCC.n17391 3.4105
R43834 VCC.n17276 VCC.n17275 3.4105
R43835 VCC.n17336 VCC.n17276 3.4105
R43836 VCC.n17357 VCC.n17273 3.4105
R43837 VCC.n17367 VCC.n17366 3.4105
R43838 VCC.n17367 VCC.n17272 3.4105
R43839 VCC.n17330 VCC.n17287 3.4105
R43840 VCC.n17330 VCC.n17329 3.4105
R43841 VCC.n17334 VCC.n17333 3.4105
R43842 VCC.n17304 VCC.n17303 3.4105
R43843 VCC.n17304 VCC.n17298 3.4105
R43844 VCC.n421 VCC.n57 3.29193
R43845 VCC.n476 VCC.n475 3.29193
R43846 VCC.n515 VCC.n20 3.29193
R43847 VCC.n973 VCC.n609 3.29193
R43848 VCC.n1028 VCC.n1027 3.29193
R43849 VCC.n1067 VCC.n572 3.29193
R43850 VCC.n1531 VCC.n1165 3.29193
R43851 VCC.n1594 VCC.n1159 3.29193
R43852 VCC.n1140 VCC.n1116 3.29193
R43853 VCC.n2082 VCC.n1718 3.29193
R43854 VCC.n2137 VCC.n2136 3.29193
R43855 VCC.n2176 VCC.n1681 3.29193
R43856 VCC.n2640 VCC.n2274 3.29193
R43857 VCC.n2703 VCC.n2268 3.29193
R43858 VCC.n2249 VCC.n2225 3.29193
R43859 VCC.n3191 VCC.n2827 3.29193
R43860 VCC.n3246 VCC.n3245 3.29193
R43861 VCC.n3285 VCC.n2790 3.29193
R43862 VCC.n3749 VCC.n3383 3.29193
R43863 VCC.n3812 VCC.n3377 3.29193
R43864 VCC.n3358 VCC.n3334 3.29193
R43865 VCC.n4300 VCC.n3936 3.29193
R43866 VCC.n4355 VCC.n4354 3.29193
R43867 VCC.n4394 VCC.n3899 3.29193
R43868 VCC.n4858 VCC.n4492 3.29193
R43869 VCC.n4921 VCC.n4486 3.29193
R43870 VCC.n4467 VCC.n4443 3.29193
R43871 VCC.n5409 VCC.n5045 3.29193
R43872 VCC.n5464 VCC.n5463 3.29193
R43873 VCC.n5503 VCC.n5008 3.29193
R43874 VCC.n5967 VCC.n5601 3.29193
R43875 VCC.n6030 VCC.n5595 3.29193
R43876 VCC.n5576 VCC.n5552 3.29193
R43877 VCC.n6518 VCC.n6154 3.29193
R43878 VCC.n6573 VCC.n6572 3.29193
R43879 VCC.n6612 VCC.n6117 3.29193
R43880 VCC.n7076 VCC.n6710 3.29193
R43881 VCC.n7139 VCC.n6704 3.29193
R43882 VCC.n6685 VCC.n6661 3.29193
R43883 VCC.n7627 VCC.n7263 3.29193
R43884 VCC.n7682 VCC.n7681 3.29193
R43885 VCC.n7721 VCC.n7226 3.29193
R43886 VCC.n8185 VCC.n7819 3.29193
R43887 VCC.n8248 VCC.n7813 3.29193
R43888 VCC.n7794 VCC.n7770 3.29193
R43889 VCC.n8736 VCC.n8372 3.29193
R43890 VCC.n8791 VCC.n8790 3.29193
R43891 VCC.n8830 VCC.n8335 3.29193
R43892 VCC.n9294 VCC.n8928 3.29193
R43893 VCC.n9357 VCC.n8922 3.29193
R43894 VCC.n8903 VCC.n8879 3.29193
R43895 VCC.n9845 VCC.n9481 3.29193
R43896 VCC.n9900 VCC.n9899 3.29193
R43897 VCC.n9939 VCC.n9444 3.29193
R43898 VCC.n10402 VCC.n10036 3.29193
R43899 VCC.n10465 VCC.n10030 3.29193
R43900 VCC.n10011 VCC.n9987 3.29193
R43901 VCC.n10952 VCC.n10588 3.29193
R43902 VCC.n11007 VCC.n11006 3.29193
R43903 VCC.n11046 VCC.n10551 3.29193
R43904 VCC.n11509 VCC.n11143 3.29193
R43905 VCC.n11572 VCC.n11137 3.29193
R43906 VCC.n11118 VCC.n11094 3.29193
R43907 VCC.n12059 VCC.n11695 3.29193
R43908 VCC.n12114 VCC.n12113 3.29193
R43909 VCC.n12153 VCC.n11658 3.29193
R43910 VCC.n12616 VCC.n12250 3.29193
R43911 VCC.n12679 VCC.n12244 3.29193
R43912 VCC.n12225 VCC.n12201 3.29193
R43913 VCC.n13166 VCC.n12802 3.29193
R43914 VCC.n13221 VCC.n13220 3.29193
R43915 VCC.n13260 VCC.n12765 3.29193
R43916 VCC.n13723 VCC.n13357 3.29193
R43917 VCC.n13786 VCC.n13351 3.29193
R43918 VCC.n13332 VCC.n13308 3.29193
R43919 VCC.n14273 VCC.n13909 3.29193
R43920 VCC.n14328 VCC.n14327 3.29193
R43921 VCC.n14367 VCC.n13872 3.29193
R43922 VCC.n14830 VCC.n14464 3.29193
R43923 VCC.n14893 VCC.n14458 3.29193
R43924 VCC.n14439 VCC.n14415 3.29193
R43925 VCC.n15380 VCC.n15016 3.29193
R43926 VCC.n15435 VCC.n15434 3.29193
R43927 VCC.n15474 VCC.n14979 3.29193
R43928 VCC.n15937 VCC.n15571 3.29193
R43929 VCC.n16000 VCC.n15565 3.29193
R43930 VCC.n15546 VCC.n15522 3.29193
R43931 VCC.n16487 VCC.n16123 3.29193
R43932 VCC.n16542 VCC.n16541 3.29193
R43933 VCC.n16581 VCC.n16086 3.29193
R43934 VCC.n17044 VCC.n16678 3.29193
R43935 VCC.n17107 VCC.n16672 3.29193
R43936 VCC.n16653 VCC.n16629 3.29193
R43937 VCC.n17407 VCC.n17230 3.29193
R43938 VCC.n17462 VCC.n17461 3.29193
R43939 VCC.n17501 VCC.n17193 3.29193
R43940 VCC.n469 VCC.n55 3.25764
R43941 VCC.n528 VCC.n6 3.25764
R43942 VCC.n1021 VCC.n607 3.25764
R43943 VCC.n1080 VCC.n560 3.25764
R43944 VCC.n1579 VCC.n1164 3.25764
R43945 VCC.n1650 VCC.n1113 3.25764
R43946 VCC.n2130 VCC.n1716 3.25764
R43947 VCC.n2189 VCC.n1669 3.25764
R43948 VCC.n2688 VCC.n2273 3.25764
R43949 VCC.n2759 VCC.n2222 3.25764
R43950 VCC.n3239 VCC.n2825 3.25764
R43951 VCC.n3298 VCC.n2778 3.25764
R43952 VCC.n3797 VCC.n3382 3.25764
R43953 VCC.n3868 VCC.n3331 3.25764
R43954 VCC.n4348 VCC.n3934 3.25764
R43955 VCC.n4407 VCC.n3887 3.25764
R43956 VCC.n4906 VCC.n4491 3.25764
R43957 VCC.n4977 VCC.n4440 3.25764
R43958 VCC.n5457 VCC.n5043 3.25764
R43959 VCC.n5516 VCC.n4996 3.25764
R43960 VCC.n6015 VCC.n5600 3.25764
R43961 VCC.n6086 VCC.n5549 3.25764
R43962 VCC.n6566 VCC.n6152 3.25764
R43963 VCC.n6625 VCC.n6105 3.25764
R43964 VCC.n7124 VCC.n6709 3.25764
R43965 VCC.n7195 VCC.n6658 3.25764
R43966 VCC.n7675 VCC.n7261 3.25764
R43967 VCC.n7734 VCC.n7214 3.25764
R43968 VCC.n8233 VCC.n7818 3.25764
R43969 VCC.n8304 VCC.n7767 3.25764
R43970 VCC.n8784 VCC.n8370 3.25764
R43971 VCC.n8843 VCC.n8323 3.25764
R43972 VCC.n9342 VCC.n8927 3.25764
R43973 VCC.n9413 VCC.n8876 3.25764
R43974 VCC.n9893 VCC.n9479 3.25764
R43975 VCC.n9952 VCC.n9432 3.25764
R43976 VCC.n10450 VCC.n10035 3.25764
R43977 VCC.n10521 VCC.n9984 3.25764
R43978 VCC.n11000 VCC.n10586 3.25764
R43979 VCC.n11059 VCC.n10539 3.25764
R43980 VCC.n11557 VCC.n11142 3.25764
R43981 VCC.n11628 VCC.n11091 3.25764
R43982 VCC.n12107 VCC.n11693 3.25764
R43983 VCC.n12166 VCC.n11646 3.25764
R43984 VCC.n12664 VCC.n12249 3.25764
R43985 VCC.n12735 VCC.n12198 3.25764
R43986 VCC.n13214 VCC.n12800 3.25764
R43987 VCC.n13273 VCC.n12753 3.25764
R43988 VCC.n13771 VCC.n13356 3.25764
R43989 VCC.n13842 VCC.n13305 3.25764
R43990 VCC.n14321 VCC.n13907 3.25764
R43991 VCC.n14380 VCC.n13860 3.25764
R43992 VCC.n14878 VCC.n14463 3.25764
R43993 VCC.n14949 VCC.n14412 3.25764
R43994 VCC.n15428 VCC.n15014 3.25764
R43995 VCC.n15487 VCC.n14967 3.25764
R43996 VCC.n15985 VCC.n15570 3.25764
R43997 VCC.n16056 VCC.n15519 3.25764
R43998 VCC.n16535 VCC.n16121 3.25764
R43999 VCC.n16594 VCC.n16074 3.25764
R44000 VCC.n17092 VCC.n16677 3.25764
R44001 VCC.n17163 VCC.n16626 3.25764
R44002 VCC.n17455 VCC.n17228 3.25764
R44003 VCC.n17514 VCC.n17181 3.25764
R44004 VCC.n545 VCC.n544 3.2005
R44005 VCC.n1099 VCC.n1098 3.2005
R44006 VCC.n1124 VCC.n1112 3.2005
R44007 VCC.n2208 VCC.n2207 3.2005
R44008 VCC.n2233 VCC.n2221 3.2005
R44009 VCC.n3317 VCC.n3316 3.2005
R44010 VCC.n3342 VCC.n3330 3.2005
R44011 VCC.n4426 VCC.n4425 3.2005
R44012 VCC.n4451 VCC.n4439 3.2005
R44013 VCC.n5535 VCC.n5534 3.2005
R44014 VCC.n5560 VCC.n5548 3.2005
R44015 VCC.n6644 VCC.n6643 3.2005
R44016 VCC.n6669 VCC.n6657 3.2005
R44017 VCC.n7753 VCC.n7752 3.2005
R44018 VCC.n7778 VCC.n7766 3.2005
R44019 VCC.n8862 VCC.n8861 3.2005
R44020 VCC.n8887 VCC.n8875 3.2005
R44021 VCC.n9971 VCC.n9970 3.2005
R44022 VCC.n9995 VCC.n9983 3.2005
R44023 VCC.n11078 VCC.n11077 3.2005
R44024 VCC.n11102 VCC.n11090 3.2005
R44025 VCC.n12185 VCC.n12184 3.2005
R44026 VCC.n12209 VCC.n12197 3.2005
R44027 VCC.n13292 VCC.n13291 3.2005
R44028 VCC.n13316 VCC.n13304 3.2005
R44029 VCC.n14399 VCC.n14398 3.2005
R44030 VCC.n14423 VCC.n14411 3.2005
R44031 VCC.n15506 VCC.n15505 3.2005
R44032 VCC.n15530 VCC.n15518 3.2005
R44033 VCC.n16613 VCC.n16612 3.2005
R44034 VCC.n16637 VCC.n16625 3.2005
R44035 VCC.n17533 VCC.n17532 3.2005
R44036 VCC.n500 VCC.n499 3.03311
R44037 VCC.n468 VCC.n467 3.03311
R44038 VCC.n1020 VCC.n1019 3.03311
R44039 VCC.n1052 VCC.n1051 3.03311
R44040 VCC.n1616 VCC.n1615 3.03311
R44041 VCC.n1577 VCC.n1576 3.03311
R44042 VCC.n2129 VCC.n2128 3.03311
R44043 VCC.n2161 VCC.n2160 3.03311
R44044 VCC.n2725 VCC.n2724 3.03311
R44045 VCC.n2686 VCC.n2685 3.03311
R44046 VCC.n3238 VCC.n3237 3.03311
R44047 VCC.n3270 VCC.n3269 3.03311
R44048 VCC.n3834 VCC.n3833 3.03311
R44049 VCC.n3795 VCC.n3794 3.03311
R44050 VCC.n4347 VCC.n4346 3.03311
R44051 VCC.n4379 VCC.n4378 3.03311
R44052 VCC.n4943 VCC.n4942 3.03311
R44053 VCC.n4904 VCC.n4903 3.03311
R44054 VCC.n5456 VCC.n5455 3.03311
R44055 VCC.n5488 VCC.n5487 3.03311
R44056 VCC.n6052 VCC.n6051 3.03311
R44057 VCC.n6013 VCC.n6012 3.03311
R44058 VCC.n6565 VCC.n6564 3.03311
R44059 VCC.n6597 VCC.n6596 3.03311
R44060 VCC.n7161 VCC.n7160 3.03311
R44061 VCC.n7122 VCC.n7121 3.03311
R44062 VCC.n7674 VCC.n7673 3.03311
R44063 VCC.n7706 VCC.n7705 3.03311
R44064 VCC.n8270 VCC.n8269 3.03311
R44065 VCC.n8231 VCC.n8230 3.03311
R44066 VCC.n8783 VCC.n8782 3.03311
R44067 VCC.n8815 VCC.n8814 3.03311
R44068 VCC.n9379 VCC.n9378 3.03311
R44069 VCC.n9340 VCC.n9339 3.03311
R44070 VCC.n9892 VCC.n9891 3.03311
R44071 VCC.n9924 VCC.n9923 3.03311
R44072 VCC.n10487 VCC.n10486 3.03311
R44073 VCC.n10448 VCC.n10447 3.03311
R44074 VCC.n10999 VCC.n10998 3.03311
R44075 VCC.n11031 VCC.n11030 3.03311
R44076 VCC.n11594 VCC.n11593 3.03311
R44077 VCC.n11555 VCC.n11554 3.03311
R44078 VCC.n12106 VCC.n12105 3.03311
R44079 VCC.n12138 VCC.n12137 3.03311
R44080 VCC.n12701 VCC.n12700 3.03311
R44081 VCC.n12662 VCC.n12661 3.03311
R44082 VCC.n13213 VCC.n13212 3.03311
R44083 VCC.n13245 VCC.n13244 3.03311
R44084 VCC.n13808 VCC.n13807 3.03311
R44085 VCC.n13769 VCC.n13768 3.03311
R44086 VCC.n14320 VCC.n14319 3.03311
R44087 VCC.n14352 VCC.n14351 3.03311
R44088 VCC.n14915 VCC.n14914 3.03311
R44089 VCC.n14876 VCC.n14875 3.03311
R44090 VCC.n15427 VCC.n15426 3.03311
R44091 VCC.n15459 VCC.n15458 3.03311
R44092 VCC.n16022 VCC.n16021 3.03311
R44093 VCC.n15983 VCC.n15982 3.03311
R44094 VCC.n16534 VCC.n16533 3.03311
R44095 VCC.n16566 VCC.n16565 3.03311
R44096 VCC.n17129 VCC.n17128 3.03311
R44097 VCC.n17090 VCC.n17089 3.03311
R44098 VCC.n17454 VCC.n17453 3.03311
R44099 VCC.n17486 VCC.n17485 3.03311
R44100 VCC.n225 VCC.n182 2.8505
R44101 VCC.n292 VCC.n140 2.8505
R44102 VCC.n338 VCC.n119 2.8505
R44103 VCC.n416 VCC.n80 2.8505
R44104 VCC.n777 VCC.n734 2.8505
R44105 VCC.n844 VCC.n692 2.8505
R44106 VCC.n890 VCC.n671 2.8505
R44107 VCC.n968 VCC.n632 2.8505
R44108 VCC.n1447 VCC.n1228 2.8505
R44109 VCC.n1525 VCC.n1189 2.8505
R44110 VCC.n1335 VCC.n1292 2.8505
R44111 VCC.n1402 VCC.n1250 2.8505
R44112 VCC.n1886 VCC.n1843 2.8505
R44113 VCC.n1953 VCC.n1801 2.8505
R44114 VCC.n1999 VCC.n1780 2.8505
R44115 VCC.n2077 VCC.n1741 2.8505
R44116 VCC.n2556 VCC.n2337 2.8505
R44117 VCC.n2634 VCC.n2298 2.8505
R44118 VCC.n2444 VCC.n2401 2.8505
R44119 VCC.n2511 VCC.n2359 2.8505
R44120 VCC.n2995 VCC.n2952 2.8505
R44121 VCC.n3062 VCC.n2910 2.8505
R44122 VCC.n3108 VCC.n2889 2.8505
R44123 VCC.n3186 VCC.n2850 2.8505
R44124 VCC.n3665 VCC.n3446 2.8505
R44125 VCC.n3743 VCC.n3407 2.8505
R44126 VCC.n3553 VCC.n3510 2.8505
R44127 VCC.n3620 VCC.n3468 2.8505
R44128 VCC.n4104 VCC.n4061 2.8505
R44129 VCC.n4171 VCC.n4019 2.8505
R44130 VCC.n4217 VCC.n3998 2.8505
R44131 VCC.n4295 VCC.n3959 2.8505
R44132 VCC.n4774 VCC.n4555 2.8505
R44133 VCC.n4852 VCC.n4516 2.8505
R44134 VCC.n4662 VCC.n4619 2.8505
R44135 VCC.n4729 VCC.n4577 2.8505
R44136 VCC.n5213 VCC.n5170 2.8505
R44137 VCC.n5280 VCC.n5128 2.8505
R44138 VCC.n5326 VCC.n5107 2.8505
R44139 VCC.n5404 VCC.n5068 2.8505
R44140 VCC.n5883 VCC.n5664 2.8505
R44141 VCC.n5961 VCC.n5625 2.8505
R44142 VCC.n5771 VCC.n5728 2.8505
R44143 VCC.n5838 VCC.n5686 2.8505
R44144 VCC.n6322 VCC.n6279 2.8505
R44145 VCC.n6389 VCC.n6237 2.8505
R44146 VCC.n6435 VCC.n6216 2.8505
R44147 VCC.n6513 VCC.n6177 2.8505
R44148 VCC.n6992 VCC.n6773 2.8505
R44149 VCC.n7070 VCC.n6734 2.8505
R44150 VCC.n6880 VCC.n6837 2.8505
R44151 VCC.n6947 VCC.n6795 2.8505
R44152 VCC.n7431 VCC.n7388 2.8505
R44153 VCC.n7498 VCC.n7346 2.8505
R44154 VCC.n7544 VCC.n7325 2.8505
R44155 VCC.n7622 VCC.n7286 2.8505
R44156 VCC.n8101 VCC.n7882 2.8505
R44157 VCC.n8179 VCC.n7843 2.8505
R44158 VCC.n7989 VCC.n7946 2.8505
R44159 VCC.n8056 VCC.n7904 2.8505
R44160 VCC.n8653 VCC.n8434 2.8505
R44161 VCC.n8731 VCC.n8395 2.8505
R44162 VCC.n8540 VCC.n8497 2.8505
R44163 VCC.n8607 VCC.n8455 2.8505
R44164 VCC.n9210 VCC.n8991 2.8505
R44165 VCC.n9288 VCC.n8952 2.8505
R44166 VCC.n9098 VCC.n9055 2.8505
R44167 VCC.n9165 VCC.n9013 2.8505
R44168 VCC.n9649 VCC.n9606 2.8505
R44169 VCC.n9716 VCC.n9564 2.8505
R44170 VCC.n9762 VCC.n9543 2.8505
R44171 VCC.n9840 VCC.n9504 2.8505
R44172 VCC.n10318 VCC.n10099 2.8505
R44173 VCC.n10396 VCC.n10060 2.8505
R44174 VCC.n10206 VCC.n10163 2.8505
R44175 VCC.n10273 VCC.n10121 2.8505
R44176 VCC.n10756 VCC.n10713 2.8505
R44177 VCC.n10823 VCC.n10671 2.8505
R44178 VCC.n10869 VCC.n10650 2.8505
R44179 VCC.n10947 VCC.n10611 2.8505
R44180 VCC.n11425 VCC.n11206 2.8505
R44181 VCC.n11503 VCC.n11167 2.8505
R44182 VCC.n11313 VCC.n11270 2.8505
R44183 VCC.n11380 VCC.n11228 2.8505
R44184 VCC.n11863 VCC.n11820 2.8505
R44185 VCC.n11930 VCC.n11778 2.8505
R44186 VCC.n11976 VCC.n11757 2.8505
R44187 VCC.n12054 VCC.n11718 2.8505
R44188 VCC.n12532 VCC.n12313 2.8505
R44189 VCC.n12610 VCC.n12274 2.8505
R44190 VCC.n12420 VCC.n12377 2.8505
R44191 VCC.n12487 VCC.n12335 2.8505
R44192 VCC.n12970 VCC.n12927 2.8505
R44193 VCC.n13037 VCC.n12885 2.8505
R44194 VCC.n13083 VCC.n12864 2.8505
R44195 VCC.n13161 VCC.n12825 2.8505
R44196 VCC.n13639 VCC.n13420 2.8505
R44197 VCC.n13717 VCC.n13381 2.8505
R44198 VCC.n13527 VCC.n13484 2.8505
R44199 VCC.n13594 VCC.n13442 2.8505
R44200 VCC.n14077 VCC.n14034 2.8505
R44201 VCC.n14144 VCC.n13992 2.8505
R44202 VCC.n14190 VCC.n13971 2.8505
R44203 VCC.n14268 VCC.n13932 2.8505
R44204 VCC.n14746 VCC.n14527 2.8505
R44205 VCC.n14824 VCC.n14488 2.8505
R44206 VCC.n14634 VCC.n14591 2.8505
R44207 VCC.n14701 VCC.n14549 2.8505
R44208 VCC.n15184 VCC.n15141 2.8505
R44209 VCC.n15251 VCC.n15099 2.8505
R44210 VCC.n15297 VCC.n15078 2.8505
R44211 VCC.n15375 VCC.n15039 2.8505
R44212 VCC.n15853 VCC.n15634 2.8505
R44213 VCC.n15931 VCC.n15595 2.8505
R44214 VCC.n15741 VCC.n15698 2.8505
R44215 VCC.n15808 VCC.n15656 2.8505
R44216 VCC.n16291 VCC.n16248 2.8505
R44217 VCC.n16358 VCC.n16206 2.8505
R44218 VCC.n16404 VCC.n16185 2.8505
R44219 VCC.n16482 VCC.n16146 2.8505
R44220 VCC.n16960 VCC.n16741 2.8505
R44221 VCC.n17038 VCC.n16702 2.8505
R44222 VCC.n16848 VCC.n16805 2.8505
R44223 VCC.n16915 VCC.n16763 2.8505
R44224 VCC.n17324 VCC.n17292 2.8505
R44225 VCC.n17402 VCC.n17253 2.8505
R44226 VCC.n272 VCC.n271 2.5605
R44227 VCC.n399 VCC.n398 2.5605
R44228 VCC.n824 VCC.n823 2.5605
R44229 VCC.n951 VCC.n950 2.5605
R44230 VCC.n1508 VCC.n1507 2.5605
R44231 VCC.n1382 VCC.n1381 2.5605
R44232 VCC.n1933 VCC.n1932 2.5605
R44233 VCC.n2060 VCC.n2059 2.5605
R44234 VCC.n2617 VCC.n2616 2.5605
R44235 VCC.n2491 VCC.n2490 2.5605
R44236 VCC.n3042 VCC.n3041 2.5605
R44237 VCC.n3169 VCC.n3168 2.5605
R44238 VCC.n3726 VCC.n3725 2.5605
R44239 VCC.n3600 VCC.n3599 2.5605
R44240 VCC.n4151 VCC.n4150 2.5605
R44241 VCC.n4278 VCC.n4277 2.5605
R44242 VCC.n4835 VCC.n4834 2.5605
R44243 VCC.n4709 VCC.n4708 2.5605
R44244 VCC.n5260 VCC.n5259 2.5605
R44245 VCC.n5387 VCC.n5386 2.5605
R44246 VCC.n5944 VCC.n5943 2.5605
R44247 VCC.n5818 VCC.n5817 2.5605
R44248 VCC.n6369 VCC.n6368 2.5605
R44249 VCC.n6496 VCC.n6495 2.5605
R44250 VCC.n7053 VCC.n7052 2.5605
R44251 VCC.n6927 VCC.n6926 2.5605
R44252 VCC.n7478 VCC.n7477 2.5605
R44253 VCC.n7605 VCC.n7604 2.5605
R44254 VCC.n8162 VCC.n8161 2.5605
R44255 VCC.n8036 VCC.n8035 2.5605
R44256 VCC.n8714 VCC.n8713 2.5605
R44257 VCC.n8587 VCC.n8586 2.5605
R44258 VCC.n9271 VCC.n9270 2.5605
R44259 VCC.n9145 VCC.n9144 2.5605
R44260 VCC.n9696 VCC.n9695 2.5605
R44261 VCC.n9823 VCC.n9822 2.5605
R44262 VCC.n10379 VCC.n10378 2.5605
R44263 VCC.n10253 VCC.n10252 2.5605
R44264 VCC.n10803 VCC.n10802 2.5605
R44265 VCC.n10930 VCC.n10929 2.5605
R44266 VCC.n11486 VCC.n11485 2.5605
R44267 VCC.n11360 VCC.n11359 2.5605
R44268 VCC.n11910 VCC.n11909 2.5605
R44269 VCC.n12037 VCC.n12036 2.5605
R44270 VCC.n12593 VCC.n12592 2.5605
R44271 VCC.n12467 VCC.n12466 2.5605
R44272 VCC.n13017 VCC.n13016 2.5605
R44273 VCC.n13144 VCC.n13143 2.5605
R44274 VCC.n13700 VCC.n13699 2.5605
R44275 VCC.n13574 VCC.n13573 2.5605
R44276 VCC.n14124 VCC.n14123 2.5605
R44277 VCC.n14251 VCC.n14250 2.5605
R44278 VCC.n14807 VCC.n14806 2.5605
R44279 VCC.n14681 VCC.n14680 2.5605
R44280 VCC.n15231 VCC.n15230 2.5605
R44281 VCC.n15358 VCC.n15357 2.5605
R44282 VCC.n15914 VCC.n15913 2.5605
R44283 VCC.n15788 VCC.n15787 2.5605
R44284 VCC.n16338 VCC.n16337 2.5605
R44285 VCC.n16465 VCC.n16464 2.5605
R44286 VCC.n17021 VCC.n17020 2.5605
R44287 VCC.n16895 VCC.n16894 2.5605
R44288 VCC.n17385 VCC.n17384 2.5605
R44289 VCC.n232 VCC.n231 2.46907
R44290 VCC.n358 VCC.n357 2.46907
R44291 VCC.n784 VCC.n783 2.46907
R44292 VCC.n910 VCC.n909 2.46907
R44293 VCC.n1467 VCC.n1466 2.46907
R44294 VCC.n1342 VCC.n1341 2.46907
R44295 VCC.n1893 VCC.n1892 2.46907
R44296 VCC.n2019 VCC.n2018 2.46907
R44297 VCC.n2576 VCC.n2575 2.46907
R44298 VCC.n2451 VCC.n2450 2.46907
R44299 VCC.n3002 VCC.n3001 2.46907
R44300 VCC.n3128 VCC.n3127 2.46907
R44301 VCC.n3685 VCC.n3684 2.46907
R44302 VCC.n3560 VCC.n3559 2.46907
R44303 VCC.n4111 VCC.n4110 2.46907
R44304 VCC.n4237 VCC.n4236 2.46907
R44305 VCC.n4794 VCC.n4793 2.46907
R44306 VCC.n4669 VCC.n4668 2.46907
R44307 VCC.n5220 VCC.n5219 2.46907
R44308 VCC.n5346 VCC.n5345 2.46907
R44309 VCC.n5903 VCC.n5902 2.46907
R44310 VCC.n5778 VCC.n5777 2.46907
R44311 VCC.n6329 VCC.n6328 2.46907
R44312 VCC.n6455 VCC.n6454 2.46907
R44313 VCC.n7012 VCC.n7011 2.46907
R44314 VCC.n6887 VCC.n6886 2.46907
R44315 VCC.n7438 VCC.n7437 2.46907
R44316 VCC.n7564 VCC.n7563 2.46907
R44317 VCC.n8121 VCC.n8120 2.46907
R44318 VCC.n7996 VCC.n7995 2.46907
R44319 VCC.n8673 VCC.n8672 2.46907
R44320 VCC.n8547 VCC.n8546 2.46907
R44321 VCC.n9230 VCC.n9229 2.46907
R44322 VCC.n9105 VCC.n9104 2.46907
R44323 VCC.n9656 VCC.n9655 2.46907
R44324 VCC.n9782 VCC.n9781 2.46907
R44325 VCC.n10338 VCC.n10337 2.46907
R44326 VCC.n10213 VCC.n10212 2.46907
R44327 VCC.n10763 VCC.n10762 2.46907
R44328 VCC.n10889 VCC.n10888 2.46907
R44329 VCC.n11445 VCC.n11444 2.46907
R44330 VCC.n11320 VCC.n11319 2.46907
R44331 VCC.n11870 VCC.n11869 2.46907
R44332 VCC.n11996 VCC.n11995 2.46907
R44333 VCC.n12552 VCC.n12551 2.46907
R44334 VCC.n12427 VCC.n12426 2.46907
R44335 VCC.n12977 VCC.n12976 2.46907
R44336 VCC.n13103 VCC.n13102 2.46907
R44337 VCC.n13659 VCC.n13658 2.46907
R44338 VCC.n13534 VCC.n13533 2.46907
R44339 VCC.n14084 VCC.n14083 2.46907
R44340 VCC.n14210 VCC.n14209 2.46907
R44341 VCC.n14766 VCC.n14765 2.46907
R44342 VCC.n14641 VCC.n14640 2.46907
R44343 VCC.n15191 VCC.n15190 2.46907
R44344 VCC.n15317 VCC.n15316 2.46907
R44345 VCC.n15873 VCC.n15872 2.46907
R44346 VCC.n15748 VCC.n15747 2.46907
R44347 VCC.n16298 VCC.n16297 2.46907
R44348 VCC.n16424 VCC.n16423 2.46907
R44349 VCC.n16980 VCC.n16979 2.46907
R44350 VCC.n16855 VCC.n16854 2.46907
R44351 VCC.n17344 VCC.n17343 2.46907
R44352 VCC.n141 VCC.n139 2.37764
R44353 VCC.n414 VCC.n78 2.37764
R44354 VCC.n693 VCC.n691 2.37764
R44355 VCC.n966 VCC.n630 2.37764
R44356 VCC.n1523 VCC.n1187 2.37764
R44357 VCC.n1251 VCC.n1249 2.37764
R44358 VCC.n1802 VCC.n1800 2.37764
R44359 VCC.n2075 VCC.n1739 2.37764
R44360 VCC.n2632 VCC.n2296 2.37764
R44361 VCC.n2360 VCC.n2358 2.37764
R44362 VCC.n2911 VCC.n2909 2.37764
R44363 VCC.n3184 VCC.n2848 2.37764
R44364 VCC.n3741 VCC.n3405 2.37764
R44365 VCC.n3469 VCC.n3467 2.37764
R44366 VCC.n4020 VCC.n4018 2.37764
R44367 VCC.n4293 VCC.n3957 2.37764
R44368 VCC.n4850 VCC.n4514 2.37764
R44369 VCC.n4578 VCC.n4576 2.37764
R44370 VCC.n5129 VCC.n5127 2.37764
R44371 VCC.n5402 VCC.n5066 2.37764
R44372 VCC.n5959 VCC.n5623 2.37764
R44373 VCC.n5687 VCC.n5685 2.37764
R44374 VCC.n6238 VCC.n6236 2.37764
R44375 VCC.n6511 VCC.n6175 2.37764
R44376 VCC.n7068 VCC.n6732 2.37764
R44377 VCC.n6796 VCC.n6794 2.37764
R44378 VCC.n7347 VCC.n7345 2.37764
R44379 VCC.n7620 VCC.n7284 2.37764
R44380 VCC.n8177 VCC.n7841 2.37764
R44381 VCC.n7905 VCC.n7903 2.37764
R44382 VCC.n8729 VCC.n8393 2.37764
R44383 VCC.n8456 VCC.n8454 2.37764
R44384 VCC.n9286 VCC.n8950 2.37764
R44385 VCC.n9014 VCC.n9012 2.37764
R44386 VCC.n9565 VCC.n9563 2.37764
R44387 VCC.n9838 VCC.n9502 2.37764
R44388 VCC.n10394 VCC.n10058 2.37764
R44389 VCC.n10122 VCC.n10120 2.37764
R44390 VCC.n10672 VCC.n10670 2.37764
R44391 VCC.n10945 VCC.n10609 2.37764
R44392 VCC.n11501 VCC.n11165 2.37764
R44393 VCC.n11229 VCC.n11227 2.37764
R44394 VCC.n11779 VCC.n11777 2.37764
R44395 VCC.n12052 VCC.n11716 2.37764
R44396 VCC.n12608 VCC.n12272 2.37764
R44397 VCC.n12336 VCC.n12334 2.37764
R44398 VCC.n12886 VCC.n12884 2.37764
R44399 VCC.n13159 VCC.n12823 2.37764
R44400 VCC.n13715 VCC.n13379 2.37764
R44401 VCC.n13443 VCC.n13441 2.37764
R44402 VCC.n13993 VCC.n13991 2.37764
R44403 VCC.n14266 VCC.n13930 2.37764
R44404 VCC.n14822 VCC.n14486 2.37764
R44405 VCC.n14550 VCC.n14548 2.37764
R44406 VCC.n15100 VCC.n15098 2.37764
R44407 VCC.n15373 VCC.n15037 2.37764
R44408 VCC.n15929 VCC.n15593 2.37764
R44409 VCC.n15657 VCC.n15655 2.37764
R44410 VCC.n16207 VCC.n16205 2.37764
R44411 VCC.n16480 VCC.n16144 2.37764
R44412 VCC.n17036 VCC.n16700 2.37764
R44413 VCC.n16764 VCC.n16762 2.37764
R44414 VCC.n17400 VCC.n17251 2.37764
R44415 VCC.n208 VCC.n194 2.34304
R44416 VCC.n81 VCC.n79 2.34304
R44417 VCC.n123 VCC.n121 2.34304
R44418 VCC.n760 VCC.n746 2.34304
R44419 VCC.n633 VCC.n631 2.34304
R44420 VCC.n675 VCC.n673 2.34304
R44421 VCC.n1190 VCC.n1188 2.34304
R44422 VCC.n1232 VCC.n1230 2.34304
R44423 VCC.n1318 VCC.n1304 2.34304
R44424 VCC.n1869 VCC.n1855 2.34304
R44425 VCC.n1742 VCC.n1740 2.34304
R44426 VCC.n1784 VCC.n1782 2.34304
R44427 VCC.n2299 VCC.n2297 2.34304
R44428 VCC.n2341 VCC.n2339 2.34304
R44429 VCC.n2427 VCC.n2413 2.34304
R44430 VCC.n2978 VCC.n2964 2.34304
R44431 VCC.n2851 VCC.n2849 2.34304
R44432 VCC.n2893 VCC.n2891 2.34304
R44433 VCC.n3408 VCC.n3406 2.34304
R44434 VCC.n3450 VCC.n3448 2.34304
R44435 VCC.n3536 VCC.n3522 2.34304
R44436 VCC.n4087 VCC.n4073 2.34304
R44437 VCC.n3960 VCC.n3958 2.34304
R44438 VCC.n4002 VCC.n4000 2.34304
R44439 VCC.n4517 VCC.n4515 2.34304
R44440 VCC.n4559 VCC.n4557 2.34304
R44441 VCC.n4645 VCC.n4631 2.34304
R44442 VCC.n5196 VCC.n5182 2.34304
R44443 VCC.n5069 VCC.n5067 2.34304
R44444 VCC.n5111 VCC.n5109 2.34304
R44445 VCC.n5626 VCC.n5624 2.34304
R44446 VCC.n5668 VCC.n5666 2.34304
R44447 VCC.n5754 VCC.n5740 2.34304
R44448 VCC.n6305 VCC.n6291 2.34304
R44449 VCC.n6178 VCC.n6176 2.34304
R44450 VCC.n6220 VCC.n6218 2.34304
R44451 VCC.n6735 VCC.n6733 2.34304
R44452 VCC.n6777 VCC.n6775 2.34304
R44453 VCC.n6863 VCC.n6849 2.34304
R44454 VCC.n7414 VCC.n7400 2.34304
R44455 VCC.n7287 VCC.n7285 2.34304
R44456 VCC.n7329 VCC.n7327 2.34304
R44457 VCC.n7844 VCC.n7842 2.34304
R44458 VCC.n7886 VCC.n7884 2.34304
R44459 VCC.n7972 VCC.n7958 2.34304
R44460 VCC.n8396 VCC.n8394 2.34304
R44461 VCC.n8438 VCC.n8436 2.34304
R44462 VCC.n8523 VCC.n8509 2.34304
R44463 VCC.n8953 VCC.n8951 2.34304
R44464 VCC.n8995 VCC.n8993 2.34304
R44465 VCC.n9081 VCC.n9067 2.34304
R44466 VCC.n9632 VCC.n9618 2.34304
R44467 VCC.n9505 VCC.n9503 2.34304
R44468 VCC.n9547 VCC.n9545 2.34304
R44469 VCC.n10061 VCC.n10059 2.34304
R44470 VCC.n10103 VCC.n10101 2.34304
R44471 VCC.n10189 VCC.n10175 2.34304
R44472 VCC.n10739 VCC.n10725 2.34304
R44473 VCC.n10612 VCC.n10610 2.34304
R44474 VCC.n10654 VCC.n10652 2.34304
R44475 VCC.n11168 VCC.n11166 2.34304
R44476 VCC.n11210 VCC.n11208 2.34304
R44477 VCC.n11296 VCC.n11282 2.34304
R44478 VCC.n11846 VCC.n11832 2.34304
R44479 VCC.n11719 VCC.n11717 2.34304
R44480 VCC.n11761 VCC.n11759 2.34304
R44481 VCC.n12275 VCC.n12273 2.34304
R44482 VCC.n12317 VCC.n12315 2.34304
R44483 VCC.n12403 VCC.n12389 2.34304
R44484 VCC.n12953 VCC.n12939 2.34304
R44485 VCC.n12826 VCC.n12824 2.34304
R44486 VCC.n12868 VCC.n12866 2.34304
R44487 VCC.n13382 VCC.n13380 2.34304
R44488 VCC.n13424 VCC.n13422 2.34304
R44489 VCC.n13510 VCC.n13496 2.34304
R44490 VCC.n14060 VCC.n14046 2.34304
R44491 VCC.n13933 VCC.n13931 2.34304
R44492 VCC.n13975 VCC.n13973 2.34304
R44493 VCC.n14489 VCC.n14487 2.34304
R44494 VCC.n14531 VCC.n14529 2.34304
R44495 VCC.n14617 VCC.n14603 2.34304
R44496 VCC.n15167 VCC.n15153 2.34304
R44497 VCC.n15040 VCC.n15038 2.34304
R44498 VCC.n15082 VCC.n15080 2.34304
R44499 VCC.n15596 VCC.n15594 2.34304
R44500 VCC.n15638 VCC.n15636 2.34304
R44501 VCC.n15724 VCC.n15710 2.34304
R44502 VCC.n16274 VCC.n16260 2.34304
R44503 VCC.n16147 VCC.n16145 2.34304
R44504 VCC.n16189 VCC.n16187 2.34304
R44505 VCC.n16703 VCC.n16701 2.34304
R44506 VCC.n16745 VCC.n16743 2.34304
R44507 VCC.n16831 VCC.n16817 2.34304
R44508 VCC.n17254 VCC.n17252 2.34304
R44509 VCC.n17296 VCC.n17294 2.34304
R44510 VCC.n1662 VCC.n1107 2.29829
R44511 VCC.n3880 VCC.n3325 2.29829
R44512 VCC.n6098 VCC.n5543 2.29829
R44513 VCC.n8316 VCC.n7761 2.29829
R44514 VCC.n17554 VCC.n17553 2.29829
R44515 VCC.n17550 VCC.n17549 2.29829
R44516 VCC.n17546 VCC.n17545 2.29829
R44517 VCC.n17542 VCC.n17541 2.29829
R44518 VCC.n201 VCC.n183 2.28621
R44519 VCC.n326 VCC.n118 2.28621
R44520 VCC.n753 VCC.n735 2.28621
R44521 VCC.n878 VCC.n670 2.28621
R44522 VCC.n1435 VCC.n1227 2.28621
R44523 VCC.n1311 VCC.n1293 2.28621
R44524 VCC.n1862 VCC.n1844 2.28621
R44525 VCC.n1987 VCC.n1779 2.28621
R44526 VCC.n2544 VCC.n2336 2.28621
R44527 VCC.n2420 VCC.n2402 2.28621
R44528 VCC.n2971 VCC.n2953 2.28621
R44529 VCC.n3096 VCC.n2888 2.28621
R44530 VCC.n3653 VCC.n3445 2.28621
R44531 VCC.n3529 VCC.n3511 2.28621
R44532 VCC.n4080 VCC.n4062 2.28621
R44533 VCC.n4205 VCC.n3997 2.28621
R44534 VCC.n4762 VCC.n4554 2.28621
R44535 VCC.n4638 VCC.n4620 2.28621
R44536 VCC.n5189 VCC.n5171 2.28621
R44537 VCC.n5314 VCC.n5106 2.28621
R44538 VCC.n5871 VCC.n5663 2.28621
R44539 VCC.n5747 VCC.n5729 2.28621
R44540 VCC.n6298 VCC.n6280 2.28621
R44541 VCC.n6423 VCC.n6215 2.28621
R44542 VCC.n6980 VCC.n6772 2.28621
R44543 VCC.n6856 VCC.n6838 2.28621
R44544 VCC.n7407 VCC.n7389 2.28621
R44545 VCC.n7532 VCC.n7324 2.28621
R44546 VCC.n8089 VCC.n7881 2.28621
R44547 VCC.n7965 VCC.n7947 2.28621
R44548 VCC.n8641 VCC.n8433 2.28621
R44549 VCC.n8516 VCC.n8498 2.28621
R44550 VCC.n9198 VCC.n8990 2.28621
R44551 VCC.n9074 VCC.n9056 2.28621
R44552 VCC.n9625 VCC.n9607 2.28621
R44553 VCC.n9750 VCC.n9542 2.28621
R44554 VCC.n10306 VCC.n10098 2.28621
R44555 VCC.n10182 VCC.n10164 2.28621
R44556 VCC.n10732 VCC.n10714 2.28621
R44557 VCC.n10857 VCC.n10649 2.28621
R44558 VCC.n11413 VCC.n11205 2.28621
R44559 VCC.n11289 VCC.n11271 2.28621
R44560 VCC.n11839 VCC.n11821 2.28621
R44561 VCC.n11964 VCC.n11756 2.28621
R44562 VCC.n12520 VCC.n12312 2.28621
R44563 VCC.n12396 VCC.n12378 2.28621
R44564 VCC.n12946 VCC.n12928 2.28621
R44565 VCC.n13071 VCC.n12863 2.28621
R44566 VCC.n13627 VCC.n13419 2.28621
R44567 VCC.n13503 VCC.n13485 2.28621
R44568 VCC.n14053 VCC.n14035 2.28621
R44569 VCC.n14178 VCC.n13970 2.28621
R44570 VCC.n14734 VCC.n14526 2.28621
R44571 VCC.n14610 VCC.n14592 2.28621
R44572 VCC.n15160 VCC.n15142 2.28621
R44573 VCC.n15285 VCC.n15077 2.28621
R44574 VCC.n15841 VCC.n15633 2.28621
R44575 VCC.n15717 VCC.n15699 2.28621
R44576 VCC.n16267 VCC.n16249 2.28621
R44577 VCC.n16392 VCC.n16184 2.28621
R44578 VCC.n16948 VCC.n16740 2.28621
R44579 VCC.n16824 VCC.n16806 2.28621
R44580 VCC.n17312 VCC.n17291 2.28621
R44581 VCC.n130 VCC.n129 2.2505
R44582 VCC.n304 VCC.n133 2.2505
R44583 VCC.n277 VCC.n149 2.2505
R44584 VCC.n193 VCC.n190 2.2505
R44585 VCC.n186 VCC.n185 2.2505
R44586 VCC.n235 VCC.n234 2.2505
R44587 VCC.n69 VCC.n68 2.2505
R44588 VCC.n439 VCC.n72 2.2505
R44589 VCC.n404 VCC.n89 2.2505
R44590 VCC.n332 VCC.n319 2.2505
R44591 VCC.n116 VCC.n115 2.2505
R44592 VCC.n351 VCC.n349 2.2505
R44593 VCC.n539 VCC.n12 2.2505
R44594 VCC.n465 VCC.n59 2.2505
R44595 VCC.n488 VCC.n487 2.2505
R44596 VCC.n28 VCC.n26 2.2505
R44597 VCC.n533 VCC.n15 2.2505
R44598 VCC.n457 VCC.n64 2.2505
R44599 VCC.n682 VCC.n681 2.2505
R44600 VCC.n856 VCC.n685 2.2505
R44601 VCC.n829 VCC.n701 2.2505
R44602 VCC.n745 VCC.n742 2.2505
R44603 VCC.n738 VCC.n737 2.2505
R44604 VCC.n787 VCC.n786 2.2505
R44605 VCC.n621 VCC.n620 2.2505
R44606 VCC.n991 VCC.n624 2.2505
R44607 VCC.n956 VCC.n641 2.2505
R44608 VCC.n884 VCC.n871 2.2505
R44609 VCC.n668 VCC.n667 2.2505
R44610 VCC.n903 VCC.n901 2.2505
R44611 VCC.n1093 VCC.n1092 2.2505
R44612 VCC.n1085 VCC.n567 2.2505
R44613 VCC.n580 VCC.n578 2.2505
R44614 VCC.n1009 VCC.n616 2.2505
R44615 VCC.n1017 VCC.n611 2.2505
R44616 VCC.n1040 VCC.n1039 2.2505
R44617 VCC.n1639 VCC.n1638 2.2505
R44618 VCC.n1590 VCC.n1589 2.2505
R44619 VCC.n1120 VCC.n1118 2.2505
R44620 VCC.n1625 VCC.n1132 2.2505
R44621 VCC.n1575 VCC.n1574 2.2505
R44622 VCC.n1568 VCC.n1173 2.2505
R44623 VCC.n1178 VCC.n1177 2.2505
R44624 VCC.n1549 VCC.n1181 2.2505
R44625 VCC.n1513 VCC.n1198 2.2505
R44626 VCC.n1460 VCC.n1458 2.2505
R44627 VCC.n1225 VCC.n1224 2.2505
R44628 VCC.n1441 VCC.n1440 2.2505
R44629 VCC.n1240 VCC.n1239 2.2505
R44630 VCC.n1414 VCC.n1243 2.2505
R44631 VCC.n1387 VCC.n1259 2.2505
R44632 VCC.n1345 VCC.n1344 2.2505
R44633 VCC.n1296 VCC.n1295 2.2505
R44634 VCC.n1303 VCC.n1300 2.2505
R44635 VCC.n1791 VCC.n1790 2.2505
R44636 VCC.n1965 VCC.n1794 2.2505
R44637 VCC.n1938 VCC.n1810 2.2505
R44638 VCC.n1854 VCC.n1851 2.2505
R44639 VCC.n1847 VCC.n1846 2.2505
R44640 VCC.n1896 VCC.n1895 2.2505
R44641 VCC.n1730 VCC.n1729 2.2505
R44642 VCC.n2100 VCC.n1733 2.2505
R44643 VCC.n2065 VCC.n1750 2.2505
R44644 VCC.n1993 VCC.n1980 2.2505
R44645 VCC.n1777 VCC.n1776 2.2505
R44646 VCC.n2012 VCC.n2010 2.2505
R44647 VCC.n2202 VCC.n2201 2.2505
R44648 VCC.n2194 VCC.n1676 2.2505
R44649 VCC.n1689 VCC.n1687 2.2505
R44650 VCC.n2118 VCC.n1725 2.2505
R44651 VCC.n2126 VCC.n1720 2.2505
R44652 VCC.n2149 VCC.n2148 2.2505
R44653 VCC.n2748 VCC.n2747 2.2505
R44654 VCC.n2699 VCC.n2698 2.2505
R44655 VCC.n2229 VCC.n2227 2.2505
R44656 VCC.n2734 VCC.n2241 2.2505
R44657 VCC.n2684 VCC.n2683 2.2505
R44658 VCC.n2677 VCC.n2282 2.2505
R44659 VCC.n2287 VCC.n2286 2.2505
R44660 VCC.n2658 VCC.n2290 2.2505
R44661 VCC.n2622 VCC.n2307 2.2505
R44662 VCC.n2569 VCC.n2567 2.2505
R44663 VCC.n2334 VCC.n2333 2.2505
R44664 VCC.n2550 VCC.n2549 2.2505
R44665 VCC.n2349 VCC.n2348 2.2505
R44666 VCC.n2523 VCC.n2352 2.2505
R44667 VCC.n2496 VCC.n2368 2.2505
R44668 VCC.n2454 VCC.n2453 2.2505
R44669 VCC.n2405 VCC.n2404 2.2505
R44670 VCC.n2412 VCC.n2409 2.2505
R44671 VCC.n2900 VCC.n2899 2.2505
R44672 VCC.n3074 VCC.n2903 2.2505
R44673 VCC.n3047 VCC.n2919 2.2505
R44674 VCC.n2963 VCC.n2960 2.2505
R44675 VCC.n2956 VCC.n2955 2.2505
R44676 VCC.n3005 VCC.n3004 2.2505
R44677 VCC.n2839 VCC.n2838 2.2505
R44678 VCC.n3209 VCC.n2842 2.2505
R44679 VCC.n3174 VCC.n2859 2.2505
R44680 VCC.n3102 VCC.n3089 2.2505
R44681 VCC.n2886 VCC.n2885 2.2505
R44682 VCC.n3121 VCC.n3119 2.2505
R44683 VCC.n3311 VCC.n3310 2.2505
R44684 VCC.n3303 VCC.n2785 2.2505
R44685 VCC.n2798 VCC.n2796 2.2505
R44686 VCC.n3227 VCC.n2834 2.2505
R44687 VCC.n3235 VCC.n2829 2.2505
R44688 VCC.n3258 VCC.n3257 2.2505
R44689 VCC.n3857 VCC.n3856 2.2505
R44690 VCC.n3808 VCC.n3807 2.2505
R44691 VCC.n3338 VCC.n3336 2.2505
R44692 VCC.n3843 VCC.n3350 2.2505
R44693 VCC.n3793 VCC.n3792 2.2505
R44694 VCC.n3786 VCC.n3391 2.2505
R44695 VCC.n3396 VCC.n3395 2.2505
R44696 VCC.n3767 VCC.n3399 2.2505
R44697 VCC.n3731 VCC.n3416 2.2505
R44698 VCC.n3678 VCC.n3676 2.2505
R44699 VCC.n3443 VCC.n3442 2.2505
R44700 VCC.n3659 VCC.n3658 2.2505
R44701 VCC.n3458 VCC.n3457 2.2505
R44702 VCC.n3632 VCC.n3461 2.2505
R44703 VCC.n3605 VCC.n3477 2.2505
R44704 VCC.n3563 VCC.n3562 2.2505
R44705 VCC.n3514 VCC.n3513 2.2505
R44706 VCC.n3521 VCC.n3518 2.2505
R44707 VCC.n4009 VCC.n4008 2.2505
R44708 VCC.n4183 VCC.n4012 2.2505
R44709 VCC.n4156 VCC.n4028 2.2505
R44710 VCC.n4072 VCC.n4069 2.2505
R44711 VCC.n4065 VCC.n4064 2.2505
R44712 VCC.n4114 VCC.n4113 2.2505
R44713 VCC.n3948 VCC.n3947 2.2505
R44714 VCC.n4318 VCC.n3951 2.2505
R44715 VCC.n4283 VCC.n3968 2.2505
R44716 VCC.n4211 VCC.n4198 2.2505
R44717 VCC.n3995 VCC.n3994 2.2505
R44718 VCC.n4230 VCC.n4228 2.2505
R44719 VCC.n4420 VCC.n4419 2.2505
R44720 VCC.n4412 VCC.n3894 2.2505
R44721 VCC.n3907 VCC.n3905 2.2505
R44722 VCC.n4336 VCC.n3943 2.2505
R44723 VCC.n4344 VCC.n3938 2.2505
R44724 VCC.n4367 VCC.n4366 2.2505
R44725 VCC.n4966 VCC.n4965 2.2505
R44726 VCC.n4917 VCC.n4916 2.2505
R44727 VCC.n4447 VCC.n4445 2.2505
R44728 VCC.n4952 VCC.n4459 2.2505
R44729 VCC.n4902 VCC.n4901 2.2505
R44730 VCC.n4895 VCC.n4500 2.2505
R44731 VCC.n4505 VCC.n4504 2.2505
R44732 VCC.n4876 VCC.n4508 2.2505
R44733 VCC.n4840 VCC.n4525 2.2505
R44734 VCC.n4787 VCC.n4785 2.2505
R44735 VCC.n4552 VCC.n4551 2.2505
R44736 VCC.n4768 VCC.n4767 2.2505
R44737 VCC.n4567 VCC.n4566 2.2505
R44738 VCC.n4741 VCC.n4570 2.2505
R44739 VCC.n4714 VCC.n4586 2.2505
R44740 VCC.n4672 VCC.n4671 2.2505
R44741 VCC.n4623 VCC.n4622 2.2505
R44742 VCC.n4630 VCC.n4627 2.2505
R44743 VCC.n5118 VCC.n5117 2.2505
R44744 VCC.n5292 VCC.n5121 2.2505
R44745 VCC.n5265 VCC.n5137 2.2505
R44746 VCC.n5181 VCC.n5178 2.2505
R44747 VCC.n5174 VCC.n5173 2.2505
R44748 VCC.n5223 VCC.n5222 2.2505
R44749 VCC.n5057 VCC.n5056 2.2505
R44750 VCC.n5427 VCC.n5060 2.2505
R44751 VCC.n5392 VCC.n5077 2.2505
R44752 VCC.n5320 VCC.n5307 2.2505
R44753 VCC.n5104 VCC.n5103 2.2505
R44754 VCC.n5339 VCC.n5337 2.2505
R44755 VCC.n5529 VCC.n5528 2.2505
R44756 VCC.n5521 VCC.n5003 2.2505
R44757 VCC.n5016 VCC.n5014 2.2505
R44758 VCC.n5445 VCC.n5052 2.2505
R44759 VCC.n5453 VCC.n5047 2.2505
R44760 VCC.n5476 VCC.n5475 2.2505
R44761 VCC.n6075 VCC.n6074 2.2505
R44762 VCC.n6026 VCC.n6025 2.2505
R44763 VCC.n5556 VCC.n5554 2.2505
R44764 VCC.n6061 VCC.n5568 2.2505
R44765 VCC.n6011 VCC.n6010 2.2505
R44766 VCC.n6004 VCC.n5609 2.2505
R44767 VCC.n5614 VCC.n5613 2.2505
R44768 VCC.n5985 VCC.n5617 2.2505
R44769 VCC.n5949 VCC.n5634 2.2505
R44770 VCC.n5896 VCC.n5894 2.2505
R44771 VCC.n5661 VCC.n5660 2.2505
R44772 VCC.n5877 VCC.n5876 2.2505
R44773 VCC.n5676 VCC.n5675 2.2505
R44774 VCC.n5850 VCC.n5679 2.2505
R44775 VCC.n5823 VCC.n5695 2.2505
R44776 VCC.n5781 VCC.n5780 2.2505
R44777 VCC.n5732 VCC.n5731 2.2505
R44778 VCC.n5739 VCC.n5736 2.2505
R44779 VCC.n6227 VCC.n6226 2.2505
R44780 VCC.n6401 VCC.n6230 2.2505
R44781 VCC.n6374 VCC.n6246 2.2505
R44782 VCC.n6290 VCC.n6287 2.2505
R44783 VCC.n6283 VCC.n6282 2.2505
R44784 VCC.n6332 VCC.n6331 2.2505
R44785 VCC.n6166 VCC.n6165 2.2505
R44786 VCC.n6536 VCC.n6169 2.2505
R44787 VCC.n6501 VCC.n6186 2.2505
R44788 VCC.n6429 VCC.n6416 2.2505
R44789 VCC.n6213 VCC.n6212 2.2505
R44790 VCC.n6448 VCC.n6446 2.2505
R44791 VCC.n6638 VCC.n6637 2.2505
R44792 VCC.n6630 VCC.n6112 2.2505
R44793 VCC.n6125 VCC.n6123 2.2505
R44794 VCC.n6554 VCC.n6161 2.2505
R44795 VCC.n6562 VCC.n6156 2.2505
R44796 VCC.n6585 VCC.n6584 2.2505
R44797 VCC.n7184 VCC.n7183 2.2505
R44798 VCC.n7135 VCC.n7134 2.2505
R44799 VCC.n6665 VCC.n6663 2.2505
R44800 VCC.n7170 VCC.n6677 2.2505
R44801 VCC.n7120 VCC.n7119 2.2505
R44802 VCC.n7113 VCC.n6718 2.2505
R44803 VCC.n6723 VCC.n6722 2.2505
R44804 VCC.n7094 VCC.n6726 2.2505
R44805 VCC.n7058 VCC.n6743 2.2505
R44806 VCC.n7005 VCC.n7003 2.2505
R44807 VCC.n6770 VCC.n6769 2.2505
R44808 VCC.n6986 VCC.n6985 2.2505
R44809 VCC.n6785 VCC.n6784 2.2505
R44810 VCC.n6959 VCC.n6788 2.2505
R44811 VCC.n6932 VCC.n6804 2.2505
R44812 VCC.n6890 VCC.n6889 2.2505
R44813 VCC.n6841 VCC.n6840 2.2505
R44814 VCC.n6848 VCC.n6845 2.2505
R44815 VCC.n7336 VCC.n7335 2.2505
R44816 VCC.n7510 VCC.n7339 2.2505
R44817 VCC.n7483 VCC.n7355 2.2505
R44818 VCC.n7399 VCC.n7396 2.2505
R44819 VCC.n7392 VCC.n7391 2.2505
R44820 VCC.n7441 VCC.n7440 2.2505
R44821 VCC.n7275 VCC.n7274 2.2505
R44822 VCC.n7645 VCC.n7278 2.2505
R44823 VCC.n7610 VCC.n7295 2.2505
R44824 VCC.n7538 VCC.n7525 2.2505
R44825 VCC.n7322 VCC.n7321 2.2505
R44826 VCC.n7557 VCC.n7555 2.2505
R44827 VCC.n7747 VCC.n7746 2.2505
R44828 VCC.n7739 VCC.n7221 2.2505
R44829 VCC.n7234 VCC.n7232 2.2505
R44830 VCC.n7663 VCC.n7270 2.2505
R44831 VCC.n7671 VCC.n7265 2.2505
R44832 VCC.n7694 VCC.n7693 2.2505
R44833 VCC.n8293 VCC.n8292 2.2505
R44834 VCC.n8244 VCC.n8243 2.2505
R44835 VCC.n7774 VCC.n7772 2.2505
R44836 VCC.n8279 VCC.n7786 2.2505
R44837 VCC.n8229 VCC.n8228 2.2505
R44838 VCC.n8222 VCC.n7827 2.2505
R44839 VCC.n7832 VCC.n7831 2.2505
R44840 VCC.n8203 VCC.n7835 2.2505
R44841 VCC.n8167 VCC.n7852 2.2505
R44842 VCC.n8114 VCC.n8112 2.2505
R44843 VCC.n7879 VCC.n7878 2.2505
R44844 VCC.n8095 VCC.n8094 2.2505
R44845 VCC.n7894 VCC.n7893 2.2505
R44846 VCC.n8068 VCC.n7897 2.2505
R44847 VCC.n8041 VCC.n7913 2.2505
R44848 VCC.n7999 VCC.n7998 2.2505
R44849 VCC.n7950 VCC.n7949 2.2505
R44850 VCC.n7957 VCC.n7954 2.2505
R44851 VCC.n8384 VCC.n8383 2.2505
R44852 VCC.n8754 VCC.n8387 2.2505
R44853 VCC.n8719 VCC.n8404 2.2505
R44854 VCC.n8647 VCC.n8634 2.2505
R44855 VCC.n8431 VCC.n8430 2.2505
R44856 VCC.n8666 VCC.n8664 2.2505
R44857 VCC.n8856 VCC.n8855 2.2505
R44858 VCC.n8848 VCC.n8330 2.2505
R44859 VCC.n8343 VCC.n8341 2.2505
R44860 VCC.n8772 VCC.n8379 2.2505
R44861 VCC.n8780 VCC.n8374 2.2505
R44862 VCC.n8803 VCC.n8802 2.2505
R44863 VCC.n8445 VCC.n8444 2.2505
R44864 VCC.n8619 VCC.n8448 2.2505
R44865 VCC.n8592 VCC.n8464 2.2505
R44866 VCC.n8550 VCC.n8549 2.2505
R44867 VCC.n8501 VCC.n8500 2.2505
R44868 VCC.n8508 VCC.n8505 2.2505
R44869 VCC.n9402 VCC.n9401 2.2505
R44870 VCC.n9353 VCC.n9352 2.2505
R44871 VCC.n8883 VCC.n8881 2.2505
R44872 VCC.n9388 VCC.n8895 2.2505
R44873 VCC.n9338 VCC.n9337 2.2505
R44874 VCC.n9331 VCC.n8936 2.2505
R44875 VCC.n8941 VCC.n8940 2.2505
R44876 VCC.n9312 VCC.n8944 2.2505
R44877 VCC.n9276 VCC.n8961 2.2505
R44878 VCC.n9223 VCC.n9221 2.2505
R44879 VCC.n8988 VCC.n8987 2.2505
R44880 VCC.n9204 VCC.n9203 2.2505
R44881 VCC.n9003 VCC.n9002 2.2505
R44882 VCC.n9177 VCC.n9006 2.2505
R44883 VCC.n9150 VCC.n9022 2.2505
R44884 VCC.n9108 VCC.n9107 2.2505
R44885 VCC.n9059 VCC.n9058 2.2505
R44886 VCC.n9066 VCC.n9063 2.2505
R44887 VCC.n9554 VCC.n9553 2.2505
R44888 VCC.n9728 VCC.n9557 2.2505
R44889 VCC.n9701 VCC.n9573 2.2505
R44890 VCC.n9617 VCC.n9614 2.2505
R44891 VCC.n9610 VCC.n9609 2.2505
R44892 VCC.n9659 VCC.n9658 2.2505
R44893 VCC.n9493 VCC.n9492 2.2505
R44894 VCC.n9863 VCC.n9496 2.2505
R44895 VCC.n9828 VCC.n9513 2.2505
R44896 VCC.n9756 VCC.n9743 2.2505
R44897 VCC.n9540 VCC.n9539 2.2505
R44898 VCC.n9775 VCC.n9773 2.2505
R44899 VCC.n9965 VCC.n9964 2.2505
R44900 VCC.n9957 VCC.n9439 2.2505
R44901 VCC.n9452 VCC.n9450 2.2505
R44902 VCC.n9881 VCC.n9488 2.2505
R44903 VCC.n9889 VCC.n9483 2.2505
R44904 VCC.n9912 VCC.n9911 2.2505
R44905 VCC.n10510 VCC.n10509 2.2505
R44906 VCC.n10461 VCC.n10460 2.2505
R44907 VCC.n9991 VCC.n9989 2.2505
R44908 VCC.n10496 VCC.n10003 2.2505
R44909 VCC.n10446 VCC.n10445 2.2505
R44910 VCC.n10439 VCC.n10044 2.2505
R44911 VCC.n10049 VCC.n10048 2.2505
R44912 VCC.n10420 VCC.n10052 2.2505
R44913 VCC.n10384 VCC.n10069 2.2505
R44914 VCC.n10331 VCC.n10329 2.2505
R44915 VCC.n10096 VCC.n10095 2.2505
R44916 VCC.n10312 VCC.n10311 2.2505
R44917 VCC.n10111 VCC.n10110 2.2505
R44918 VCC.n10285 VCC.n10114 2.2505
R44919 VCC.n10258 VCC.n10130 2.2505
R44920 VCC.n10216 VCC.n10215 2.2505
R44921 VCC.n10167 VCC.n10166 2.2505
R44922 VCC.n10174 VCC.n10171 2.2505
R44923 VCC.n10661 VCC.n10660 2.2505
R44924 VCC.n10835 VCC.n10664 2.2505
R44925 VCC.n10808 VCC.n10680 2.2505
R44926 VCC.n10724 VCC.n10721 2.2505
R44927 VCC.n10717 VCC.n10716 2.2505
R44928 VCC.n10766 VCC.n10765 2.2505
R44929 VCC.n10600 VCC.n10599 2.2505
R44930 VCC.n10970 VCC.n10603 2.2505
R44931 VCC.n10935 VCC.n10620 2.2505
R44932 VCC.n10863 VCC.n10850 2.2505
R44933 VCC.n10647 VCC.n10646 2.2505
R44934 VCC.n10882 VCC.n10880 2.2505
R44935 VCC.n11072 VCC.n11071 2.2505
R44936 VCC.n11064 VCC.n10546 2.2505
R44937 VCC.n10559 VCC.n10557 2.2505
R44938 VCC.n10988 VCC.n10595 2.2505
R44939 VCC.n10996 VCC.n10590 2.2505
R44940 VCC.n11019 VCC.n11018 2.2505
R44941 VCC.n11617 VCC.n11616 2.2505
R44942 VCC.n11568 VCC.n11567 2.2505
R44943 VCC.n11098 VCC.n11096 2.2505
R44944 VCC.n11603 VCC.n11110 2.2505
R44945 VCC.n11553 VCC.n11552 2.2505
R44946 VCC.n11546 VCC.n11151 2.2505
R44947 VCC.n11156 VCC.n11155 2.2505
R44948 VCC.n11527 VCC.n11159 2.2505
R44949 VCC.n11491 VCC.n11176 2.2505
R44950 VCC.n11438 VCC.n11436 2.2505
R44951 VCC.n11203 VCC.n11202 2.2505
R44952 VCC.n11419 VCC.n11418 2.2505
R44953 VCC.n11218 VCC.n11217 2.2505
R44954 VCC.n11392 VCC.n11221 2.2505
R44955 VCC.n11365 VCC.n11237 2.2505
R44956 VCC.n11323 VCC.n11322 2.2505
R44957 VCC.n11274 VCC.n11273 2.2505
R44958 VCC.n11281 VCC.n11278 2.2505
R44959 VCC.n11768 VCC.n11767 2.2505
R44960 VCC.n11942 VCC.n11771 2.2505
R44961 VCC.n11915 VCC.n11787 2.2505
R44962 VCC.n11831 VCC.n11828 2.2505
R44963 VCC.n11824 VCC.n11823 2.2505
R44964 VCC.n11873 VCC.n11872 2.2505
R44965 VCC.n11707 VCC.n11706 2.2505
R44966 VCC.n12077 VCC.n11710 2.2505
R44967 VCC.n12042 VCC.n11727 2.2505
R44968 VCC.n11970 VCC.n11957 2.2505
R44969 VCC.n11754 VCC.n11753 2.2505
R44970 VCC.n11989 VCC.n11987 2.2505
R44971 VCC.n12179 VCC.n12178 2.2505
R44972 VCC.n12171 VCC.n11653 2.2505
R44973 VCC.n11666 VCC.n11664 2.2505
R44974 VCC.n12095 VCC.n11702 2.2505
R44975 VCC.n12103 VCC.n11697 2.2505
R44976 VCC.n12126 VCC.n12125 2.2505
R44977 VCC.n12724 VCC.n12723 2.2505
R44978 VCC.n12675 VCC.n12674 2.2505
R44979 VCC.n12205 VCC.n12203 2.2505
R44980 VCC.n12710 VCC.n12217 2.2505
R44981 VCC.n12660 VCC.n12659 2.2505
R44982 VCC.n12653 VCC.n12258 2.2505
R44983 VCC.n12263 VCC.n12262 2.2505
R44984 VCC.n12634 VCC.n12266 2.2505
R44985 VCC.n12598 VCC.n12283 2.2505
R44986 VCC.n12545 VCC.n12543 2.2505
R44987 VCC.n12310 VCC.n12309 2.2505
R44988 VCC.n12526 VCC.n12525 2.2505
R44989 VCC.n12325 VCC.n12324 2.2505
R44990 VCC.n12499 VCC.n12328 2.2505
R44991 VCC.n12472 VCC.n12344 2.2505
R44992 VCC.n12430 VCC.n12429 2.2505
R44993 VCC.n12381 VCC.n12380 2.2505
R44994 VCC.n12388 VCC.n12385 2.2505
R44995 VCC.n12875 VCC.n12874 2.2505
R44996 VCC.n13049 VCC.n12878 2.2505
R44997 VCC.n13022 VCC.n12894 2.2505
R44998 VCC.n12938 VCC.n12935 2.2505
R44999 VCC.n12931 VCC.n12930 2.2505
R45000 VCC.n12980 VCC.n12979 2.2505
R45001 VCC.n12814 VCC.n12813 2.2505
R45002 VCC.n13184 VCC.n12817 2.2505
R45003 VCC.n13149 VCC.n12834 2.2505
R45004 VCC.n13077 VCC.n13064 2.2505
R45005 VCC.n12861 VCC.n12860 2.2505
R45006 VCC.n13096 VCC.n13094 2.2505
R45007 VCC.n13286 VCC.n13285 2.2505
R45008 VCC.n13278 VCC.n12760 2.2505
R45009 VCC.n12773 VCC.n12771 2.2505
R45010 VCC.n13202 VCC.n12809 2.2505
R45011 VCC.n13210 VCC.n12804 2.2505
R45012 VCC.n13233 VCC.n13232 2.2505
R45013 VCC.n13831 VCC.n13830 2.2505
R45014 VCC.n13782 VCC.n13781 2.2505
R45015 VCC.n13312 VCC.n13310 2.2505
R45016 VCC.n13817 VCC.n13324 2.2505
R45017 VCC.n13767 VCC.n13766 2.2505
R45018 VCC.n13760 VCC.n13365 2.2505
R45019 VCC.n13370 VCC.n13369 2.2505
R45020 VCC.n13741 VCC.n13373 2.2505
R45021 VCC.n13705 VCC.n13390 2.2505
R45022 VCC.n13652 VCC.n13650 2.2505
R45023 VCC.n13417 VCC.n13416 2.2505
R45024 VCC.n13633 VCC.n13632 2.2505
R45025 VCC.n13432 VCC.n13431 2.2505
R45026 VCC.n13606 VCC.n13435 2.2505
R45027 VCC.n13579 VCC.n13451 2.2505
R45028 VCC.n13537 VCC.n13536 2.2505
R45029 VCC.n13488 VCC.n13487 2.2505
R45030 VCC.n13495 VCC.n13492 2.2505
R45031 VCC.n13982 VCC.n13981 2.2505
R45032 VCC.n14156 VCC.n13985 2.2505
R45033 VCC.n14129 VCC.n14001 2.2505
R45034 VCC.n14045 VCC.n14042 2.2505
R45035 VCC.n14038 VCC.n14037 2.2505
R45036 VCC.n14087 VCC.n14086 2.2505
R45037 VCC.n13921 VCC.n13920 2.2505
R45038 VCC.n14291 VCC.n13924 2.2505
R45039 VCC.n14256 VCC.n13941 2.2505
R45040 VCC.n14184 VCC.n14171 2.2505
R45041 VCC.n13968 VCC.n13967 2.2505
R45042 VCC.n14203 VCC.n14201 2.2505
R45043 VCC.n14393 VCC.n14392 2.2505
R45044 VCC.n14385 VCC.n13867 2.2505
R45045 VCC.n13880 VCC.n13878 2.2505
R45046 VCC.n14309 VCC.n13916 2.2505
R45047 VCC.n14317 VCC.n13911 2.2505
R45048 VCC.n14340 VCC.n14339 2.2505
R45049 VCC.n14938 VCC.n14937 2.2505
R45050 VCC.n14889 VCC.n14888 2.2505
R45051 VCC.n14419 VCC.n14417 2.2505
R45052 VCC.n14924 VCC.n14431 2.2505
R45053 VCC.n14874 VCC.n14873 2.2505
R45054 VCC.n14867 VCC.n14472 2.2505
R45055 VCC.n14477 VCC.n14476 2.2505
R45056 VCC.n14848 VCC.n14480 2.2505
R45057 VCC.n14812 VCC.n14497 2.2505
R45058 VCC.n14759 VCC.n14757 2.2505
R45059 VCC.n14524 VCC.n14523 2.2505
R45060 VCC.n14740 VCC.n14739 2.2505
R45061 VCC.n14539 VCC.n14538 2.2505
R45062 VCC.n14713 VCC.n14542 2.2505
R45063 VCC.n14686 VCC.n14558 2.2505
R45064 VCC.n14644 VCC.n14643 2.2505
R45065 VCC.n14595 VCC.n14594 2.2505
R45066 VCC.n14602 VCC.n14599 2.2505
R45067 VCC.n15089 VCC.n15088 2.2505
R45068 VCC.n15263 VCC.n15092 2.2505
R45069 VCC.n15236 VCC.n15108 2.2505
R45070 VCC.n15152 VCC.n15149 2.2505
R45071 VCC.n15145 VCC.n15144 2.2505
R45072 VCC.n15194 VCC.n15193 2.2505
R45073 VCC.n15028 VCC.n15027 2.2505
R45074 VCC.n15398 VCC.n15031 2.2505
R45075 VCC.n15363 VCC.n15048 2.2505
R45076 VCC.n15291 VCC.n15278 2.2505
R45077 VCC.n15075 VCC.n15074 2.2505
R45078 VCC.n15310 VCC.n15308 2.2505
R45079 VCC.n15500 VCC.n15499 2.2505
R45080 VCC.n15492 VCC.n14974 2.2505
R45081 VCC.n14987 VCC.n14985 2.2505
R45082 VCC.n15416 VCC.n15023 2.2505
R45083 VCC.n15424 VCC.n15018 2.2505
R45084 VCC.n15447 VCC.n15446 2.2505
R45085 VCC.n16045 VCC.n16044 2.2505
R45086 VCC.n15996 VCC.n15995 2.2505
R45087 VCC.n15526 VCC.n15524 2.2505
R45088 VCC.n16031 VCC.n15538 2.2505
R45089 VCC.n15981 VCC.n15980 2.2505
R45090 VCC.n15974 VCC.n15579 2.2505
R45091 VCC.n15584 VCC.n15583 2.2505
R45092 VCC.n15955 VCC.n15587 2.2505
R45093 VCC.n15919 VCC.n15604 2.2505
R45094 VCC.n15866 VCC.n15864 2.2505
R45095 VCC.n15631 VCC.n15630 2.2505
R45096 VCC.n15847 VCC.n15846 2.2505
R45097 VCC.n15646 VCC.n15645 2.2505
R45098 VCC.n15820 VCC.n15649 2.2505
R45099 VCC.n15793 VCC.n15665 2.2505
R45100 VCC.n15751 VCC.n15750 2.2505
R45101 VCC.n15702 VCC.n15701 2.2505
R45102 VCC.n15709 VCC.n15706 2.2505
R45103 VCC.n16196 VCC.n16195 2.2505
R45104 VCC.n16370 VCC.n16199 2.2505
R45105 VCC.n16343 VCC.n16215 2.2505
R45106 VCC.n16259 VCC.n16256 2.2505
R45107 VCC.n16252 VCC.n16251 2.2505
R45108 VCC.n16301 VCC.n16300 2.2505
R45109 VCC.n16135 VCC.n16134 2.2505
R45110 VCC.n16505 VCC.n16138 2.2505
R45111 VCC.n16470 VCC.n16155 2.2505
R45112 VCC.n16398 VCC.n16385 2.2505
R45113 VCC.n16182 VCC.n16181 2.2505
R45114 VCC.n16417 VCC.n16415 2.2505
R45115 VCC.n16607 VCC.n16606 2.2505
R45116 VCC.n16599 VCC.n16081 2.2505
R45117 VCC.n16094 VCC.n16092 2.2505
R45118 VCC.n16523 VCC.n16130 2.2505
R45119 VCC.n16531 VCC.n16125 2.2505
R45120 VCC.n16554 VCC.n16553 2.2505
R45121 VCC.n17152 VCC.n17151 2.2505
R45122 VCC.n17103 VCC.n17102 2.2505
R45123 VCC.n16633 VCC.n16631 2.2505
R45124 VCC.n17138 VCC.n16645 2.2505
R45125 VCC.n17088 VCC.n17087 2.2505
R45126 VCC.n17081 VCC.n16686 2.2505
R45127 VCC.n16691 VCC.n16690 2.2505
R45128 VCC.n17062 VCC.n16694 2.2505
R45129 VCC.n17026 VCC.n16711 2.2505
R45130 VCC.n16973 VCC.n16971 2.2505
R45131 VCC.n16738 VCC.n16737 2.2505
R45132 VCC.n16954 VCC.n16953 2.2505
R45133 VCC.n16753 VCC.n16752 2.2505
R45134 VCC.n16927 VCC.n16756 2.2505
R45135 VCC.n16900 VCC.n16772 2.2505
R45136 VCC.n16858 VCC.n16857 2.2505
R45137 VCC.n16809 VCC.n16808 2.2505
R45138 VCC.n16816 VCC.n16813 2.2505
R45139 VCC.n17242 VCC.n17241 2.2505
R45140 VCC.n17425 VCC.n17245 2.2505
R45141 VCC.n17390 VCC.n17262 2.2505
R45142 VCC.n17318 VCC.n17305 2.2505
R45143 VCC.n17289 VCC.n17288 2.2505
R45144 VCC.n17337 VCC.n17335 2.2505
R45145 VCC.n17527 VCC.n17526 2.2505
R45146 VCC.n17519 VCC.n17188 2.2505
R45147 VCC.n17201 VCC.n17199 2.2505
R45148 VCC.n17443 VCC.n17237 2.2505
R45149 VCC.n17451 VCC.n17232 2.2505
R45150 VCC.n17474 VCC.n17473 2.2505
R45151 VCC.n17541 VCC 2.24163
R45152 VCC.n2216 VCC.n1662 2.21741
R45153 VCC.n4434 VCC.n3880 2.21741
R45154 VCC.n6652 VCC.n6098 2.21741
R45155 VCC.n8870 VCC.n8316 2.21741
R45156 VCC.n17553 VCC.n17552 2.21741
R45157 VCC.n17549 VCC.n17548 2.21741
R45158 VCC.n17545 VCC.n17544 2.21741
R45159 VCC.n264 VCC.n263 2.10336
R45160 VCC.n386 VCC.n385 2.10336
R45161 VCC.n816 VCC.n815 2.10336
R45162 VCC.n938 VCC.n937 2.10336
R45163 VCC.n1495 VCC.n1494 2.10336
R45164 VCC.n1374 VCC.n1373 2.10336
R45165 VCC.n1925 VCC.n1924 2.10336
R45166 VCC.n2047 VCC.n2046 2.10336
R45167 VCC.n2604 VCC.n2603 2.10336
R45168 VCC.n2483 VCC.n2482 2.10336
R45169 VCC.n3034 VCC.n3033 2.10336
R45170 VCC.n3156 VCC.n3155 2.10336
R45171 VCC.n3713 VCC.n3712 2.10336
R45172 VCC.n3592 VCC.n3591 2.10336
R45173 VCC.n4143 VCC.n4142 2.10336
R45174 VCC.n4265 VCC.n4264 2.10336
R45175 VCC.n4822 VCC.n4821 2.10336
R45176 VCC.n4701 VCC.n4700 2.10336
R45177 VCC.n5252 VCC.n5251 2.10336
R45178 VCC.n5374 VCC.n5373 2.10336
R45179 VCC.n5931 VCC.n5930 2.10336
R45180 VCC.n5810 VCC.n5809 2.10336
R45181 VCC.n6361 VCC.n6360 2.10336
R45182 VCC.n6483 VCC.n6482 2.10336
R45183 VCC.n7040 VCC.n7039 2.10336
R45184 VCC.n6919 VCC.n6918 2.10336
R45185 VCC.n7470 VCC.n7469 2.10336
R45186 VCC.n7592 VCC.n7591 2.10336
R45187 VCC.n8149 VCC.n8148 2.10336
R45188 VCC.n8028 VCC.n8027 2.10336
R45189 VCC.n8701 VCC.n8700 2.10336
R45190 VCC.n8579 VCC.n8578 2.10336
R45191 VCC.n9258 VCC.n9257 2.10336
R45192 VCC.n9137 VCC.n9136 2.10336
R45193 VCC.n9688 VCC.n9687 2.10336
R45194 VCC.n9810 VCC.n9809 2.10336
R45195 VCC.n10366 VCC.n10365 2.10336
R45196 VCC.n10245 VCC.n10244 2.10336
R45197 VCC.n10795 VCC.n10794 2.10336
R45198 VCC.n10917 VCC.n10916 2.10336
R45199 VCC.n11473 VCC.n11472 2.10336
R45200 VCC.n11352 VCC.n11351 2.10336
R45201 VCC.n11902 VCC.n11901 2.10336
R45202 VCC.n12024 VCC.n12023 2.10336
R45203 VCC.n12580 VCC.n12579 2.10336
R45204 VCC.n12459 VCC.n12458 2.10336
R45205 VCC.n13009 VCC.n13008 2.10336
R45206 VCC.n13131 VCC.n13130 2.10336
R45207 VCC.n13687 VCC.n13686 2.10336
R45208 VCC.n13566 VCC.n13565 2.10336
R45209 VCC.n14116 VCC.n14115 2.10336
R45210 VCC.n14238 VCC.n14237 2.10336
R45211 VCC.n14794 VCC.n14793 2.10336
R45212 VCC.n14673 VCC.n14672 2.10336
R45213 VCC.n15223 VCC.n15222 2.10336
R45214 VCC.n15345 VCC.n15344 2.10336
R45215 VCC.n15901 VCC.n15900 2.10336
R45216 VCC.n15780 VCC.n15779 2.10336
R45217 VCC.n16330 VCC.n16329 2.10336
R45218 VCC.n16452 VCC.n16451 2.10336
R45219 VCC.n17008 VCC.n17007 2.10336
R45220 VCC.n16887 VCC.n16886 2.10336
R45221 VCC.n17372 VCC.n17371 2.10336
R45222 VCC.n264 VCC.n155 2.01193
R45223 VCC.n385 VCC.n384 2.01193
R45224 VCC.n816 VCC.n707 2.01193
R45225 VCC.n937 VCC.n936 2.01193
R45226 VCC.n1494 VCC.n1493 2.01193
R45227 VCC.n1374 VCC.n1265 2.01193
R45228 VCC.n1925 VCC.n1816 2.01193
R45229 VCC.n2046 VCC.n2045 2.01193
R45230 VCC.n2603 VCC.n2602 2.01193
R45231 VCC.n2483 VCC.n2374 2.01193
R45232 VCC.n3034 VCC.n2925 2.01193
R45233 VCC.n3155 VCC.n3154 2.01193
R45234 VCC.n3712 VCC.n3711 2.01193
R45235 VCC.n3592 VCC.n3483 2.01193
R45236 VCC.n4143 VCC.n4034 2.01193
R45237 VCC.n4264 VCC.n4263 2.01193
R45238 VCC.n4821 VCC.n4820 2.01193
R45239 VCC.n4701 VCC.n4592 2.01193
R45240 VCC.n5252 VCC.n5143 2.01193
R45241 VCC.n5373 VCC.n5372 2.01193
R45242 VCC.n5930 VCC.n5929 2.01193
R45243 VCC.n5810 VCC.n5701 2.01193
R45244 VCC.n6361 VCC.n6252 2.01193
R45245 VCC.n6482 VCC.n6481 2.01193
R45246 VCC.n7039 VCC.n7038 2.01193
R45247 VCC.n6919 VCC.n6810 2.01193
R45248 VCC.n7470 VCC.n7361 2.01193
R45249 VCC.n7591 VCC.n7590 2.01193
R45250 VCC.n8148 VCC.n8147 2.01193
R45251 VCC.n8028 VCC.n7919 2.01193
R45252 VCC.n8700 VCC.n8699 2.01193
R45253 VCC.n8579 VCC.n8470 2.01193
R45254 VCC.n9257 VCC.n9256 2.01193
R45255 VCC.n9137 VCC.n9028 2.01193
R45256 VCC.n9688 VCC.n9579 2.01193
R45257 VCC.n9809 VCC.n9808 2.01193
R45258 VCC.n10365 VCC.n10364 2.01193
R45259 VCC.n10245 VCC.n10136 2.01193
R45260 VCC.n10795 VCC.n10686 2.01193
R45261 VCC.n10916 VCC.n10915 2.01193
R45262 VCC.n11472 VCC.n11471 2.01193
R45263 VCC.n11352 VCC.n11243 2.01193
R45264 VCC.n11902 VCC.n11793 2.01193
R45265 VCC.n12023 VCC.n12022 2.01193
R45266 VCC.n12579 VCC.n12578 2.01193
R45267 VCC.n12459 VCC.n12350 2.01193
R45268 VCC.n13009 VCC.n12900 2.01193
R45269 VCC.n13130 VCC.n13129 2.01193
R45270 VCC.n13686 VCC.n13685 2.01193
R45271 VCC.n13566 VCC.n13457 2.01193
R45272 VCC.n14116 VCC.n14007 2.01193
R45273 VCC.n14237 VCC.n14236 2.01193
R45274 VCC.n14793 VCC.n14792 2.01193
R45275 VCC.n14673 VCC.n14564 2.01193
R45276 VCC.n15223 VCC.n15114 2.01193
R45277 VCC.n15344 VCC.n15343 2.01193
R45278 VCC.n15900 VCC.n15899 2.01193
R45279 VCC.n15780 VCC.n15671 2.01193
R45280 VCC.n16330 VCC.n16221 2.01193
R45281 VCC.n16451 VCC.n16450 2.01193
R45282 VCC.n17007 VCC.n17006 2.01193
R45283 VCC.n16887 VCC.n16778 2.01193
R45284 VCC.n17371 VCC.n17370 2.01193
R45285 VCC.n550 VCC.n549 2.00996
R45286 VCC.n1104 VCC.n1103 2.00996
R45287 VCC.n1658 VCC.n1657 2.00996
R45288 VCC.n2213 VCC.n2212 2.00996
R45289 VCC.n2767 VCC.n2766 2.00996
R45290 VCC.n3322 VCC.n3321 2.00996
R45291 VCC.n3876 VCC.n3875 2.00996
R45292 VCC.n4431 VCC.n4430 2.00996
R45293 VCC.n4985 VCC.n4984 2.00996
R45294 VCC.n5540 VCC.n5539 2.00996
R45295 VCC.n6094 VCC.n6093 2.00996
R45296 VCC.n6649 VCC.n6648 2.00996
R45297 VCC.n7203 VCC.n7202 2.00996
R45298 VCC.n7758 VCC.n7757 2.00996
R45299 VCC.n8312 VCC.n8311 2.00996
R45300 VCC.n8867 VCC.n8866 2.00996
R45301 VCC.n9421 VCC.n9420 2.00996
R45302 VCC.n9976 VCC.n9975 2.00996
R45303 VCC.n10529 VCC.n10528 2.00996
R45304 VCC.n11083 VCC.n11082 2.00996
R45305 VCC.n11636 VCC.n11635 2.00996
R45306 VCC.n12190 VCC.n12189 2.00996
R45307 VCC.n12743 VCC.n12742 2.00996
R45308 VCC.n13297 VCC.n13296 2.00996
R45309 VCC.n13850 VCC.n13849 2.00996
R45310 VCC.n14404 VCC.n14403 2.00996
R45311 VCC.n14957 VCC.n14956 2.00996
R45312 VCC.n15511 VCC.n15510 2.00996
R45313 VCC.n16064 VCC.n16063 2.00996
R45314 VCC.n16618 VCC.n16617 2.00996
R45315 VCC.n17171 VCC.n17170 2.00996
R45316 VCC.n17538 VCC.n17537 2.00996
R45317 VCC VCC.n2216 1.98947
R45318 VCC VCC.n6652 1.98947
R45319 VCC.n17552 VCC 1.98947
R45320 VCC.n17544 VCC 1.98947
R45321 VCC.n451 VCC.n65 1.98102
R45322 VCC.n1003 VCC.n617 1.98102
R45323 VCC.n2112 VCC.n1726 1.98102
R45324 VCC.n3221 VCC.n2835 1.98102
R45325 VCC.n4330 VCC.n3944 1.98102
R45326 VCC.n5439 VCC.n5053 1.98102
R45327 VCC.n6548 VCC.n6162 1.98102
R45328 VCC.n7657 VCC.n7271 1.98102
R45329 VCC.n8766 VCC.n8380 1.98102
R45330 VCC.n9875 VCC.n9489 1.98102
R45331 VCC.n10982 VCC.n10596 1.98102
R45332 VCC.n12089 VCC.n11703 1.98102
R45333 VCC.n13196 VCC.n12810 1.98102
R45334 VCC.n14303 VCC.n13917 1.98102
R45335 VCC.n15410 VCC.n15024 1.98102
R45336 VCC.n16517 VCC.n16131 1.98102
R45337 VCC.n17437 VCC.n17238 1.98102
R45338 VCC.n1561 VCC.n1174 1.98071
R45339 VCC.n2670 VCC.n2283 1.98071
R45340 VCC.n3779 VCC.n3392 1.98071
R45341 VCC.n4888 VCC.n4501 1.98071
R45342 VCC.n5997 VCC.n5610 1.98071
R45343 VCC.n7106 VCC.n6719 1.98071
R45344 VCC.n8215 VCC.n7828 1.98071
R45345 VCC.n9324 VCC.n8937 1.98071
R45346 VCC.n10432 VCC.n10045 1.98071
R45347 VCC.n11539 VCC.n11152 1.98071
R45348 VCC.n12646 VCC.n12259 1.98071
R45349 VCC.n13753 VCC.n13366 1.98071
R45350 VCC.n14860 VCC.n14473 1.98071
R45351 VCC.n15967 VCC.n15580 1.98071
R45352 VCC.n17074 VCC.n16687 1.98071
R45353 VCC.n1107 VCC 1.87918
R45354 VCC.n3325 VCC 1.87918
R45355 VCC.n5543 VCC 1.87918
R45356 VCC.n7761 VCC 1.87918
R45357 VCC VCC.n17554 1.87918
R45358 VCC VCC.n17550 1.87918
R45359 VCC VCC.n17546 1.87918
R45360 VCC VCC.n17542 1.87918
R45361 VCC.n229 VCC.n228 1.82742
R45362 VCC.n268 VCC.n142 1.82742
R45363 VCC.n361 VCC.n360 1.82742
R45364 VCC.n396 VCC.n395 1.82742
R45365 VCC.n781 VCC.n780 1.82742
R45366 VCC.n820 VCC.n694 1.82742
R45367 VCC.n913 VCC.n912 1.82742
R45368 VCC.n948 VCC.n947 1.82742
R45369 VCC.n1470 VCC.n1469 1.82742
R45370 VCC.n1505 VCC.n1504 1.82742
R45371 VCC.n1339 VCC.n1338 1.82742
R45372 VCC.n1378 VCC.n1252 1.82742
R45373 VCC.n1890 VCC.n1889 1.82742
R45374 VCC.n1929 VCC.n1803 1.82742
R45375 VCC.n2022 VCC.n2021 1.82742
R45376 VCC.n2057 VCC.n2056 1.82742
R45377 VCC.n2579 VCC.n2578 1.82742
R45378 VCC.n2614 VCC.n2613 1.82742
R45379 VCC.n2448 VCC.n2447 1.82742
R45380 VCC.n2487 VCC.n2361 1.82742
R45381 VCC.n2999 VCC.n2998 1.82742
R45382 VCC.n3038 VCC.n2912 1.82742
R45383 VCC.n3131 VCC.n3130 1.82742
R45384 VCC.n3166 VCC.n3165 1.82742
R45385 VCC.n3688 VCC.n3687 1.82742
R45386 VCC.n3723 VCC.n3722 1.82742
R45387 VCC.n3557 VCC.n3556 1.82742
R45388 VCC.n3596 VCC.n3470 1.82742
R45389 VCC.n4108 VCC.n4107 1.82742
R45390 VCC.n4147 VCC.n4021 1.82742
R45391 VCC.n4240 VCC.n4239 1.82742
R45392 VCC.n4275 VCC.n4274 1.82742
R45393 VCC.n4797 VCC.n4796 1.82742
R45394 VCC.n4832 VCC.n4831 1.82742
R45395 VCC.n4666 VCC.n4665 1.82742
R45396 VCC.n4705 VCC.n4579 1.82742
R45397 VCC.n5217 VCC.n5216 1.82742
R45398 VCC.n5256 VCC.n5130 1.82742
R45399 VCC.n5349 VCC.n5348 1.82742
R45400 VCC.n5384 VCC.n5383 1.82742
R45401 VCC.n5906 VCC.n5905 1.82742
R45402 VCC.n5941 VCC.n5940 1.82742
R45403 VCC.n5775 VCC.n5774 1.82742
R45404 VCC.n5814 VCC.n5688 1.82742
R45405 VCC.n6326 VCC.n6325 1.82742
R45406 VCC.n6365 VCC.n6239 1.82742
R45407 VCC.n6458 VCC.n6457 1.82742
R45408 VCC.n6493 VCC.n6492 1.82742
R45409 VCC.n7015 VCC.n7014 1.82742
R45410 VCC.n7050 VCC.n7049 1.82742
R45411 VCC.n6884 VCC.n6883 1.82742
R45412 VCC.n6923 VCC.n6797 1.82742
R45413 VCC.n7435 VCC.n7434 1.82742
R45414 VCC.n7474 VCC.n7348 1.82742
R45415 VCC.n7567 VCC.n7566 1.82742
R45416 VCC.n7602 VCC.n7601 1.82742
R45417 VCC.n8124 VCC.n8123 1.82742
R45418 VCC.n8159 VCC.n8158 1.82742
R45419 VCC.n7993 VCC.n7992 1.82742
R45420 VCC.n8032 VCC.n7906 1.82742
R45421 VCC.n8676 VCC.n8675 1.82742
R45422 VCC.n8711 VCC.n8710 1.82742
R45423 VCC.n8544 VCC.n8543 1.82742
R45424 VCC.n8583 VCC.n8457 1.82742
R45425 VCC.n9233 VCC.n9232 1.82742
R45426 VCC.n9268 VCC.n9267 1.82742
R45427 VCC.n9102 VCC.n9101 1.82742
R45428 VCC.n9141 VCC.n9015 1.82742
R45429 VCC.n9653 VCC.n9652 1.82742
R45430 VCC.n9692 VCC.n9566 1.82742
R45431 VCC.n9785 VCC.n9784 1.82742
R45432 VCC.n9820 VCC.n9819 1.82742
R45433 VCC.n10341 VCC.n10340 1.82742
R45434 VCC.n10376 VCC.n10375 1.82742
R45435 VCC.n10210 VCC.n10209 1.82742
R45436 VCC.n10249 VCC.n10123 1.82742
R45437 VCC.n10760 VCC.n10759 1.82742
R45438 VCC.n10799 VCC.n10673 1.82742
R45439 VCC.n10892 VCC.n10891 1.82742
R45440 VCC.n10927 VCC.n10926 1.82742
R45441 VCC.n11448 VCC.n11447 1.82742
R45442 VCC.n11483 VCC.n11482 1.82742
R45443 VCC.n11317 VCC.n11316 1.82742
R45444 VCC.n11356 VCC.n11230 1.82742
R45445 VCC.n11867 VCC.n11866 1.82742
R45446 VCC.n11906 VCC.n11780 1.82742
R45447 VCC.n11999 VCC.n11998 1.82742
R45448 VCC.n12034 VCC.n12033 1.82742
R45449 VCC.n12555 VCC.n12554 1.82742
R45450 VCC.n12590 VCC.n12589 1.82742
R45451 VCC.n12424 VCC.n12423 1.82742
R45452 VCC.n12463 VCC.n12337 1.82742
R45453 VCC.n12974 VCC.n12973 1.82742
R45454 VCC.n13013 VCC.n12887 1.82742
R45455 VCC.n13106 VCC.n13105 1.82742
R45456 VCC.n13141 VCC.n13140 1.82742
R45457 VCC.n13662 VCC.n13661 1.82742
R45458 VCC.n13697 VCC.n13696 1.82742
R45459 VCC.n13531 VCC.n13530 1.82742
R45460 VCC.n13570 VCC.n13444 1.82742
R45461 VCC.n14081 VCC.n14080 1.82742
R45462 VCC.n14120 VCC.n13994 1.82742
R45463 VCC.n14213 VCC.n14212 1.82742
R45464 VCC.n14248 VCC.n14247 1.82742
R45465 VCC.n14769 VCC.n14768 1.82742
R45466 VCC.n14804 VCC.n14803 1.82742
R45467 VCC.n14638 VCC.n14637 1.82742
R45468 VCC.n14677 VCC.n14551 1.82742
R45469 VCC.n15188 VCC.n15187 1.82742
R45470 VCC.n15227 VCC.n15101 1.82742
R45471 VCC.n15320 VCC.n15319 1.82742
R45472 VCC.n15355 VCC.n15354 1.82742
R45473 VCC.n15876 VCC.n15875 1.82742
R45474 VCC.n15911 VCC.n15910 1.82742
R45475 VCC.n15745 VCC.n15744 1.82742
R45476 VCC.n15784 VCC.n15658 1.82742
R45477 VCC.n16295 VCC.n16294 1.82742
R45478 VCC.n16334 VCC.n16208 1.82742
R45479 VCC.n16427 VCC.n16426 1.82742
R45480 VCC.n16462 VCC.n16461 1.82742
R45481 VCC.n16983 VCC.n16982 1.82742
R45482 VCC.n17018 VCC.n17017 1.82742
R45483 VCC.n16852 VCC.n16851 1.82742
R45484 VCC.n16891 VCC.n16765 1.82742
R45485 VCC.n17347 VCC.n17346 1.82742
R45486 VCC.n17382 VCC.n17381 1.82742
R45487 VCC VCC.n8870 1.82403
R45488 VCC VCC.n4434 1.67697
R45489 VCC.n17548 VCC 1.67697
R45490 VCC.n492 VCC.n42 1.62907
R45491 VCC.n524 VCC.n23 1.62907
R45492 VCC.n1044 VCC.n594 1.62907
R45493 VCC.n1076 VCC.n575 1.62907
R45494 VCC.n1586 VCC.n1162 1.62907
R45495 VCC.n1622 VCC.n1142 1.62907
R45496 VCC.n2153 VCC.n1703 1.62907
R45497 VCC.n2185 VCC.n1684 1.62907
R45498 VCC.n2695 VCC.n2271 1.62907
R45499 VCC.n2731 VCC.n2251 1.62907
R45500 VCC.n3262 VCC.n2812 1.62907
R45501 VCC.n3294 VCC.n2793 1.62907
R45502 VCC.n3804 VCC.n3380 1.62907
R45503 VCC.n3840 VCC.n3360 1.62907
R45504 VCC.n4371 VCC.n3921 1.62907
R45505 VCC.n4403 VCC.n3902 1.62907
R45506 VCC.n4913 VCC.n4489 1.62907
R45507 VCC.n4949 VCC.n4469 1.62907
R45508 VCC.n5480 VCC.n5030 1.62907
R45509 VCC.n5512 VCC.n5011 1.62907
R45510 VCC.n6022 VCC.n5598 1.62907
R45511 VCC.n6058 VCC.n5578 1.62907
R45512 VCC.n6589 VCC.n6139 1.62907
R45513 VCC.n6621 VCC.n6120 1.62907
R45514 VCC.n7131 VCC.n6707 1.62907
R45515 VCC.n7167 VCC.n6687 1.62907
R45516 VCC.n7698 VCC.n7248 1.62907
R45517 VCC.n7730 VCC.n7229 1.62907
R45518 VCC.n8240 VCC.n7816 1.62907
R45519 VCC.n8276 VCC.n7796 1.62907
R45520 VCC.n8807 VCC.n8357 1.62907
R45521 VCC.n8839 VCC.n8338 1.62907
R45522 VCC.n9349 VCC.n8925 1.62907
R45523 VCC.n9385 VCC.n8905 1.62907
R45524 VCC.n9916 VCC.n9466 1.62907
R45525 VCC.n9948 VCC.n9447 1.62907
R45526 VCC.n10457 VCC.n10033 1.62907
R45527 VCC.n10493 VCC.n10013 1.62907
R45528 VCC.n11023 VCC.n10573 1.62907
R45529 VCC.n11055 VCC.n10554 1.62907
R45530 VCC.n11564 VCC.n11140 1.62907
R45531 VCC.n11600 VCC.n11120 1.62907
R45532 VCC.n12130 VCC.n11680 1.62907
R45533 VCC.n12162 VCC.n11661 1.62907
R45534 VCC.n12671 VCC.n12247 1.62907
R45535 VCC.n12707 VCC.n12227 1.62907
R45536 VCC.n13237 VCC.n12787 1.62907
R45537 VCC.n13269 VCC.n12768 1.62907
R45538 VCC.n13778 VCC.n13354 1.62907
R45539 VCC.n13814 VCC.n13334 1.62907
R45540 VCC.n14344 VCC.n13894 1.62907
R45541 VCC.n14376 VCC.n13875 1.62907
R45542 VCC.n14885 VCC.n14461 1.62907
R45543 VCC.n14921 VCC.n14441 1.62907
R45544 VCC.n15451 VCC.n15001 1.62907
R45545 VCC.n15483 VCC.n14982 1.62907
R45546 VCC.n15992 VCC.n15568 1.62907
R45547 VCC.n16028 VCC.n15548 1.62907
R45548 VCC.n16558 VCC.n16108 1.62907
R45549 VCC.n16590 VCC.n16089 1.62907
R45550 VCC.n17099 VCC.n16675 1.62907
R45551 VCC.n17135 VCC.n16655 1.62907
R45552 VCC.n17478 VCC.n17215 1.62907
R45553 VCC.n17510 VCC.n17196 1.62907
R45554 VCC.n468 VCC.n57 1.55479
R45555 VCC.n1020 VCC.n609 1.55479
R45556 VCC.n1577 VCC.n1165 1.55479
R45557 VCC.n2129 VCC.n1718 1.55479
R45558 VCC.n2686 VCC.n2274 1.55479
R45559 VCC.n3238 VCC.n2827 1.55479
R45560 VCC.n3795 VCC.n3383 1.55479
R45561 VCC.n4347 VCC.n3936 1.55479
R45562 VCC.n4904 VCC.n4492 1.55479
R45563 VCC.n5456 VCC.n5045 1.55479
R45564 VCC.n6013 VCC.n5601 1.55479
R45565 VCC.n6565 VCC.n6154 1.55479
R45566 VCC.n7122 VCC.n6710 1.55479
R45567 VCC.n7674 VCC.n7263 1.55479
R45568 VCC.n8231 VCC.n7819 1.55479
R45569 VCC.n8783 VCC.n8372 1.55479
R45570 VCC.n9340 VCC.n8928 1.55479
R45571 VCC.n9892 VCC.n9481 1.55479
R45572 VCC.n10448 VCC.n10036 1.55479
R45573 VCC.n10999 VCC.n10588 1.55479
R45574 VCC.n11555 VCC.n11143 1.55479
R45575 VCC.n12106 VCC.n11695 1.55479
R45576 VCC.n12662 VCC.n12250 1.55479
R45577 VCC.n13213 VCC.n12802 1.55479
R45578 VCC.n13769 VCC.n13357 1.55479
R45579 VCC.n14320 VCC.n13909 1.55479
R45580 VCC.n14876 VCC.n14464 1.55479
R45581 VCC.n15427 VCC.n15016 1.55479
R45582 VCC.n15983 VCC.n15571 1.55479
R45583 VCC.n16534 VCC.n16123 1.55479
R45584 VCC.n17090 VCC.n16678 1.55479
R45585 VCC.n17454 VCC.n17230 1.55479
R45586 VCC.n253 VCC.n252 1.5005
R45587 VCC.n805 VCC.n804 1.5005
R45588 VCC.n1363 VCC.n1362 1.5005
R45589 VCC.n1914 VCC.n1913 1.5005
R45590 VCC.n2472 VCC.n2471 1.5005
R45591 VCC.n3023 VCC.n3022 1.5005
R45592 VCC.n3581 VCC.n3580 1.5005
R45593 VCC.n4132 VCC.n4131 1.5005
R45594 VCC.n4690 VCC.n4689 1.5005
R45595 VCC.n5241 VCC.n5240 1.5005
R45596 VCC.n5799 VCC.n5798 1.5005
R45597 VCC.n6350 VCC.n6349 1.5005
R45598 VCC.n6908 VCC.n6907 1.5005
R45599 VCC.n7459 VCC.n7458 1.5005
R45600 VCC.n8017 VCC.n8016 1.5005
R45601 VCC.n8568 VCC.n8567 1.5005
R45602 VCC.n9126 VCC.n9125 1.5005
R45603 VCC.n9677 VCC.n9676 1.5005
R45604 VCC.n10234 VCC.n10233 1.5005
R45605 VCC.n10784 VCC.n10783 1.5005
R45606 VCC.n11341 VCC.n11340 1.5005
R45607 VCC.n11891 VCC.n11890 1.5005
R45608 VCC.n12448 VCC.n12447 1.5005
R45609 VCC.n12998 VCC.n12997 1.5005
R45610 VCC.n13555 VCC.n13554 1.5005
R45611 VCC.n14105 VCC.n14104 1.5005
R45612 VCC.n14662 VCC.n14661 1.5005
R45613 VCC.n15212 VCC.n15211 1.5005
R45614 VCC.n15769 VCC.n15768 1.5005
R45615 VCC.n16319 VCC.n16318 1.5005
R45616 VCC.n16876 VCC.n16875 1.5005
R45617 VCC.n178 VCC.n169 1.46336
R45618 VCC.n270 VCC.n151 1.46336
R45619 VCC.n364 VCC.n106 1.46336
R45620 VCC.n392 VCC.n91 1.46336
R45621 VCC.n530 VCC.n7 1.46336
R45622 VCC.n730 VCC.n721 1.46336
R45623 VCC.n822 VCC.n703 1.46336
R45624 VCC.n916 VCC.n658 1.46336
R45625 VCC.n944 VCC.n643 1.46336
R45626 VCC.n1082 VCC.n561 1.46336
R45627 VCC.n1123 VCC.n1117 1.46336
R45628 VCC.n1473 VCC.n1215 1.46336
R45629 VCC.n1501 VCC.n1200 1.46336
R45630 VCC.n1288 VCC.n1279 1.46336
R45631 VCC.n1380 VCC.n1261 1.46336
R45632 VCC.n1839 VCC.n1830 1.46336
R45633 VCC.n1931 VCC.n1812 1.46336
R45634 VCC.n2025 VCC.n1767 1.46336
R45635 VCC.n2053 VCC.n1752 1.46336
R45636 VCC.n2191 VCC.n1670 1.46336
R45637 VCC.n2232 VCC.n2226 1.46336
R45638 VCC.n2582 VCC.n2324 1.46336
R45639 VCC.n2610 VCC.n2309 1.46336
R45640 VCC.n2397 VCC.n2388 1.46336
R45641 VCC.n2489 VCC.n2370 1.46336
R45642 VCC.n2948 VCC.n2939 1.46336
R45643 VCC.n3040 VCC.n2921 1.46336
R45644 VCC.n3134 VCC.n2876 1.46336
R45645 VCC.n3162 VCC.n2861 1.46336
R45646 VCC.n3300 VCC.n2779 1.46336
R45647 VCC.n3341 VCC.n3335 1.46336
R45648 VCC.n3691 VCC.n3433 1.46336
R45649 VCC.n3719 VCC.n3418 1.46336
R45650 VCC.n3506 VCC.n3497 1.46336
R45651 VCC.n3598 VCC.n3479 1.46336
R45652 VCC.n4057 VCC.n4048 1.46336
R45653 VCC.n4149 VCC.n4030 1.46336
R45654 VCC.n4243 VCC.n3985 1.46336
R45655 VCC.n4271 VCC.n3970 1.46336
R45656 VCC.n4409 VCC.n3888 1.46336
R45657 VCC.n4450 VCC.n4444 1.46336
R45658 VCC.n4800 VCC.n4542 1.46336
R45659 VCC.n4828 VCC.n4527 1.46336
R45660 VCC.n4615 VCC.n4606 1.46336
R45661 VCC.n4707 VCC.n4588 1.46336
R45662 VCC.n5166 VCC.n5157 1.46336
R45663 VCC.n5258 VCC.n5139 1.46336
R45664 VCC.n5352 VCC.n5094 1.46336
R45665 VCC.n5380 VCC.n5079 1.46336
R45666 VCC.n5518 VCC.n4997 1.46336
R45667 VCC.n5559 VCC.n5553 1.46336
R45668 VCC.n5909 VCC.n5651 1.46336
R45669 VCC.n5937 VCC.n5636 1.46336
R45670 VCC.n5724 VCC.n5715 1.46336
R45671 VCC.n5816 VCC.n5697 1.46336
R45672 VCC.n6275 VCC.n6266 1.46336
R45673 VCC.n6367 VCC.n6248 1.46336
R45674 VCC.n6461 VCC.n6203 1.46336
R45675 VCC.n6489 VCC.n6188 1.46336
R45676 VCC.n6627 VCC.n6106 1.46336
R45677 VCC.n6668 VCC.n6662 1.46336
R45678 VCC.n7018 VCC.n6760 1.46336
R45679 VCC.n7046 VCC.n6745 1.46336
R45680 VCC.n6833 VCC.n6824 1.46336
R45681 VCC.n6925 VCC.n6806 1.46336
R45682 VCC.n7384 VCC.n7375 1.46336
R45683 VCC.n7476 VCC.n7357 1.46336
R45684 VCC.n7570 VCC.n7312 1.46336
R45685 VCC.n7598 VCC.n7297 1.46336
R45686 VCC.n7736 VCC.n7215 1.46336
R45687 VCC.n7777 VCC.n7771 1.46336
R45688 VCC.n8127 VCC.n7869 1.46336
R45689 VCC.n8155 VCC.n7854 1.46336
R45690 VCC.n7942 VCC.n7933 1.46336
R45691 VCC.n8034 VCC.n7915 1.46336
R45692 VCC.n8679 VCC.n8421 1.46336
R45693 VCC.n8707 VCC.n8406 1.46336
R45694 VCC.n8845 VCC.n8324 1.46336
R45695 VCC.n8493 VCC.n8484 1.46336
R45696 VCC.n8585 VCC.n8466 1.46336
R45697 VCC.n8886 VCC.n8880 1.46336
R45698 VCC.n9236 VCC.n8978 1.46336
R45699 VCC.n9264 VCC.n8963 1.46336
R45700 VCC.n9051 VCC.n9042 1.46336
R45701 VCC.n9143 VCC.n9024 1.46336
R45702 VCC.n9602 VCC.n9593 1.46336
R45703 VCC.n9694 VCC.n9575 1.46336
R45704 VCC.n9788 VCC.n9530 1.46336
R45705 VCC.n9816 VCC.n9515 1.46336
R45706 VCC.n9954 VCC.n9433 1.46336
R45707 VCC.n9994 VCC.n9988 1.46336
R45708 VCC.n10344 VCC.n10086 1.46336
R45709 VCC.n10372 VCC.n10071 1.46336
R45710 VCC.n10159 VCC.n10150 1.46336
R45711 VCC.n10251 VCC.n10132 1.46336
R45712 VCC.n10709 VCC.n10700 1.46336
R45713 VCC.n10801 VCC.n10682 1.46336
R45714 VCC.n10895 VCC.n10637 1.46336
R45715 VCC.n10923 VCC.n10622 1.46336
R45716 VCC.n11061 VCC.n10540 1.46336
R45717 VCC.n11101 VCC.n11095 1.46336
R45718 VCC.n11451 VCC.n11193 1.46336
R45719 VCC.n11479 VCC.n11178 1.46336
R45720 VCC.n11266 VCC.n11257 1.46336
R45721 VCC.n11358 VCC.n11239 1.46336
R45722 VCC.n11816 VCC.n11807 1.46336
R45723 VCC.n11908 VCC.n11789 1.46336
R45724 VCC.n12002 VCC.n11744 1.46336
R45725 VCC.n12030 VCC.n11729 1.46336
R45726 VCC.n12168 VCC.n11647 1.46336
R45727 VCC.n12208 VCC.n12202 1.46336
R45728 VCC.n12558 VCC.n12300 1.46336
R45729 VCC.n12586 VCC.n12285 1.46336
R45730 VCC.n12373 VCC.n12364 1.46336
R45731 VCC.n12465 VCC.n12346 1.46336
R45732 VCC.n12923 VCC.n12914 1.46336
R45733 VCC.n13015 VCC.n12896 1.46336
R45734 VCC.n13109 VCC.n12851 1.46336
R45735 VCC.n13137 VCC.n12836 1.46336
R45736 VCC.n13275 VCC.n12754 1.46336
R45737 VCC.n13315 VCC.n13309 1.46336
R45738 VCC.n13665 VCC.n13407 1.46336
R45739 VCC.n13693 VCC.n13392 1.46336
R45740 VCC.n13480 VCC.n13471 1.46336
R45741 VCC.n13572 VCC.n13453 1.46336
R45742 VCC.n14030 VCC.n14021 1.46336
R45743 VCC.n14122 VCC.n14003 1.46336
R45744 VCC.n14216 VCC.n13958 1.46336
R45745 VCC.n14244 VCC.n13943 1.46336
R45746 VCC.n14382 VCC.n13861 1.46336
R45747 VCC.n14422 VCC.n14416 1.46336
R45748 VCC.n14772 VCC.n14514 1.46336
R45749 VCC.n14800 VCC.n14499 1.46336
R45750 VCC.n14587 VCC.n14578 1.46336
R45751 VCC.n14679 VCC.n14560 1.46336
R45752 VCC.n15137 VCC.n15128 1.46336
R45753 VCC.n15229 VCC.n15110 1.46336
R45754 VCC.n15323 VCC.n15065 1.46336
R45755 VCC.n15351 VCC.n15050 1.46336
R45756 VCC.n15489 VCC.n14968 1.46336
R45757 VCC.n15529 VCC.n15523 1.46336
R45758 VCC.n15879 VCC.n15621 1.46336
R45759 VCC.n15907 VCC.n15606 1.46336
R45760 VCC.n15694 VCC.n15685 1.46336
R45761 VCC.n15786 VCC.n15667 1.46336
R45762 VCC.n16244 VCC.n16235 1.46336
R45763 VCC.n16336 VCC.n16217 1.46336
R45764 VCC.n16430 VCC.n16172 1.46336
R45765 VCC.n16458 VCC.n16157 1.46336
R45766 VCC.n16596 VCC.n16075 1.46336
R45767 VCC.n16636 VCC.n16630 1.46336
R45768 VCC.n16986 VCC.n16728 1.46336
R45769 VCC.n17014 VCC.n16713 1.46336
R45770 VCC.n16801 VCC.n16792 1.46336
R45771 VCC.n16893 VCC.n16774 1.46336
R45772 VCC.n17350 VCC.n17279 1.46336
R45773 VCC.n17378 VCC.n17264 1.46336
R45774 VCC.n17516 VCC.n17182 1.46336
R45775 VCC.n476 VCC.n43 1.37193
R45776 VCC.n491 VCC.n39 1.37193
R45777 VCC.n498 VCC.n24 1.37193
R45778 VCC.n515 VCC.n25 1.37193
R45779 VCC.n1028 VCC.n595 1.37193
R45780 VCC.n1043 VCC.n591 1.37193
R45781 VCC.n1050 VCC.n576 1.37193
R45782 VCC.n1067 VCC.n577 1.37193
R45783 VCC.n1594 VCC.n1593 1.37193
R45784 VCC.n1160 VCC.n1145 1.37193
R45785 VCC.n1617 VCC.n1135 1.37193
R45786 VCC.n1141 VCC.n1140 1.37193
R45787 VCC.n2137 VCC.n1704 1.37193
R45788 VCC.n2152 VCC.n1700 1.37193
R45789 VCC.n2159 VCC.n1685 1.37193
R45790 VCC.n2176 VCC.n1686 1.37193
R45791 VCC.n2703 VCC.n2702 1.37193
R45792 VCC.n2269 VCC.n2254 1.37193
R45793 VCC.n2726 VCC.n2244 1.37193
R45794 VCC.n2250 VCC.n2249 1.37193
R45795 VCC.n3246 VCC.n2813 1.37193
R45796 VCC.n3261 VCC.n2809 1.37193
R45797 VCC.n3268 VCC.n2794 1.37193
R45798 VCC.n3285 VCC.n2795 1.37193
R45799 VCC.n3812 VCC.n3811 1.37193
R45800 VCC.n3378 VCC.n3363 1.37193
R45801 VCC.n3835 VCC.n3353 1.37193
R45802 VCC.n3359 VCC.n3358 1.37193
R45803 VCC.n4355 VCC.n3922 1.37193
R45804 VCC.n4370 VCC.n3918 1.37193
R45805 VCC.n4377 VCC.n3903 1.37193
R45806 VCC.n4394 VCC.n3904 1.37193
R45807 VCC.n4921 VCC.n4920 1.37193
R45808 VCC.n4487 VCC.n4472 1.37193
R45809 VCC.n4944 VCC.n4462 1.37193
R45810 VCC.n4468 VCC.n4467 1.37193
R45811 VCC.n5464 VCC.n5031 1.37193
R45812 VCC.n5479 VCC.n5027 1.37193
R45813 VCC.n5486 VCC.n5012 1.37193
R45814 VCC.n5503 VCC.n5013 1.37193
R45815 VCC.n6030 VCC.n6029 1.37193
R45816 VCC.n5596 VCC.n5581 1.37193
R45817 VCC.n6053 VCC.n5571 1.37193
R45818 VCC.n5577 VCC.n5576 1.37193
R45819 VCC.n6573 VCC.n6140 1.37193
R45820 VCC.n6588 VCC.n6136 1.37193
R45821 VCC.n6595 VCC.n6121 1.37193
R45822 VCC.n6612 VCC.n6122 1.37193
R45823 VCC.n7139 VCC.n7138 1.37193
R45824 VCC.n6705 VCC.n6690 1.37193
R45825 VCC.n7162 VCC.n6680 1.37193
R45826 VCC.n6686 VCC.n6685 1.37193
R45827 VCC.n7682 VCC.n7249 1.37193
R45828 VCC.n7697 VCC.n7245 1.37193
R45829 VCC.n7704 VCC.n7230 1.37193
R45830 VCC.n7721 VCC.n7231 1.37193
R45831 VCC.n8248 VCC.n8247 1.37193
R45832 VCC.n7814 VCC.n7799 1.37193
R45833 VCC.n8271 VCC.n7789 1.37193
R45834 VCC.n7795 VCC.n7794 1.37193
R45835 VCC.n8791 VCC.n8358 1.37193
R45836 VCC.n8806 VCC.n8354 1.37193
R45837 VCC.n8813 VCC.n8339 1.37193
R45838 VCC.n8830 VCC.n8340 1.37193
R45839 VCC.n9357 VCC.n9356 1.37193
R45840 VCC.n8923 VCC.n8908 1.37193
R45841 VCC.n9380 VCC.n8898 1.37193
R45842 VCC.n8904 VCC.n8903 1.37193
R45843 VCC.n9900 VCC.n9467 1.37193
R45844 VCC.n9915 VCC.n9463 1.37193
R45845 VCC.n9922 VCC.n9448 1.37193
R45846 VCC.n9939 VCC.n9449 1.37193
R45847 VCC.n10465 VCC.n10464 1.37193
R45848 VCC.n10031 VCC.n10016 1.37193
R45849 VCC.n10488 VCC.n10006 1.37193
R45850 VCC.n10012 VCC.n10011 1.37193
R45851 VCC.n11007 VCC.n10574 1.37193
R45852 VCC.n11022 VCC.n10570 1.37193
R45853 VCC.n11029 VCC.n10555 1.37193
R45854 VCC.n11046 VCC.n10556 1.37193
R45855 VCC.n11572 VCC.n11571 1.37193
R45856 VCC.n11138 VCC.n11123 1.37193
R45857 VCC.n11595 VCC.n11113 1.37193
R45858 VCC.n11119 VCC.n11118 1.37193
R45859 VCC.n12114 VCC.n11681 1.37193
R45860 VCC.n12129 VCC.n11677 1.37193
R45861 VCC.n12136 VCC.n11662 1.37193
R45862 VCC.n12153 VCC.n11663 1.37193
R45863 VCC.n12679 VCC.n12678 1.37193
R45864 VCC.n12245 VCC.n12230 1.37193
R45865 VCC.n12702 VCC.n12220 1.37193
R45866 VCC.n12226 VCC.n12225 1.37193
R45867 VCC.n13221 VCC.n12788 1.37193
R45868 VCC.n13236 VCC.n12784 1.37193
R45869 VCC.n13243 VCC.n12769 1.37193
R45870 VCC.n13260 VCC.n12770 1.37193
R45871 VCC.n13786 VCC.n13785 1.37193
R45872 VCC.n13352 VCC.n13337 1.37193
R45873 VCC.n13809 VCC.n13327 1.37193
R45874 VCC.n13333 VCC.n13332 1.37193
R45875 VCC.n14328 VCC.n13895 1.37193
R45876 VCC.n14343 VCC.n13891 1.37193
R45877 VCC.n14350 VCC.n13876 1.37193
R45878 VCC.n14367 VCC.n13877 1.37193
R45879 VCC.n14893 VCC.n14892 1.37193
R45880 VCC.n14459 VCC.n14444 1.37193
R45881 VCC.n14916 VCC.n14434 1.37193
R45882 VCC.n14440 VCC.n14439 1.37193
R45883 VCC.n15435 VCC.n15002 1.37193
R45884 VCC.n15450 VCC.n14998 1.37193
R45885 VCC.n15457 VCC.n14983 1.37193
R45886 VCC.n15474 VCC.n14984 1.37193
R45887 VCC.n16000 VCC.n15999 1.37193
R45888 VCC.n15566 VCC.n15551 1.37193
R45889 VCC.n16023 VCC.n15541 1.37193
R45890 VCC.n15547 VCC.n15546 1.37193
R45891 VCC.n16542 VCC.n16109 1.37193
R45892 VCC.n16557 VCC.n16105 1.37193
R45893 VCC.n16564 VCC.n16090 1.37193
R45894 VCC.n16581 VCC.n16091 1.37193
R45895 VCC.n17107 VCC.n17106 1.37193
R45896 VCC.n16673 VCC.n16658 1.37193
R45897 VCC.n17130 VCC.n16648 1.37193
R45898 VCC.n16654 VCC.n16653 1.37193
R45899 VCC.n17462 VCC.n17216 1.37193
R45900 VCC.n17477 VCC.n17212 1.37193
R45901 VCC.n17484 VCC.n17197 1.37193
R45902 VCC.n17501 VCC.n17198 1.37193
R45903 VCC.n224 VCC.n223 1.2805
R45904 VCC.n287 VCC.n286 1.2805
R45905 VCC.n341 VCC.n339 1.2805
R45906 VCC.n415 VCC.n413 1.2805
R45907 VCC.n776 VCC.n775 1.2805
R45908 VCC.n839 VCC.n838 1.2805
R45909 VCC.n893 VCC.n891 1.2805
R45910 VCC.n967 VCC.n965 1.2805
R45911 VCC.n1450 VCC.n1448 1.2805
R45912 VCC.n1524 VCC.n1522 1.2805
R45913 VCC.n1334 VCC.n1333 1.2805
R45914 VCC.n1397 VCC.n1396 1.2805
R45915 VCC.n1885 VCC.n1884 1.2805
R45916 VCC.n1948 VCC.n1947 1.2805
R45917 VCC.n2002 VCC.n2000 1.2805
R45918 VCC.n2076 VCC.n2074 1.2805
R45919 VCC.n2559 VCC.n2557 1.2805
R45920 VCC.n2633 VCC.n2631 1.2805
R45921 VCC.n2443 VCC.n2442 1.2805
R45922 VCC.n2506 VCC.n2505 1.2805
R45923 VCC.n2994 VCC.n2993 1.2805
R45924 VCC.n3057 VCC.n3056 1.2805
R45925 VCC.n3111 VCC.n3109 1.2805
R45926 VCC.n3185 VCC.n3183 1.2805
R45927 VCC.n3668 VCC.n3666 1.2805
R45928 VCC.n3742 VCC.n3740 1.2805
R45929 VCC.n3552 VCC.n3551 1.2805
R45930 VCC.n3615 VCC.n3614 1.2805
R45931 VCC.n4103 VCC.n4102 1.2805
R45932 VCC.n4166 VCC.n4165 1.2805
R45933 VCC.n4220 VCC.n4218 1.2805
R45934 VCC.n4294 VCC.n4292 1.2805
R45935 VCC.n4777 VCC.n4775 1.2805
R45936 VCC.n4851 VCC.n4849 1.2805
R45937 VCC.n4661 VCC.n4660 1.2805
R45938 VCC.n4724 VCC.n4723 1.2805
R45939 VCC.n5212 VCC.n5211 1.2805
R45940 VCC.n5275 VCC.n5274 1.2805
R45941 VCC.n5329 VCC.n5327 1.2805
R45942 VCC.n5403 VCC.n5401 1.2805
R45943 VCC.n5886 VCC.n5884 1.2805
R45944 VCC.n5960 VCC.n5958 1.2805
R45945 VCC.n5770 VCC.n5769 1.2805
R45946 VCC.n5833 VCC.n5832 1.2805
R45947 VCC.n6321 VCC.n6320 1.2805
R45948 VCC.n6384 VCC.n6383 1.2805
R45949 VCC.n6438 VCC.n6436 1.2805
R45950 VCC.n6512 VCC.n6510 1.2805
R45951 VCC.n6995 VCC.n6993 1.2805
R45952 VCC.n7069 VCC.n7067 1.2805
R45953 VCC.n6879 VCC.n6878 1.2805
R45954 VCC.n6942 VCC.n6941 1.2805
R45955 VCC.n7430 VCC.n7429 1.2805
R45956 VCC.n7493 VCC.n7492 1.2805
R45957 VCC.n7547 VCC.n7545 1.2805
R45958 VCC.n7621 VCC.n7619 1.2805
R45959 VCC.n8104 VCC.n8102 1.2805
R45960 VCC.n8178 VCC.n8176 1.2805
R45961 VCC.n7988 VCC.n7987 1.2805
R45962 VCC.n8051 VCC.n8050 1.2805
R45963 VCC.n8656 VCC.n8654 1.2805
R45964 VCC.n8730 VCC.n8728 1.2805
R45965 VCC.n8539 VCC.n8538 1.2805
R45966 VCC.n8602 VCC.n8601 1.2805
R45967 VCC.n9213 VCC.n9211 1.2805
R45968 VCC.n9287 VCC.n9285 1.2805
R45969 VCC.n9097 VCC.n9096 1.2805
R45970 VCC.n9160 VCC.n9159 1.2805
R45971 VCC.n9648 VCC.n9647 1.2805
R45972 VCC.n9711 VCC.n9710 1.2805
R45973 VCC.n9765 VCC.n9763 1.2805
R45974 VCC.n9839 VCC.n9837 1.2805
R45975 VCC.n10321 VCC.n10319 1.2805
R45976 VCC.n10395 VCC.n10393 1.2805
R45977 VCC.n10205 VCC.n10204 1.2805
R45978 VCC.n10268 VCC.n10267 1.2805
R45979 VCC.n10755 VCC.n10754 1.2805
R45980 VCC.n10818 VCC.n10817 1.2805
R45981 VCC.n10872 VCC.n10870 1.2805
R45982 VCC.n10946 VCC.n10944 1.2805
R45983 VCC.n11428 VCC.n11426 1.2805
R45984 VCC.n11502 VCC.n11500 1.2805
R45985 VCC.n11312 VCC.n11311 1.2805
R45986 VCC.n11375 VCC.n11374 1.2805
R45987 VCC.n11862 VCC.n11861 1.2805
R45988 VCC.n11925 VCC.n11924 1.2805
R45989 VCC.n11979 VCC.n11977 1.2805
R45990 VCC.n12053 VCC.n12051 1.2805
R45991 VCC.n12535 VCC.n12533 1.2805
R45992 VCC.n12609 VCC.n12607 1.2805
R45993 VCC.n12419 VCC.n12418 1.2805
R45994 VCC.n12482 VCC.n12481 1.2805
R45995 VCC.n12969 VCC.n12968 1.2805
R45996 VCC.n13032 VCC.n13031 1.2805
R45997 VCC.n13086 VCC.n13084 1.2805
R45998 VCC.n13160 VCC.n13158 1.2805
R45999 VCC.n13642 VCC.n13640 1.2805
R46000 VCC.n13716 VCC.n13714 1.2805
R46001 VCC.n13526 VCC.n13525 1.2805
R46002 VCC.n13589 VCC.n13588 1.2805
R46003 VCC.n14076 VCC.n14075 1.2805
R46004 VCC.n14139 VCC.n14138 1.2805
R46005 VCC.n14193 VCC.n14191 1.2805
R46006 VCC.n14267 VCC.n14265 1.2805
R46007 VCC.n14749 VCC.n14747 1.2805
R46008 VCC.n14823 VCC.n14821 1.2805
R46009 VCC.n14633 VCC.n14632 1.2805
R46010 VCC.n14696 VCC.n14695 1.2805
R46011 VCC.n15183 VCC.n15182 1.2805
R46012 VCC.n15246 VCC.n15245 1.2805
R46013 VCC.n15300 VCC.n15298 1.2805
R46014 VCC.n15374 VCC.n15372 1.2805
R46015 VCC.n15856 VCC.n15854 1.2805
R46016 VCC.n15930 VCC.n15928 1.2805
R46017 VCC.n15740 VCC.n15739 1.2805
R46018 VCC.n15803 VCC.n15802 1.2805
R46019 VCC.n16290 VCC.n16289 1.2805
R46020 VCC.n16353 VCC.n16352 1.2805
R46021 VCC.n16407 VCC.n16405 1.2805
R46022 VCC.n16481 VCC.n16479 1.2805
R46023 VCC.n16963 VCC.n16961 1.2805
R46024 VCC.n17037 VCC.n17035 1.2805
R46025 VCC.n16847 VCC.n16846 1.2805
R46026 VCC.n16910 VCC.n16909 1.2805
R46027 VCC.n17327 VCC.n17325 1.2805
R46028 VCC.n17401 VCC.n17399 1.2805
R46029 VCC.n475 VCC.n54 1.18907
R46030 VCC.n529 VCC.n20 1.18907
R46031 VCC.n1027 VCC.n606 1.18907
R46032 VCC.n1081 VCC.n572 1.18907
R46033 VCC.n1578 VCC.n1159 1.18907
R46034 VCC.n1649 VCC.n1116 1.18907
R46035 VCC.n2136 VCC.n1715 1.18907
R46036 VCC.n2190 VCC.n1681 1.18907
R46037 VCC.n2687 VCC.n2268 1.18907
R46038 VCC.n2758 VCC.n2225 1.18907
R46039 VCC.n3245 VCC.n2824 1.18907
R46040 VCC.n3299 VCC.n2790 1.18907
R46041 VCC.n3796 VCC.n3377 1.18907
R46042 VCC.n3867 VCC.n3334 1.18907
R46043 VCC.n4354 VCC.n3933 1.18907
R46044 VCC.n4408 VCC.n3899 1.18907
R46045 VCC.n4905 VCC.n4486 1.18907
R46046 VCC.n4976 VCC.n4443 1.18907
R46047 VCC.n5463 VCC.n5042 1.18907
R46048 VCC.n5517 VCC.n5008 1.18907
R46049 VCC.n6014 VCC.n5595 1.18907
R46050 VCC.n6085 VCC.n5552 1.18907
R46051 VCC.n6572 VCC.n6151 1.18907
R46052 VCC.n6626 VCC.n6117 1.18907
R46053 VCC.n7123 VCC.n6704 1.18907
R46054 VCC.n7194 VCC.n6661 1.18907
R46055 VCC.n7681 VCC.n7260 1.18907
R46056 VCC.n7735 VCC.n7226 1.18907
R46057 VCC.n8232 VCC.n7813 1.18907
R46058 VCC.n8303 VCC.n7770 1.18907
R46059 VCC.n8790 VCC.n8369 1.18907
R46060 VCC.n8844 VCC.n8335 1.18907
R46061 VCC.n9341 VCC.n8922 1.18907
R46062 VCC.n9412 VCC.n8879 1.18907
R46063 VCC.n9899 VCC.n9478 1.18907
R46064 VCC.n9953 VCC.n9444 1.18907
R46065 VCC.n10449 VCC.n10030 1.18907
R46066 VCC.n10520 VCC.n9987 1.18907
R46067 VCC.n11006 VCC.n10585 1.18907
R46068 VCC.n11060 VCC.n10551 1.18907
R46069 VCC.n11556 VCC.n11137 1.18907
R46070 VCC.n11627 VCC.n11094 1.18907
R46071 VCC.n12113 VCC.n11692 1.18907
R46072 VCC.n12167 VCC.n11658 1.18907
R46073 VCC.n12663 VCC.n12244 1.18907
R46074 VCC.n12734 VCC.n12201 1.18907
R46075 VCC.n13220 VCC.n12799 1.18907
R46076 VCC.n13274 VCC.n12765 1.18907
R46077 VCC.n13770 VCC.n13351 1.18907
R46078 VCC.n13841 VCC.n13308 1.18907
R46079 VCC.n14327 VCC.n13906 1.18907
R46080 VCC.n14381 VCC.n13872 1.18907
R46081 VCC.n14877 VCC.n14458 1.18907
R46082 VCC.n14948 VCC.n14415 1.18907
R46083 VCC.n15434 VCC.n15013 1.18907
R46084 VCC.n15488 VCC.n14979 1.18907
R46085 VCC.n15984 VCC.n15565 1.18907
R46086 VCC.n16055 VCC.n15522 1.18907
R46087 VCC.n16541 VCC.n16120 1.18907
R46088 VCC.n16595 VCC.n16086 1.18907
R46089 VCC.n17091 VCC.n16672 1.18907
R46090 VCC.n17162 VCC.n16629 1.18907
R46091 VCC.n17461 VCC.n17227 1.18907
R46092 VCC.n17515 VCC.n17193 1.18907
R46093 VCC.n1 VCC.n0 1.13717
R46094 VCC.n189 VCC.n188 1.13717
R46095 VCC.n187 VCC.n173 1.13717
R46096 VCC.n244 VCC.n243 1.13717
R46097 VCC.n164 VCC.n147 1.13717
R46098 VCC.n132 VCC.n131 1.13717
R46099 VCC.n128 VCC.n127 1.13717
R46100 VCC.n316 VCC.n126 1.13717
R46101 VCC.n346 VCC.n345 1.13717
R46102 VCC.n370 VCC.n369 1.13717
R46103 VCC.n373 VCC.n87 1.13717
R46104 VCC.n71 VCC.n70 1.13717
R46105 VCC.n67 VCC.n66 1.13717
R46106 VCC.n63 VCC.n62 1.13717
R46107 VCC.n61 VCC.n49 1.13717
R46108 VCC.n484 VCC.n483 1.13717
R46109 VCC.n34 VCC.n30 1.13717
R46110 VCC.n14 VCC.n13 1.13717
R46111 VCC.n741 VCC.n740 1.13717
R46112 VCC.n739 VCC.n725 1.13717
R46113 VCC.n796 VCC.n795 1.13717
R46114 VCC.n716 VCC.n699 1.13717
R46115 VCC.n684 VCC.n683 1.13717
R46116 VCC.n680 VCC.n679 1.13717
R46117 VCC.n868 VCC.n678 1.13717
R46118 VCC.n898 VCC.n897 1.13717
R46119 VCC.n922 VCC.n921 1.13717
R46120 VCC.n925 VCC.n639 1.13717
R46121 VCC.n623 VCC.n622 1.13717
R46122 VCC.n619 VCC.n618 1.13717
R46123 VCC.n615 VCC.n614 1.13717
R46124 VCC.n613 VCC.n601 1.13717
R46125 VCC.n1036 VCC.n1035 1.13717
R46126 VCC.n586 VCC.n582 1.13717
R46127 VCC.n566 VCC.n565 1.13717
R46128 VCC.n555 VCC.n554 1.13717
R46129 VCC.n1299 VCC.n1298 1.13717
R46130 VCC.n1297 VCC.n1283 1.13717
R46131 VCC.n1354 VCC.n1353 1.13717
R46132 VCC.n1274 VCC.n1257 1.13717
R46133 VCC.n1242 VCC.n1241 1.13717
R46134 VCC.n1238 VCC.n1237 1.13717
R46135 VCC.n1426 VCC.n1236 1.13717
R46136 VCC.n1170 VCC.n1154 1.13717
R46137 VCC.n1602 VCC.n1601 1.13717
R46138 VCC.n1609 VCC.n1130 1.13717
R46139 VCC.n1127 VCC.n1126 1.13717
R46140 VCC.n1109 VCC.n1108 1.13717
R46141 VCC.n1172 VCC.n1171 1.13717
R46142 VCC.n1455 VCC.n1454 1.13717
R46143 VCC.n1479 VCC.n1478 1.13717
R46144 VCC.n1482 VCC.n1196 1.13717
R46145 VCC.n1180 VCC.n1179 1.13717
R46146 VCC.n1176 VCC.n1175 1.13717
R46147 VCC.n1850 VCC.n1849 1.13717
R46148 VCC.n1848 VCC.n1834 1.13717
R46149 VCC.n1905 VCC.n1904 1.13717
R46150 VCC.n1825 VCC.n1808 1.13717
R46151 VCC.n1793 VCC.n1792 1.13717
R46152 VCC.n1789 VCC.n1788 1.13717
R46153 VCC.n1977 VCC.n1787 1.13717
R46154 VCC.n2007 VCC.n2006 1.13717
R46155 VCC.n2031 VCC.n2030 1.13717
R46156 VCC.n2034 VCC.n1748 1.13717
R46157 VCC.n1732 VCC.n1731 1.13717
R46158 VCC.n1728 VCC.n1727 1.13717
R46159 VCC.n1724 VCC.n1723 1.13717
R46160 VCC.n1722 VCC.n1710 1.13717
R46161 VCC.n2145 VCC.n2144 1.13717
R46162 VCC.n1695 VCC.n1691 1.13717
R46163 VCC.n1675 VCC.n1674 1.13717
R46164 VCC.n1664 VCC.n1663 1.13717
R46165 VCC.n2408 VCC.n2407 1.13717
R46166 VCC.n2406 VCC.n2392 1.13717
R46167 VCC.n2463 VCC.n2462 1.13717
R46168 VCC.n2383 VCC.n2366 1.13717
R46169 VCC.n2351 VCC.n2350 1.13717
R46170 VCC.n2347 VCC.n2346 1.13717
R46171 VCC.n2535 VCC.n2345 1.13717
R46172 VCC.n2279 VCC.n2263 1.13717
R46173 VCC.n2711 VCC.n2710 1.13717
R46174 VCC.n2718 VCC.n2239 1.13717
R46175 VCC.n2236 VCC.n2235 1.13717
R46176 VCC.n2218 VCC.n2217 1.13717
R46177 VCC.n2281 VCC.n2280 1.13717
R46178 VCC.n2564 VCC.n2563 1.13717
R46179 VCC.n2588 VCC.n2587 1.13717
R46180 VCC.n2591 VCC.n2305 1.13717
R46181 VCC.n2289 VCC.n2288 1.13717
R46182 VCC.n2285 VCC.n2284 1.13717
R46183 VCC.n2959 VCC.n2958 1.13717
R46184 VCC.n2957 VCC.n2943 1.13717
R46185 VCC.n3014 VCC.n3013 1.13717
R46186 VCC.n2934 VCC.n2917 1.13717
R46187 VCC.n2902 VCC.n2901 1.13717
R46188 VCC.n2898 VCC.n2897 1.13717
R46189 VCC.n3086 VCC.n2896 1.13717
R46190 VCC.n3116 VCC.n3115 1.13717
R46191 VCC.n3140 VCC.n3139 1.13717
R46192 VCC.n3143 VCC.n2857 1.13717
R46193 VCC.n2841 VCC.n2840 1.13717
R46194 VCC.n2837 VCC.n2836 1.13717
R46195 VCC.n2833 VCC.n2832 1.13717
R46196 VCC.n2831 VCC.n2819 1.13717
R46197 VCC.n3254 VCC.n3253 1.13717
R46198 VCC.n2804 VCC.n2800 1.13717
R46199 VCC.n2784 VCC.n2783 1.13717
R46200 VCC.n2773 VCC.n2772 1.13717
R46201 VCC.n3517 VCC.n3516 1.13717
R46202 VCC.n3515 VCC.n3501 1.13717
R46203 VCC.n3572 VCC.n3571 1.13717
R46204 VCC.n3492 VCC.n3475 1.13717
R46205 VCC.n3460 VCC.n3459 1.13717
R46206 VCC.n3456 VCC.n3455 1.13717
R46207 VCC.n3644 VCC.n3454 1.13717
R46208 VCC.n3388 VCC.n3372 1.13717
R46209 VCC.n3820 VCC.n3819 1.13717
R46210 VCC.n3827 VCC.n3348 1.13717
R46211 VCC.n3345 VCC.n3344 1.13717
R46212 VCC.n3327 VCC.n3326 1.13717
R46213 VCC.n3390 VCC.n3389 1.13717
R46214 VCC.n3673 VCC.n3672 1.13717
R46215 VCC.n3697 VCC.n3696 1.13717
R46216 VCC.n3700 VCC.n3414 1.13717
R46217 VCC.n3398 VCC.n3397 1.13717
R46218 VCC.n3394 VCC.n3393 1.13717
R46219 VCC.n4068 VCC.n4067 1.13717
R46220 VCC.n4066 VCC.n4052 1.13717
R46221 VCC.n4123 VCC.n4122 1.13717
R46222 VCC.n4043 VCC.n4026 1.13717
R46223 VCC.n4011 VCC.n4010 1.13717
R46224 VCC.n4007 VCC.n4006 1.13717
R46225 VCC.n4195 VCC.n4005 1.13717
R46226 VCC.n4225 VCC.n4224 1.13717
R46227 VCC.n4249 VCC.n4248 1.13717
R46228 VCC.n4252 VCC.n3966 1.13717
R46229 VCC.n3950 VCC.n3949 1.13717
R46230 VCC.n3946 VCC.n3945 1.13717
R46231 VCC.n3942 VCC.n3941 1.13717
R46232 VCC.n3940 VCC.n3928 1.13717
R46233 VCC.n4363 VCC.n4362 1.13717
R46234 VCC.n3913 VCC.n3909 1.13717
R46235 VCC.n3893 VCC.n3892 1.13717
R46236 VCC.n3882 VCC.n3881 1.13717
R46237 VCC.n4626 VCC.n4625 1.13717
R46238 VCC.n4624 VCC.n4610 1.13717
R46239 VCC.n4681 VCC.n4680 1.13717
R46240 VCC.n4601 VCC.n4584 1.13717
R46241 VCC.n4569 VCC.n4568 1.13717
R46242 VCC.n4565 VCC.n4564 1.13717
R46243 VCC.n4753 VCC.n4563 1.13717
R46244 VCC.n4497 VCC.n4481 1.13717
R46245 VCC.n4929 VCC.n4928 1.13717
R46246 VCC.n4936 VCC.n4457 1.13717
R46247 VCC.n4454 VCC.n4453 1.13717
R46248 VCC.n4436 VCC.n4435 1.13717
R46249 VCC.n4499 VCC.n4498 1.13717
R46250 VCC.n4782 VCC.n4781 1.13717
R46251 VCC.n4806 VCC.n4805 1.13717
R46252 VCC.n4809 VCC.n4523 1.13717
R46253 VCC.n4507 VCC.n4506 1.13717
R46254 VCC.n4503 VCC.n4502 1.13717
R46255 VCC.n5177 VCC.n5176 1.13717
R46256 VCC.n5175 VCC.n5161 1.13717
R46257 VCC.n5232 VCC.n5231 1.13717
R46258 VCC.n5152 VCC.n5135 1.13717
R46259 VCC.n5120 VCC.n5119 1.13717
R46260 VCC.n5116 VCC.n5115 1.13717
R46261 VCC.n5304 VCC.n5114 1.13717
R46262 VCC.n5334 VCC.n5333 1.13717
R46263 VCC.n5358 VCC.n5357 1.13717
R46264 VCC.n5361 VCC.n5075 1.13717
R46265 VCC.n5059 VCC.n5058 1.13717
R46266 VCC.n5055 VCC.n5054 1.13717
R46267 VCC.n5051 VCC.n5050 1.13717
R46268 VCC.n5049 VCC.n5037 1.13717
R46269 VCC.n5472 VCC.n5471 1.13717
R46270 VCC.n5022 VCC.n5018 1.13717
R46271 VCC.n5002 VCC.n5001 1.13717
R46272 VCC.n4991 VCC.n4990 1.13717
R46273 VCC.n5735 VCC.n5734 1.13717
R46274 VCC.n5733 VCC.n5719 1.13717
R46275 VCC.n5790 VCC.n5789 1.13717
R46276 VCC.n5710 VCC.n5693 1.13717
R46277 VCC.n5678 VCC.n5677 1.13717
R46278 VCC.n5674 VCC.n5673 1.13717
R46279 VCC.n5862 VCC.n5672 1.13717
R46280 VCC.n5606 VCC.n5590 1.13717
R46281 VCC.n6038 VCC.n6037 1.13717
R46282 VCC.n6045 VCC.n5566 1.13717
R46283 VCC.n5563 VCC.n5562 1.13717
R46284 VCC.n5545 VCC.n5544 1.13717
R46285 VCC.n5608 VCC.n5607 1.13717
R46286 VCC.n5891 VCC.n5890 1.13717
R46287 VCC.n5915 VCC.n5914 1.13717
R46288 VCC.n5918 VCC.n5632 1.13717
R46289 VCC.n5616 VCC.n5615 1.13717
R46290 VCC.n5612 VCC.n5611 1.13717
R46291 VCC.n6286 VCC.n6285 1.13717
R46292 VCC.n6284 VCC.n6270 1.13717
R46293 VCC.n6341 VCC.n6340 1.13717
R46294 VCC.n6261 VCC.n6244 1.13717
R46295 VCC.n6229 VCC.n6228 1.13717
R46296 VCC.n6225 VCC.n6224 1.13717
R46297 VCC.n6413 VCC.n6223 1.13717
R46298 VCC.n6443 VCC.n6442 1.13717
R46299 VCC.n6467 VCC.n6466 1.13717
R46300 VCC.n6470 VCC.n6184 1.13717
R46301 VCC.n6168 VCC.n6167 1.13717
R46302 VCC.n6164 VCC.n6163 1.13717
R46303 VCC.n6160 VCC.n6159 1.13717
R46304 VCC.n6158 VCC.n6146 1.13717
R46305 VCC.n6581 VCC.n6580 1.13717
R46306 VCC.n6131 VCC.n6127 1.13717
R46307 VCC.n6111 VCC.n6110 1.13717
R46308 VCC.n6100 VCC.n6099 1.13717
R46309 VCC.n6844 VCC.n6843 1.13717
R46310 VCC.n6842 VCC.n6828 1.13717
R46311 VCC.n6899 VCC.n6898 1.13717
R46312 VCC.n6819 VCC.n6802 1.13717
R46313 VCC.n6787 VCC.n6786 1.13717
R46314 VCC.n6783 VCC.n6782 1.13717
R46315 VCC.n6971 VCC.n6781 1.13717
R46316 VCC.n6715 VCC.n6699 1.13717
R46317 VCC.n7147 VCC.n7146 1.13717
R46318 VCC.n7154 VCC.n6675 1.13717
R46319 VCC.n6672 VCC.n6671 1.13717
R46320 VCC.n6654 VCC.n6653 1.13717
R46321 VCC.n6717 VCC.n6716 1.13717
R46322 VCC.n7000 VCC.n6999 1.13717
R46323 VCC.n7024 VCC.n7023 1.13717
R46324 VCC.n7027 VCC.n6741 1.13717
R46325 VCC.n6725 VCC.n6724 1.13717
R46326 VCC.n6721 VCC.n6720 1.13717
R46327 VCC.n7395 VCC.n7394 1.13717
R46328 VCC.n7393 VCC.n7379 1.13717
R46329 VCC.n7450 VCC.n7449 1.13717
R46330 VCC.n7370 VCC.n7353 1.13717
R46331 VCC.n7338 VCC.n7337 1.13717
R46332 VCC.n7334 VCC.n7333 1.13717
R46333 VCC.n7522 VCC.n7332 1.13717
R46334 VCC.n7552 VCC.n7551 1.13717
R46335 VCC.n7576 VCC.n7575 1.13717
R46336 VCC.n7579 VCC.n7293 1.13717
R46337 VCC.n7277 VCC.n7276 1.13717
R46338 VCC.n7273 VCC.n7272 1.13717
R46339 VCC.n7269 VCC.n7268 1.13717
R46340 VCC.n7267 VCC.n7255 1.13717
R46341 VCC.n7690 VCC.n7689 1.13717
R46342 VCC.n7240 VCC.n7236 1.13717
R46343 VCC.n7220 VCC.n7219 1.13717
R46344 VCC.n7209 VCC.n7208 1.13717
R46345 VCC.n7953 VCC.n7952 1.13717
R46346 VCC.n7951 VCC.n7937 1.13717
R46347 VCC.n8008 VCC.n8007 1.13717
R46348 VCC.n7928 VCC.n7911 1.13717
R46349 VCC.n7896 VCC.n7895 1.13717
R46350 VCC.n7892 VCC.n7891 1.13717
R46351 VCC.n8080 VCC.n7890 1.13717
R46352 VCC.n7824 VCC.n7808 1.13717
R46353 VCC.n8256 VCC.n8255 1.13717
R46354 VCC.n8263 VCC.n7784 1.13717
R46355 VCC.n7781 VCC.n7780 1.13717
R46356 VCC.n7763 VCC.n7762 1.13717
R46357 VCC.n7826 VCC.n7825 1.13717
R46358 VCC.n8109 VCC.n8108 1.13717
R46359 VCC.n8133 VCC.n8132 1.13717
R46360 VCC.n8136 VCC.n7850 1.13717
R46361 VCC.n7834 VCC.n7833 1.13717
R46362 VCC.n7830 VCC.n7829 1.13717
R46363 VCC.n8504 VCC.n8503 1.13717
R46364 VCC.n8502 VCC.n8488 1.13717
R46365 VCC.n8559 VCC.n8558 1.13717
R46366 VCC.n8479 VCC.n8462 1.13717
R46367 VCC.n8447 VCC.n8446 1.13717
R46368 VCC.n8443 VCC.n8442 1.13717
R46369 VCC.n8631 VCC.n8441 1.13717
R46370 VCC.n8661 VCC.n8660 1.13717
R46371 VCC.n8685 VCC.n8684 1.13717
R46372 VCC.n8688 VCC.n8402 1.13717
R46373 VCC.n8386 VCC.n8385 1.13717
R46374 VCC.n8382 VCC.n8381 1.13717
R46375 VCC.n8378 VCC.n8377 1.13717
R46376 VCC.n8376 VCC.n8364 1.13717
R46377 VCC.n8799 VCC.n8798 1.13717
R46378 VCC.n8349 VCC.n8345 1.13717
R46379 VCC.n8329 VCC.n8328 1.13717
R46380 VCC.n8318 VCC.n8317 1.13717
R46381 VCC.n9062 VCC.n9061 1.13717
R46382 VCC.n9060 VCC.n9046 1.13717
R46383 VCC.n9117 VCC.n9116 1.13717
R46384 VCC.n9037 VCC.n9020 1.13717
R46385 VCC.n9005 VCC.n9004 1.13717
R46386 VCC.n9001 VCC.n9000 1.13717
R46387 VCC.n9189 VCC.n8999 1.13717
R46388 VCC.n8933 VCC.n8917 1.13717
R46389 VCC.n9365 VCC.n9364 1.13717
R46390 VCC.n9372 VCC.n8893 1.13717
R46391 VCC.n8890 VCC.n8889 1.13717
R46392 VCC.n8872 VCC.n8871 1.13717
R46393 VCC.n8935 VCC.n8934 1.13717
R46394 VCC.n9218 VCC.n9217 1.13717
R46395 VCC.n9242 VCC.n9241 1.13717
R46396 VCC.n9245 VCC.n8959 1.13717
R46397 VCC.n8943 VCC.n8942 1.13717
R46398 VCC.n8939 VCC.n8938 1.13717
R46399 VCC.n9613 VCC.n9612 1.13717
R46400 VCC.n9611 VCC.n9597 1.13717
R46401 VCC.n9668 VCC.n9667 1.13717
R46402 VCC.n9588 VCC.n9571 1.13717
R46403 VCC.n9556 VCC.n9555 1.13717
R46404 VCC.n9552 VCC.n9551 1.13717
R46405 VCC.n9740 VCC.n9550 1.13717
R46406 VCC.n9770 VCC.n9769 1.13717
R46407 VCC.n9794 VCC.n9793 1.13717
R46408 VCC.n9797 VCC.n9511 1.13717
R46409 VCC.n9495 VCC.n9494 1.13717
R46410 VCC.n9491 VCC.n9490 1.13717
R46411 VCC.n9487 VCC.n9486 1.13717
R46412 VCC.n9485 VCC.n9473 1.13717
R46413 VCC.n9908 VCC.n9907 1.13717
R46414 VCC.n9458 VCC.n9454 1.13717
R46415 VCC.n9438 VCC.n9437 1.13717
R46416 VCC.n9427 VCC.n9426 1.13717
R46417 VCC.n10170 VCC.n10169 1.13717
R46418 VCC.n10168 VCC.n10154 1.13717
R46419 VCC.n10225 VCC.n10224 1.13717
R46420 VCC.n10145 VCC.n10128 1.13717
R46421 VCC.n10113 VCC.n10112 1.13717
R46422 VCC.n10109 VCC.n10108 1.13717
R46423 VCC.n10297 VCC.n10107 1.13717
R46424 VCC.n10041 VCC.n10025 1.13717
R46425 VCC.n10473 VCC.n10472 1.13717
R46426 VCC.n10480 VCC.n10001 1.13717
R46427 VCC.n9998 VCC.n9997 1.13717
R46428 VCC.n9980 VCC.n9979 1.13717
R46429 VCC.n10043 VCC.n10042 1.13717
R46430 VCC.n10326 VCC.n10325 1.13717
R46431 VCC.n10350 VCC.n10349 1.13717
R46432 VCC.n10353 VCC.n10067 1.13717
R46433 VCC.n10051 VCC.n10050 1.13717
R46434 VCC.n10047 VCC.n10046 1.13717
R46435 VCC.n10720 VCC.n10719 1.13717
R46436 VCC.n10718 VCC.n10704 1.13717
R46437 VCC.n10775 VCC.n10774 1.13717
R46438 VCC.n10695 VCC.n10678 1.13717
R46439 VCC.n10663 VCC.n10662 1.13717
R46440 VCC.n10659 VCC.n10658 1.13717
R46441 VCC.n10847 VCC.n10657 1.13717
R46442 VCC.n10877 VCC.n10876 1.13717
R46443 VCC.n10901 VCC.n10900 1.13717
R46444 VCC.n10904 VCC.n10618 1.13717
R46445 VCC.n10602 VCC.n10601 1.13717
R46446 VCC.n10598 VCC.n10597 1.13717
R46447 VCC.n10594 VCC.n10593 1.13717
R46448 VCC.n10592 VCC.n10580 1.13717
R46449 VCC.n11015 VCC.n11014 1.13717
R46450 VCC.n10565 VCC.n10561 1.13717
R46451 VCC.n10545 VCC.n10544 1.13717
R46452 VCC.n10534 VCC.n10533 1.13717
R46453 VCC.n11277 VCC.n11276 1.13717
R46454 VCC.n11275 VCC.n11261 1.13717
R46455 VCC.n11332 VCC.n11331 1.13717
R46456 VCC.n11252 VCC.n11235 1.13717
R46457 VCC.n11220 VCC.n11219 1.13717
R46458 VCC.n11216 VCC.n11215 1.13717
R46459 VCC.n11404 VCC.n11214 1.13717
R46460 VCC.n11148 VCC.n11132 1.13717
R46461 VCC.n11580 VCC.n11579 1.13717
R46462 VCC.n11587 VCC.n11108 1.13717
R46463 VCC.n11105 VCC.n11104 1.13717
R46464 VCC.n11087 VCC.n11086 1.13717
R46465 VCC.n11150 VCC.n11149 1.13717
R46466 VCC.n11433 VCC.n11432 1.13717
R46467 VCC.n11457 VCC.n11456 1.13717
R46468 VCC.n11460 VCC.n11174 1.13717
R46469 VCC.n11158 VCC.n11157 1.13717
R46470 VCC.n11154 VCC.n11153 1.13717
R46471 VCC.n11827 VCC.n11826 1.13717
R46472 VCC.n11825 VCC.n11811 1.13717
R46473 VCC.n11882 VCC.n11881 1.13717
R46474 VCC.n11802 VCC.n11785 1.13717
R46475 VCC.n11770 VCC.n11769 1.13717
R46476 VCC.n11766 VCC.n11765 1.13717
R46477 VCC.n11954 VCC.n11764 1.13717
R46478 VCC.n11984 VCC.n11983 1.13717
R46479 VCC.n12008 VCC.n12007 1.13717
R46480 VCC.n12011 VCC.n11725 1.13717
R46481 VCC.n11709 VCC.n11708 1.13717
R46482 VCC.n11705 VCC.n11704 1.13717
R46483 VCC.n11701 VCC.n11700 1.13717
R46484 VCC.n11699 VCC.n11687 1.13717
R46485 VCC.n12122 VCC.n12121 1.13717
R46486 VCC.n11672 VCC.n11668 1.13717
R46487 VCC.n11652 VCC.n11651 1.13717
R46488 VCC.n11641 VCC.n11640 1.13717
R46489 VCC.n12384 VCC.n12383 1.13717
R46490 VCC.n12382 VCC.n12368 1.13717
R46491 VCC.n12439 VCC.n12438 1.13717
R46492 VCC.n12359 VCC.n12342 1.13717
R46493 VCC.n12327 VCC.n12326 1.13717
R46494 VCC.n12323 VCC.n12322 1.13717
R46495 VCC.n12511 VCC.n12321 1.13717
R46496 VCC.n12255 VCC.n12239 1.13717
R46497 VCC.n12687 VCC.n12686 1.13717
R46498 VCC.n12694 VCC.n12215 1.13717
R46499 VCC.n12212 VCC.n12211 1.13717
R46500 VCC.n12194 VCC.n12193 1.13717
R46501 VCC.n12257 VCC.n12256 1.13717
R46502 VCC.n12540 VCC.n12539 1.13717
R46503 VCC.n12564 VCC.n12563 1.13717
R46504 VCC.n12567 VCC.n12281 1.13717
R46505 VCC.n12265 VCC.n12264 1.13717
R46506 VCC.n12261 VCC.n12260 1.13717
R46507 VCC.n12934 VCC.n12933 1.13717
R46508 VCC.n12932 VCC.n12918 1.13717
R46509 VCC.n12989 VCC.n12988 1.13717
R46510 VCC.n12909 VCC.n12892 1.13717
R46511 VCC.n12877 VCC.n12876 1.13717
R46512 VCC.n12873 VCC.n12872 1.13717
R46513 VCC.n13061 VCC.n12871 1.13717
R46514 VCC.n13091 VCC.n13090 1.13717
R46515 VCC.n13115 VCC.n13114 1.13717
R46516 VCC.n13118 VCC.n12832 1.13717
R46517 VCC.n12816 VCC.n12815 1.13717
R46518 VCC.n12812 VCC.n12811 1.13717
R46519 VCC.n12808 VCC.n12807 1.13717
R46520 VCC.n12806 VCC.n12794 1.13717
R46521 VCC.n13229 VCC.n13228 1.13717
R46522 VCC.n12779 VCC.n12775 1.13717
R46523 VCC.n12759 VCC.n12758 1.13717
R46524 VCC.n12748 VCC.n12747 1.13717
R46525 VCC.n13491 VCC.n13490 1.13717
R46526 VCC.n13489 VCC.n13475 1.13717
R46527 VCC.n13546 VCC.n13545 1.13717
R46528 VCC.n13466 VCC.n13449 1.13717
R46529 VCC.n13434 VCC.n13433 1.13717
R46530 VCC.n13430 VCC.n13429 1.13717
R46531 VCC.n13618 VCC.n13428 1.13717
R46532 VCC.n13362 VCC.n13346 1.13717
R46533 VCC.n13794 VCC.n13793 1.13717
R46534 VCC.n13801 VCC.n13322 1.13717
R46535 VCC.n13319 VCC.n13318 1.13717
R46536 VCC.n13301 VCC.n13300 1.13717
R46537 VCC.n13364 VCC.n13363 1.13717
R46538 VCC.n13647 VCC.n13646 1.13717
R46539 VCC.n13671 VCC.n13670 1.13717
R46540 VCC.n13674 VCC.n13388 1.13717
R46541 VCC.n13372 VCC.n13371 1.13717
R46542 VCC.n13368 VCC.n13367 1.13717
R46543 VCC.n14041 VCC.n14040 1.13717
R46544 VCC.n14039 VCC.n14025 1.13717
R46545 VCC.n14096 VCC.n14095 1.13717
R46546 VCC.n14016 VCC.n13999 1.13717
R46547 VCC.n13984 VCC.n13983 1.13717
R46548 VCC.n13980 VCC.n13979 1.13717
R46549 VCC.n14168 VCC.n13978 1.13717
R46550 VCC.n14198 VCC.n14197 1.13717
R46551 VCC.n14222 VCC.n14221 1.13717
R46552 VCC.n14225 VCC.n13939 1.13717
R46553 VCC.n13923 VCC.n13922 1.13717
R46554 VCC.n13919 VCC.n13918 1.13717
R46555 VCC.n13915 VCC.n13914 1.13717
R46556 VCC.n13913 VCC.n13901 1.13717
R46557 VCC.n14336 VCC.n14335 1.13717
R46558 VCC.n13886 VCC.n13882 1.13717
R46559 VCC.n13866 VCC.n13865 1.13717
R46560 VCC.n13855 VCC.n13854 1.13717
R46561 VCC.n14598 VCC.n14597 1.13717
R46562 VCC.n14596 VCC.n14582 1.13717
R46563 VCC.n14653 VCC.n14652 1.13717
R46564 VCC.n14573 VCC.n14556 1.13717
R46565 VCC.n14541 VCC.n14540 1.13717
R46566 VCC.n14537 VCC.n14536 1.13717
R46567 VCC.n14725 VCC.n14535 1.13717
R46568 VCC.n14469 VCC.n14453 1.13717
R46569 VCC.n14901 VCC.n14900 1.13717
R46570 VCC.n14908 VCC.n14429 1.13717
R46571 VCC.n14426 VCC.n14425 1.13717
R46572 VCC.n14408 VCC.n14407 1.13717
R46573 VCC.n14471 VCC.n14470 1.13717
R46574 VCC.n14754 VCC.n14753 1.13717
R46575 VCC.n14778 VCC.n14777 1.13717
R46576 VCC.n14781 VCC.n14495 1.13717
R46577 VCC.n14479 VCC.n14478 1.13717
R46578 VCC.n14475 VCC.n14474 1.13717
R46579 VCC.n15148 VCC.n15147 1.13717
R46580 VCC.n15146 VCC.n15132 1.13717
R46581 VCC.n15203 VCC.n15202 1.13717
R46582 VCC.n15123 VCC.n15106 1.13717
R46583 VCC.n15091 VCC.n15090 1.13717
R46584 VCC.n15087 VCC.n15086 1.13717
R46585 VCC.n15275 VCC.n15085 1.13717
R46586 VCC.n15305 VCC.n15304 1.13717
R46587 VCC.n15329 VCC.n15328 1.13717
R46588 VCC.n15332 VCC.n15046 1.13717
R46589 VCC.n15030 VCC.n15029 1.13717
R46590 VCC.n15026 VCC.n15025 1.13717
R46591 VCC.n15022 VCC.n15021 1.13717
R46592 VCC.n15020 VCC.n15008 1.13717
R46593 VCC.n15443 VCC.n15442 1.13717
R46594 VCC.n14993 VCC.n14989 1.13717
R46595 VCC.n14973 VCC.n14972 1.13717
R46596 VCC.n14962 VCC.n14961 1.13717
R46597 VCC.n15705 VCC.n15704 1.13717
R46598 VCC.n15703 VCC.n15689 1.13717
R46599 VCC.n15760 VCC.n15759 1.13717
R46600 VCC.n15680 VCC.n15663 1.13717
R46601 VCC.n15648 VCC.n15647 1.13717
R46602 VCC.n15644 VCC.n15643 1.13717
R46603 VCC.n15832 VCC.n15642 1.13717
R46604 VCC.n15576 VCC.n15560 1.13717
R46605 VCC.n16008 VCC.n16007 1.13717
R46606 VCC.n16015 VCC.n15536 1.13717
R46607 VCC.n15533 VCC.n15532 1.13717
R46608 VCC.n15515 VCC.n15514 1.13717
R46609 VCC.n15578 VCC.n15577 1.13717
R46610 VCC.n15861 VCC.n15860 1.13717
R46611 VCC.n15885 VCC.n15884 1.13717
R46612 VCC.n15888 VCC.n15602 1.13717
R46613 VCC.n15586 VCC.n15585 1.13717
R46614 VCC.n15582 VCC.n15581 1.13717
R46615 VCC.n16255 VCC.n16254 1.13717
R46616 VCC.n16253 VCC.n16239 1.13717
R46617 VCC.n16310 VCC.n16309 1.13717
R46618 VCC.n16230 VCC.n16213 1.13717
R46619 VCC.n16198 VCC.n16197 1.13717
R46620 VCC.n16194 VCC.n16193 1.13717
R46621 VCC.n16382 VCC.n16192 1.13717
R46622 VCC.n16412 VCC.n16411 1.13717
R46623 VCC.n16436 VCC.n16435 1.13717
R46624 VCC.n16439 VCC.n16153 1.13717
R46625 VCC.n16137 VCC.n16136 1.13717
R46626 VCC.n16133 VCC.n16132 1.13717
R46627 VCC.n16129 VCC.n16128 1.13717
R46628 VCC.n16127 VCC.n16115 1.13717
R46629 VCC.n16550 VCC.n16549 1.13717
R46630 VCC.n16100 VCC.n16096 1.13717
R46631 VCC.n16080 VCC.n16079 1.13717
R46632 VCC.n16069 VCC.n16068 1.13717
R46633 VCC.n16812 VCC.n16811 1.13717
R46634 VCC.n16810 VCC.n16796 1.13717
R46635 VCC.n16867 VCC.n16866 1.13717
R46636 VCC.n16787 VCC.n16770 1.13717
R46637 VCC.n16755 VCC.n16754 1.13717
R46638 VCC.n16751 VCC.n16750 1.13717
R46639 VCC.n16939 VCC.n16749 1.13717
R46640 VCC.n16683 VCC.n16667 1.13717
R46641 VCC.n17115 VCC.n17114 1.13717
R46642 VCC.n17122 VCC.n16643 1.13717
R46643 VCC.n16640 VCC.n16639 1.13717
R46644 VCC.n16622 VCC.n16621 1.13717
R46645 VCC.n16685 VCC.n16684 1.13717
R46646 VCC.n16968 VCC.n16967 1.13717
R46647 VCC.n16992 VCC.n16991 1.13717
R46648 VCC.n16995 VCC.n16709 1.13717
R46649 VCC.n16693 VCC.n16692 1.13717
R46650 VCC.n16689 VCC.n16688 1.13717
R46651 VCC.n17302 VCC.n17299 1.13717
R46652 VCC.n17332 VCC.n17331 1.13717
R46653 VCC.n17356 VCC.n17355 1.13717
R46654 VCC.n17359 VCC.n17260 1.13717
R46655 VCC.n17244 VCC.n17243 1.13717
R46656 VCC.n17240 VCC.n17239 1.13717
R46657 VCC.n17236 VCC.n17235 1.13717
R46658 VCC.n17234 VCC.n17222 1.13717
R46659 VCC.n17470 VCC.n17469 1.13717
R46660 VCC.n17207 VCC.n17203 1.13717
R46661 VCC.n17187 VCC.n17186 1.13717
R46662 VCC.n17176 VCC.n17175 1.13717
R46663 VCC.n376 VCC.n101 1.1255
R46664 VCC.n500 VCC.n37 1.1255
R46665 VCC.n928 VCC.n653 1.1255
R46666 VCC.n1052 VCC.n589 1.1255
R46667 VCC.n1615 VCC.n1147 1.1255
R46668 VCC.n1485 VCC.n1210 1.1255
R46669 VCC.n2037 VCC.n1762 1.1255
R46670 VCC.n2161 VCC.n1698 1.1255
R46671 VCC.n2724 VCC.n2256 1.1255
R46672 VCC.n2594 VCC.n2319 1.1255
R46673 VCC.n3146 VCC.n2871 1.1255
R46674 VCC.n3270 VCC.n2807 1.1255
R46675 VCC.n3833 VCC.n3365 1.1255
R46676 VCC.n3703 VCC.n3428 1.1255
R46677 VCC.n4255 VCC.n3980 1.1255
R46678 VCC.n4379 VCC.n3916 1.1255
R46679 VCC.n4942 VCC.n4474 1.1255
R46680 VCC.n4812 VCC.n4537 1.1255
R46681 VCC.n5364 VCC.n5089 1.1255
R46682 VCC.n5488 VCC.n5025 1.1255
R46683 VCC.n6051 VCC.n5583 1.1255
R46684 VCC.n5921 VCC.n5646 1.1255
R46685 VCC.n6473 VCC.n6198 1.1255
R46686 VCC.n6597 VCC.n6134 1.1255
R46687 VCC.n7160 VCC.n6692 1.1255
R46688 VCC.n7030 VCC.n6755 1.1255
R46689 VCC.n7582 VCC.n7307 1.1255
R46690 VCC.n7706 VCC.n7243 1.1255
R46691 VCC.n8269 VCC.n7801 1.1255
R46692 VCC.n8139 VCC.n7864 1.1255
R46693 VCC.n8691 VCC.n8416 1.1255
R46694 VCC.n8815 VCC.n8352 1.1255
R46695 VCC.n9378 VCC.n8910 1.1255
R46696 VCC.n9248 VCC.n8973 1.1255
R46697 VCC.n9800 VCC.n9525 1.1255
R46698 VCC.n9924 VCC.n9461 1.1255
R46699 VCC.n10486 VCC.n10018 1.1255
R46700 VCC.n10356 VCC.n10081 1.1255
R46701 VCC.n10907 VCC.n10632 1.1255
R46702 VCC.n11031 VCC.n10568 1.1255
R46703 VCC.n11593 VCC.n11125 1.1255
R46704 VCC.n11463 VCC.n11188 1.1255
R46705 VCC.n12014 VCC.n11739 1.1255
R46706 VCC.n12138 VCC.n11675 1.1255
R46707 VCC.n12700 VCC.n12232 1.1255
R46708 VCC.n12570 VCC.n12295 1.1255
R46709 VCC.n13121 VCC.n12846 1.1255
R46710 VCC.n13245 VCC.n12782 1.1255
R46711 VCC.n13807 VCC.n13339 1.1255
R46712 VCC.n13677 VCC.n13402 1.1255
R46713 VCC.n14228 VCC.n13953 1.1255
R46714 VCC.n14352 VCC.n13889 1.1255
R46715 VCC.n14914 VCC.n14446 1.1255
R46716 VCC.n14784 VCC.n14509 1.1255
R46717 VCC.n15335 VCC.n15060 1.1255
R46718 VCC.n15459 VCC.n14996 1.1255
R46719 VCC.n16021 VCC.n15553 1.1255
R46720 VCC.n15891 VCC.n15616 1.1255
R46721 VCC.n16442 VCC.n16167 1.1255
R46722 VCC.n16566 VCC.n16103 1.1255
R46723 VCC.n17128 VCC.n16660 1.1255
R46724 VCC.n16998 VCC.n16723 1.1255
R46725 VCC.n17362 VCC.n17274 1.1255
R46726 VCC.n17486 VCC.n17210 1.1255
R46727 VCC.n213 VCC.n207 1.00621
R46728 VCC.n201 VCC.n195 1.00621
R46729 VCC.n160 VCC.n159 1.00621
R46730 VCC.n333 VCC.n124 1.00621
R46731 VCC.n326 VCC.n325 1.00621
R46732 VCC.n391 VCC.n95 1.00621
R46733 VCC.n422 VCC.n421 1.00621
R46734 VCC.n545 VCC.n3 1.00621
R46735 VCC.n765 VCC.n759 1.00621
R46736 VCC.n753 VCC.n747 1.00621
R46737 VCC.n712 VCC.n711 1.00621
R46738 VCC.n885 VCC.n676 1.00621
R46739 VCC.n878 VCC.n877 1.00621
R46740 VCC.n943 VCC.n647 1.00621
R46741 VCC.n974 VCC.n973 1.00621
R46742 VCC.n1099 VCC.n557 1.00621
R46743 VCC.n1532 VCC.n1531 1.00621
R46744 VCC.n1656 VCC.n1112 1.00621
R46745 VCC.n1442 VCC.n1233 1.00621
R46746 VCC.n1435 VCC.n1434 1.00621
R46747 VCC.n1500 VCC.n1204 1.00621
R46748 VCC.n1323 VCC.n1317 1.00621
R46749 VCC.n1311 VCC.n1305 1.00621
R46750 VCC.n1270 VCC.n1269 1.00621
R46751 VCC.n1874 VCC.n1868 1.00621
R46752 VCC.n1862 VCC.n1856 1.00621
R46753 VCC.n1821 VCC.n1820 1.00621
R46754 VCC.n1994 VCC.n1785 1.00621
R46755 VCC.n1987 VCC.n1986 1.00621
R46756 VCC.n2052 VCC.n1756 1.00621
R46757 VCC.n2083 VCC.n2082 1.00621
R46758 VCC.n2208 VCC.n1666 1.00621
R46759 VCC.n2641 VCC.n2640 1.00621
R46760 VCC.n2765 VCC.n2221 1.00621
R46761 VCC.n2551 VCC.n2342 1.00621
R46762 VCC.n2544 VCC.n2543 1.00621
R46763 VCC.n2609 VCC.n2313 1.00621
R46764 VCC.n2432 VCC.n2426 1.00621
R46765 VCC.n2420 VCC.n2414 1.00621
R46766 VCC.n2379 VCC.n2378 1.00621
R46767 VCC.n2983 VCC.n2977 1.00621
R46768 VCC.n2971 VCC.n2965 1.00621
R46769 VCC.n2930 VCC.n2929 1.00621
R46770 VCC.n3103 VCC.n2894 1.00621
R46771 VCC.n3096 VCC.n3095 1.00621
R46772 VCC.n3161 VCC.n2865 1.00621
R46773 VCC.n3192 VCC.n3191 1.00621
R46774 VCC.n3317 VCC.n2775 1.00621
R46775 VCC.n3750 VCC.n3749 1.00621
R46776 VCC.n3874 VCC.n3330 1.00621
R46777 VCC.n3660 VCC.n3451 1.00621
R46778 VCC.n3653 VCC.n3652 1.00621
R46779 VCC.n3718 VCC.n3422 1.00621
R46780 VCC.n3541 VCC.n3535 1.00621
R46781 VCC.n3529 VCC.n3523 1.00621
R46782 VCC.n3488 VCC.n3487 1.00621
R46783 VCC.n4092 VCC.n4086 1.00621
R46784 VCC.n4080 VCC.n4074 1.00621
R46785 VCC.n4039 VCC.n4038 1.00621
R46786 VCC.n4212 VCC.n4003 1.00621
R46787 VCC.n4205 VCC.n4204 1.00621
R46788 VCC.n4270 VCC.n3974 1.00621
R46789 VCC.n4301 VCC.n4300 1.00621
R46790 VCC.n4426 VCC.n3884 1.00621
R46791 VCC.n4859 VCC.n4858 1.00621
R46792 VCC.n4983 VCC.n4439 1.00621
R46793 VCC.n4769 VCC.n4560 1.00621
R46794 VCC.n4762 VCC.n4761 1.00621
R46795 VCC.n4827 VCC.n4531 1.00621
R46796 VCC.n4650 VCC.n4644 1.00621
R46797 VCC.n4638 VCC.n4632 1.00621
R46798 VCC.n4597 VCC.n4596 1.00621
R46799 VCC.n5201 VCC.n5195 1.00621
R46800 VCC.n5189 VCC.n5183 1.00621
R46801 VCC.n5148 VCC.n5147 1.00621
R46802 VCC.n5321 VCC.n5112 1.00621
R46803 VCC.n5314 VCC.n5313 1.00621
R46804 VCC.n5379 VCC.n5083 1.00621
R46805 VCC.n5410 VCC.n5409 1.00621
R46806 VCC.n5535 VCC.n4993 1.00621
R46807 VCC.n5968 VCC.n5967 1.00621
R46808 VCC.n6092 VCC.n5548 1.00621
R46809 VCC.n5878 VCC.n5669 1.00621
R46810 VCC.n5871 VCC.n5870 1.00621
R46811 VCC.n5936 VCC.n5640 1.00621
R46812 VCC.n5759 VCC.n5753 1.00621
R46813 VCC.n5747 VCC.n5741 1.00621
R46814 VCC.n5706 VCC.n5705 1.00621
R46815 VCC.n6310 VCC.n6304 1.00621
R46816 VCC.n6298 VCC.n6292 1.00621
R46817 VCC.n6257 VCC.n6256 1.00621
R46818 VCC.n6430 VCC.n6221 1.00621
R46819 VCC.n6423 VCC.n6422 1.00621
R46820 VCC.n6488 VCC.n6192 1.00621
R46821 VCC.n6519 VCC.n6518 1.00621
R46822 VCC.n6644 VCC.n6102 1.00621
R46823 VCC.n7077 VCC.n7076 1.00621
R46824 VCC.n7201 VCC.n6657 1.00621
R46825 VCC.n6987 VCC.n6778 1.00621
R46826 VCC.n6980 VCC.n6979 1.00621
R46827 VCC.n7045 VCC.n6749 1.00621
R46828 VCC.n6868 VCC.n6862 1.00621
R46829 VCC.n6856 VCC.n6850 1.00621
R46830 VCC.n6815 VCC.n6814 1.00621
R46831 VCC.n7419 VCC.n7413 1.00621
R46832 VCC.n7407 VCC.n7401 1.00621
R46833 VCC.n7366 VCC.n7365 1.00621
R46834 VCC.n7539 VCC.n7330 1.00621
R46835 VCC.n7532 VCC.n7531 1.00621
R46836 VCC.n7597 VCC.n7301 1.00621
R46837 VCC.n7628 VCC.n7627 1.00621
R46838 VCC.n7753 VCC.n7211 1.00621
R46839 VCC.n8186 VCC.n8185 1.00621
R46840 VCC.n8310 VCC.n7766 1.00621
R46841 VCC.n8096 VCC.n7887 1.00621
R46842 VCC.n8089 VCC.n8088 1.00621
R46843 VCC.n8154 VCC.n7858 1.00621
R46844 VCC.n7977 VCC.n7971 1.00621
R46845 VCC.n7965 VCC.n7959 1.00621
R46846 VCC.n7924 VCC.n7923 1.00621
R46847 VCC.n8648 VCC.n8439 1.00621
R46848 VCC.n8641 VCC.n8640 1.00621
R46849 VCC.n8706 VCC.n8410 1.00621
R46850 VCC.n8737 VCC.n8736 1.00621
R46851 VCC.n8862 VCC.n8320 1.00621
R46852 VCC.n8528 VCC.n8522 1.00621
R46853 VCC.n8516 VCC.n8510 1.00621
R46854 VCC.n8475 VCC.n8474 1.00621
R46855 VCC.n9295 VCC.n9294 1.00621
R46856 VCC.n9419 VCC.n8875 1.00621
R46857 VCC.n9205 VCC.n8996 1.00621
R46858 VCC.n9198 VCC.n9197 1.00621
R46859 VCC.n9263 VCC.n8967 1.00621
R46860 VCC.n9086 VCC.n9080 1.00621
R46861 VCC.n9074 VCC.n9068 1.00621
R46862 VCC.n9033 VCC.n9032 1.00621
R46863 VCC.n9637 VCC.n9631 1.00621
R46864 VCC.n9625 VCC.n9619 1.00621
R46865 VCC.n9584 VCC.n9583 1.00621
R46866 VCC.n9757 VCC.n9548 1.00621
R46867 VCC.n9750 VCC.n9749 1.00621
R46868 VCC.n9815 VCC.n9519 1.00621
R46869 VCC.n9846 VCC.n9845 1.00621
R46870 VCC.n9971 VCC.n9429 1.00621
R46871 VCC.n10403 VCC.n10402 1.00621
R46872 VCC.n10527 VCC.n9983 1.00621
R46873 VCC.n10313 VCC.n10104 1.00621
R46874 VCC.n10306 VCC.n10305 1.00621
R46875 VCC.n10371 VCC.n10075 1.00621
R46876 VCC.n10194 VCC.n10188 1.00621
R46877 VCC.n10182 VCC.n10176 1.00621
R46878 VCC.n10141 VCC.n10140 1.00621
R46879 VCC.n10744 VCC.n10738 1.00621
R46880 VCC.n10732 VCC.n10726 1.00621
R46881 VCC.n10691 VCC.n10690 1.00621
R46882 VCC.n10864 VCC.n10655 1.00621
R46883 VCC.n10857 VCC.n10856 1.00621
R46884 VCC.n10922 VCC.n10626 1.00621
R46885 VCC.n10953 VCC.n10952 1.00621
R46886 VCC.n11078 VCC.n10536 1.00621
R46887 VCC.n11510 VCC.n11509 1.00621
R46888 VCC.n11634 VCC.n11090 1.00621
R46889 VCC.n11420 VCC.n11211 1.00621
R46890 VCC.n11413 VCC.n11412 1.00621
R46891 VCC.n11478 VCC.n11182 1.00621
R46892 VCC.n11301 VCC.n11295 1.00621
R46893 VCC.n11289 VCC.n11283 1.00621
R46894 VCC.n11248 VCC.n11247 1.00621
R46895 VCC.n11851 VCC.n11845 1.00621
R46896 VCC.n11839 VCC.n11833 1.00621
R46897 VCC.n11798 VCC.n11797 1.00621
R46898 VCC.n11971 VCC.n11762 1.00621
R46899 VCC.n11964 VCC.n11963 1.00621
R46900 VCC.n12029 VCC.n11733 1.00621
R46901 VCC.n12060 VCC.n12059 1.00621
R46902 VCC.n12185 VCC.n11643 1.00621
R46903 VCC.n12617 VCC.n12616 1.00621
R46904 VCC.n12741 VCC.n12197 1.00621
R46905 VCC.n12527 VCC.n12318 1.00621
R46906 VCC.n12520 VCC.n12519 1.00621
R46907 VCC.n12585 VCC.n12289 1.00621
R46908 VCC.n12408 VCC.n12402 1.00621
R46909 VCC.n12396 VCC.n12390 1.00621
R46910 VCC.n12355 VCC.n12354 1.00621
R46911 VCC.n12958 VCC.n12952 1.00621
R46912 VCC.n12946 VCC.n12940 1.00621
R46913 VCC.n12905 VCC.n12904 1.00621
R46914 VCC.n13078 VCC.n12869 1.00621
R46915 VCC.n13071 VCC.n13070 1.00621
R46916 VCC.n13136 VCC.n12840 1.00621
R46917 VCC.n13167 VCC.n13166 1.00621
R46918 VCC.n13292 VCC.n12750 1.00621
R46919 VCC.n13724 VCC.n13723 1.00621
R46920 VCC.n13848 VCC.n13304 1.00621
R46921 VCC.n13634 VCC.n13425 1.00621
R46922 VCC.n13627 VCC.n13626 1.00621
R46923 VCC.n13692 VCC.n13396 1.00621
R46924 VCC.n13515 VCC.n13509 1.00621
R46925 VCC.n13503 VCC.n13497 1.00621
R46926 VCC.n13462 VCC.n13461 1.00621
R46927 VCC.n14065 VCC.n14059 1.00621
R46928 VCC.n14053 VCC.n14047 1.00621
R46929 VCC.n14012 VCC.n14011 1.00621
R46930 VCC.n14185 VCC.n13976 1.00621
R46931 VCC.n14178 VCC.n14177 1.00621
R46932 VCC.n14243 VCC.n13947 1.00621
R46933 VCC.n14274 VCC.n14273 1.00621
R46934 VCC.n14399 VCC.n13857 1.00621
R46935 VCC.n14831 VCC.n14830 1.00621
R46936 VCC.n14955 VCC.n14411 1.00621
R46937 VCC.n14741 VCC.n14532 1.00621
R46938 VCC.n14734 VCC.n14733 1.00621
R46939 VCC.n14799 VCC.n14503 1.00621
R46940 VCC.n14622 VCC.n14616 1.00621
R46941 VCC.n14610 VCC.n14604 1.00621
R46942 VCC.n14569 VCC.n14568 1.00621
R46943 VCC.n15172 VCC.n15166 1.00621
R46944 VCC.n15160 VCC.n15154 1.00621
R46945 VCC.n15119 VCC.n15118 1.00621
R46946 VCC.n15292 VCC.n15083 1.00621
R46947 VCC.n15285 VCC.n15284 1.00621
R46948 VCC.n15350 VCC.n15054 1.00621
R46949 VCC.n15381 VCC.n15380 1.00621
R46950 VCC.n15506 VCC.n14964 1.00621
R46951 VCC.n15938 VCC.n15937 1.00621
R46952 VCC.n16062 VCC.n15518 1.00621
R46953 VCC.n15848 VCC.n15639 1.00621
R46954 VCC.n15841 VCC.n15840 1.00621
R46955 VCC.n15906 VCC.n15610 1.00621
R46956 VCC.n15729 VCC.n15723 1.00621
R46957 VCC.n15717 VCC.n15711 1.00621
R46958 VCC.n15676 VCC.n15675 1.00621
R46959 VCC.n16279 VCC.n16273 1.00621
R46960 VCC.n16267 VCC.n16261 1.00621
R46961 VCC.n16226 VCC.n16225 1.00621
R46962 VCC.n16399 VCC.n16190 1.00621
R46963 VCC.n16392 VCC.n16391 1.00621
R46964 VCC.n16457 VCC.n16161 1.00621
R46965 VCC.n16488 VCC.n16487 1.00621
R46966 VCC.n16613 VCC.n16071 1.00621
R46967 VCC.n17045 VCC.n17044 1.00621
R46968 VCC.n17169 VCC.n16625 1.00621
R46969 VCC.n16955 VCC.n16746 1.00621
R46970 VCC.n16948 VCC.n16947 1.00621
R46971 VCC.n17013 VCC.n16717 1.00621
R46972 VCC.n16836 VCC.n16830 1.00621
R46973 VCC.n16824 VCC.n16818 1.00621
R46974 VCC.n16783 VCC.n16782 1.00621
R46975 VCC.n17319 VCC.n17297 1.00621
R46976 VCC.n17312 VCC.n17311 1.00621
R46977 VCC.n17377 VCC.n17268 1.00621
R46978 VCC.n17408 VCC.n17407 1.00621
R46979 VCC.n17533 VCC.n17178 1.00621
R46980 VCC.n230 VCC.n180 0.9505
R46981 VCC.n269 VCC.n143 0.9505
R46982 VCC.n359 VCC.n107 0.9505
R46983 VCC.n397 VCC.n92 0.9505
R46984 VCC.n782 VCC.n732 0.9505
R46985 VCC.n821 VCC.n695 0.9505
R46986 VCC.n911 VCC.n659 0.9505
R46987 VCC.n949 VCC.n644 0.9505
R46988 VCC.n1468 VCC.n1216 0.9505
R46989 VCC.n1506 VCC.n1201 0.9505
R46990 VCC.n1340 VCC.n1290 0.9505
R46991 VCC.n1379 VCC.n1253 0.9505
R46992 VCC.n1891 VCC.n1841 0.9505
R46993 VCC.n1930 VCC.n1804 0.9505
R46994 VCC.n2020 VCC.n1768 0.9505
R46995 VCC.n2058 VCC.n1753 0.9505
R46996 VCC.n2577 VCC.n2325 0.9505
R46997 VCC.n2615 VCC.n2310 0.9505
R46998 VCC.n2449 VCC.n2399 0.9505
R46999 VCC.n2488 VCC.n2362 0.9505
R47000 VCC.n3000 VCC.n2950 0.9505
R47001 VCC.n3039 VCC.n2913 0.9505
R47002 VCC.n3129 VCC.n2877 0.9505
R47003 VCC.n3167 VCC.n2862 0.9505
R47004 VCC.n3686 VCC.n3434 0.9505
R47005 VCC.n3724 VCC.n3419 0.9505
R47006 VCC.n3558 VCC.n3508 0.9505
R47007 VCC.n3597 VCC.n3471 0.9505
R47008 VCC.n4109 VCC.n4059 0.9505
R47009 VCC.n4148 VCC.n4022 0.9505
R47010 VCC.n4238 VCC.n3986 0.9505
R47011 VCC.n4276 VCC.n3971 0.9505
R47012 VCC.n4795 VCC.n4543 0.9505
R47013 VCC.n4833 VCC.n4528 0.9505
R47014 VCC.n4667 VCC.n4617 0.9505
R47015 VCC.n4706 VCC.n4580 0.9505
R47016 VCC.n5218 VCC.n5168 0.9505
R47017 VCC.n5257 VCC.n5131 0.9505
R47018 VCC.n5347 VCC.n5095 0.9505
R47019 VCC.n5385 VCC.n5080 0.9505
R47020 VCC.n5904 VCC.n5652 0.9505
R47021 VCC.n5942 VCC.n5637 0.9505
R47022 VCC.n5776 VCC.n5726 0.9505
R47023 VCC.n5815 VCC.n5689 0.9505
R47024 VCC.n6327 VCC.n6277 0.9505
R47025 VCC.n6366 VCC.n6240 0.9505
R47026 VCC.n6456 VCC.n6204 0.9505
R47027 VCC.n6494 VCC.n6189 0.9505
R47028 VCC.n7013 VCC.n6761 0.9505
R47029 VCC.n7051 VCC.n6746 0.9505
R47030 VCC.n6885 VCC.n6835 0.9505
R47031 VCC.n6924 VCC.n6798 0.9505
R47032 VCC.n7436 VCC.n7386 0.9505
R47033 VCC.n7475 VCC.n7349 0.9505
R47034 VCC.n7565 VCC.n7313 0.9505
R47035 VCC.n7603 VCC.n7298 0.9505
R47036 VCC.n8122 VCC.n7870 0.9505
R47037 VCC.n8160 VCC.n7855 0.9505
R47038 VCC.n7994 VCC.n7944 0.9505
R47039 VCC.n8033 VCC.n7907 0.9505
R47040 VCC.n8674 VCC.n8422 0.9505
R47041 VCC.n8712 VCC.n8407 0.9505
R47042 VCC.n8545 VCC.n8495 0.9505
R47043 VCC.n8584 VCC.n8458 0.9505
R47044 VCC.n9231 VCC.n8979 0.9505
R47045 VCC.n9269 VCC.n8964 0.9505
R47046 VCC.n9103 VCC.n9053 0.9505
R47047 VCC.n9142 VCC.n9016 0.9505
R47048 VCC.n9654 VCC.n9604 0.9505
R47049 VCC.n9693 VCC.n9567 0.9505
R47050 VCC.n9783 VCC.n9531 0.9505
R47051 VCC.n9821 VCC.n9516 0.9505
R47052 VCC.n10339 VCC.n10087 0.9505
R47053 VCC.n10377 VCC.n10072 0.9505
R47054 VCC.n10211 VCC.n10161 0.9505
R47055 VCC.n10250 VCC.n10124 0.9505
R47056 VCC.n10761 VCC.n10711 0.9505
R47057 VCC.n10800 VCC.n10674 0.9505
R47058 VCC.n10890 VCC.n10638 0.9505
R47059 VCC.n10928 VCC.n10623 0.9505
R47060 VCC.n11446 VCC.n11194 0.9505
R47061 VCC.n11484 VCC.n11179 0.9505
R47062 VCC.n11318 VCC.n11268 0.9505
R47063 VCC.n11357 VCC.n11231 0.9505
R47064 VCC.n11868 VCC.n11818 0.9505
R47065 VCC.n11907 VCC.n11781 0.9505
R47066 VCC.n11997 VCC.n11745 0.9505
R47067 VCC.n12035 VCC.n11730 0.9505
R47068 VCC.n12553 VCC.n12301 0.9505
R47069 VCC.n12591 VCC.n12286 0.9505
R47070 VCC.n12425 VCC.n12375 0.9505
R47071 VCC.n12464 VCC.n12338 0.9505
R47072 VCC.n12975 VCC.n12925 0.9505
R47073 VCC.n13014 VCC.n12888 0.9505
R47074 VCC.n13104 VCC.n12852 0.9505
R47075 VCC.n13142 VCC.n12837 0.9505
R47076 VCC.n13660 VCC.n13408 0.9505
R47077 VCC.n13698 VCC.n13393 0.9505
R47078 VCC.n13532 VCC.n13482 0.9505
R47079 VCC.n13571 VCC.n13445 0.9505
R47080 VCC.n14082 VCC.n14032 0.9505
R47081 VCC.n14121 VCC.n13995 0.9505
R47082 VCC.n14211 VCC.n13959 0.9505
R47083 VCC.n14249 VCC.n13944 0.9505
R47084 VCC.n14767 VCC.n14515 0.9505
R47085 VCC.n14805 VCC.n14500 0.9505
R47086 VCC.n14639 VCC.n14589 0.9505
R47087 VCC.n14678 VCC.n14552 0.9505
R47088 VCC.n15189 VCC.n15139 0.9505
R47089 VCC.n15228 VCC.n15102 0.9505
R47090 VCC.n15318 VCC.n15066 0.9505
R47091 VCC.n15356 VCC.n15051 0.9505
R47092 VCC.n15874 VCC.n15622 0.9505
R47093 VCC.n15912 VCC.n15607 0.9505
R47094 VCC.n15746 VCC.n15696 0.9505
R47095 VCC.n15785 VCC.n15659 0.9505
R47096 VCC.n16296 VCC.n16246 0.9505
R47097 VCC.n16335 VCC.n16209 0.9505
R47098 VCC.n16425 VCC.n16173 0.9505
R47099 VCC.n16463 VCC.n16158 0.9505
R47100 VCC.n16981 VCC.n16729 0.9505
R47101 VCC.n17019 VCC.n16714 0.9505
R47102 VCC.n16853 VCC.n16803 0.9505
R47103 VCC.n16892 VCC.n16766 0.9505
R47104 VCC.n17345 VCC.n17280 0.9505
R47105 VCC.n17383 VCC.n17265 0.9505
R47106 VCC.n248 VCC.n247 0.914786
R47107 VCC.n263 VCC.n156 0.914786
R47108 VCC.n297 VCC.n139 0.914786
R47109 VCC.n296 VCC.n295 0.914786
R47110 VCC.n366 VCC.n365 0.914786
R47111 VCC.n384 VCC.n97 0.914786
R47112 VCC.n432 VCC.n78 0.914786
R47113 VCC.n431 VCC.n430 0.914786
R47114 VCC.n800 VCC.n799 0.914786
R47115 VCC.n815 VCC.n708 0.914786
R47116 VCC.n849 VCC.n691 0.914786
R47117 VCC.n848 VCC.n847 0.914786
R47118 VCC.n918 VCC.n917 0.914786
R47119 VCC.n936 VCC.n649 0.914786
R47120 VCC.n984 VCC.n630 0.914786
R47121 VCC.n983 VCC.n982 0.914786
R47122 VCC.n1475 VCC.n1474 0.914786
R47123 VCC.n1493 VCC.n1206 0.914786
R47124 VCC.n1542 VCC.n1187 0.914786
R47125 VCC.n1541 VCC.n1540 0.914786
R47126 VCC.n1358 VCC.n1357 0.914786
R47127 VCC.n1373 VCC.n1266 0.914786
R47128 VCC.n1407 VCC.n1249 0.914786
R47129 VCC.n1406 VCC.n1405 0.914786
R47130 VCC.n1909 VCC.n1908 0.914786
R47131 VCC.n1924 VCC.n1817 0.914786
R47132 VCC.n1958 VCC.n1800 0.914786
R47133 VCC.n1957 VCC.n1956 0.914786
R47134 VCC.n2027 VCC.n2026 0.914786
R47135 VCC.n2045 VCC.n1758 0.914786
R47136 VCC.n2093 VCC.n1739 0.914786
R47137 VCC.n2092 VCC.n2091 0.914786
R47138 VCC.n2584 VCC.n2583 0.914786
R47139 VCC.n2602 VCC.n2315 0.914786
R47140 VCC.n2651 VCC.n2296 0.914786
R47141 VCC.n2650 VCC.n2649 0.914786
R47142 VCC.n2467 VCC.n2466 0.914786
R47143 VCC.n2482 VCC.n2375 0.914786
R47144 VCC.n2516 VCC.n2358 0.914786
R47145 VCC.n2515 VCC.n2514 0.914786
R47146 VCC.n3018 VCC.n3017 0.914786
R47147 VCC.n3033 VCC.n2926 0.914786
R47148 VCC.n3067 VCC.n2909 0.914786
R47149 VCC.n3066 VCC.n3065 0.914786
R47150 VCC.n3136 VCC.n3135 0.914786
R47151 VCC.n3154 VCC.n2867 0.914786
R47152 VCC.n3202 VCC.n2848 0.914786
R47153 VCC.n3201 VCC.n3200 0.914786
R47154 VCC.n3693 VCC.n3692 0.914786
R47155 VCC.n3711 VCC.n3424 0.914786
R47156 VCC.n3760 VCC.n3405 0.914786
R47157 VCC.n3759 VCC.n3758 0.914786
R47158 VCC.n3576 VCC.n3575 0.914786
R47159 VCC.n3591 VCC.n3484 0.914786
R47160 VCC.n3625 VCC.n3467 0.914786
R47161 VCC.n3624 VCC.n3623 0.914786
R47162 VCC.n4127 VCC.n4126 0.914786
R47163 VCC.n4142 VCC.n4035 0.914786
R47164 VCC.n4176 VCC.n4018 0.914786
R47165 VCC.n4175 VCC.n4174 0.914786
R47166 VCC.n4245 VCC.n4244 0.914786
R47167 VCC.n4263 VCC.n3976 0.914786
R47168 VCC.n4311 VCC.n3957 0.914786
R47169 VCC.n4310 VCC.n4309 0.914786
R47170 VCC.n4802 VCC.n4801 0.914786
R47171 VCC.n4820 VCC.n4533 0.914786
R47172 VCC.n4869 VCC.n4514 0.914786
R47173 VCC.n4868 VCC.n4867 0.914786
R47174 VCC.n4685 VCC.n4684 0.914786
R47175 VCC.n4700 VCC.n4593 0.914786
R47176 VCC.n4734 VCC.n4576 0.914786
R47177 VCC.n4733 VCC.n4732 0.914786
R47178 VCC.n5236 VCC.n5235 0.914786
R47179 VCC.n5251 VCC.n5144 0.914786
R47180 VCC.n5285 VCC.n5127 0.914786
R47181 VCC.n5284 VCC.n5283 0.914786
R47182 VCC.n5354 VCC.n5353 0.914786
R47183 VCC.n5372 VCC.n5085 0.914786
R47184 VCC.n5420 VCC.n5066 0.914786
R47185 VCC.n5419 VCC.n5418 0.914786
R47186 VCC.n5911 VCC.n5910 0.914786
R47187 VCC.n5929 VCC.n5642 0.914786
R47188 VCC.n5978 VCC.n5623 0.914786
R47189 VCC.n5977 VCC.n5976 0.914786
R47190 VCC.n5794 VCC.n5793 0.914786
R47191 VCC.n5809 VCC.n5702 0.914786
R47192 VCC.n5843 VCC.n5685 0.914786
R47193 VCC.n5842 VCC.n5841 0.914786
R47194 VCC.n6345 VCC.n6344 0.914786
R47195 VCC.n6360 VCC.n6253 0.914786
R47196 VCC.n6394 VCC.n6236 0.914786
R47197 VCC.n6393 VCC.n6392 0.914786
R47198 VCC.n6463 VCC.n6462 0.914786
R47199 VCC.n6481 VCC.n6194 0.914786
R47200 VCC.n6529 VCC.n6175 0.914786
R47201 VCC.n6528 VCC.n6527 0.914786
R47202 VCC.n7020 VCC.n7019 0.914786
R47203 VCC.n7038 VCC.n6751 0.914786
R47204 VCC.n7087 VCC.n6732 0.914786
R47205 VCC.n7086 VCC.n7085 0.914786
R47206 VCC.n6903 VCC.n6902 0.914786
R47207 VCC.n6918 VCC.n6811 0.914786
R47208 VCC.n6952 VCC.n6794 0.914786
R47209 VCC.n6951 VCC.n6950 0.914786
R47210 VCC.n7454 VCC.n7453 0.914786
R47211 VCC.n7469 VCC.n7362 0.914786
R47212 VCC.n7503 VCC.n7345 0.914786
R47213 VCC.n7502 VCC.n7501 0.914786
R47214 VCC.n7572 VCC.n7571 0.914786
R47215 VCC.n7590 VCC.n7303 0.914786
R47216 VCC.n7638 VCC.n7284 0.914786
R47217 VCC.n7637 VCC.n7636 0.914786
R47218 VCC.n8129 VCC.n8128 0.914786
R47219 VCC.n8147 VCC.n7860 0.914786
R47220 VCC.n8196 VCC.n7841 0.914786
R47221 VCC.n8195 VCC.n8194 0.914786
R47222 VCC.n8012 VCC.n8011 0.914786
R47223 VCC.n8027 VCC.n7920 0.914786
R47224 VCC.n8061 VCC.n7903 0.914786
R47225 VCC.n8060 VCC.n8059 0.914786
R47226 VCC.n8681 VCC.n8680 0.914786
R47227 VCC.n8699 VCC.n8412 0.914786
R47228 VCC.n8747 VCC.n8393 0.914786
R47229 VCC.n8746 VCC.n8745 0.914786
R47230 VCC.n8563 VCC.n8562 0.914786
R47231 VCC.n8578 VCC.n8471 0.914786
R47232 VCC.n8612 VCC.n8454 0.914786
R47233 VCC.n8611 VCC.n8610 0.914786
R47234 VCC.n9238 VCC.n9237 0.914786
R47235 VCC.n9256 VCC.n8969 0.914786
R47236 VCC.n9305 VCC.n8950 0.914786
R47237 VCC.n9304 VCC.n9303 0.914786
R47238 VCC.n9121 VCC.n9120 0.914786
R47239 VCC.n9136 VCC.n9029 0.914786
R47240 VCC.n9170 VCC.n9012 0.914786
R47241 VCC.n9169 VCC.n9168 0.914786
R47242 VCC.n9672 VCC.n9671 0.914786
R47243 VCC.n9687 VCC.n9580 0.914786
R47244 VCC.n9721 VCC.n9563 0.914786
R47245 VCC.n9720 VCC.n9719 0.914786
R47246 VCC.n9790 VCC.n9789 0.914786
R47247 VCC.n9808 VCC.n9521 0.914786
R47248 VCC.n9856 VCC.n9502 0.914786
R47249 VCC.n9855 VCC.n9854 0.914786
R47250 VCC.n10346 VCC.n10345 0.914786
R47251 VCC.n10364 VCC.n10077 0.914786
R47252 VCC.n10413 VCC.n10058 0.914786
R47253 VCC.n10412 VCC.n10411 0.914786
R47254 VCC.n10229 VCC.n10228 0.914786
R47255 VCC.n10244 VCC.n10137 0.914786
R47256 VCC.n10278 VCC.n10120 0.914786
R47257 VCC.n10277 VCC.n10276 0.914786
R47258 VCC.n10779 VCC.n10778 0.914786
R47259 VCC.n10794 VCC.n10687 0.914786
R47260 VCC.n10828 VCC.n10670 0.914786
R47261 VCC.n10827 VCC.n10826 0.914786
R47262 VCC.n10897 VCC.n10896 0.914786
R47263 VCC.n10915 VCC.n10628 0.914786
R47264 VCC.n10963 VCC.n10609 0.914786
R47265 VCC.n10962 VCC.n10961 0.914786
R47266 VCC.n11453 VCC.n11452 0.914786
R47267 VCC.n11471 VCC.n11184 0.914786
R47268 VCC.n11520 VCC.n11165 0.914786
R47269 VCC.n11519 VCC.n11518 0.914786
R47270 VCC.n11336 VCC.n11335 0.914786
R47271 VCC.n11351 VCC.n11244 0.914786
R47272 VCC.n11385 VCC.n11227 0.914786
R47273 VCC.n11384 VCC.n11383 0.914786
R47274 VCC.n11886 VCC.n11885 0.914786
R47275 VCC.n11901 VCC.n11794 0.914786
R47276 VCC.n11935 VCC.n11777 0.914786
R47277 VCC.n11934 VCC.n11933 0.914786
R47278 VCC.n12004 VCC.n12003 0.914786
R47279 VCC.n12022 VCC.n11735 0.914786
R47280 VCC.n12070 VCC.n11716 0.914786
R47281 VCC.n12069 VCC.n12068 0.914786
R47282 VCC.n12560 VCC.n12559 0.914786
R47283 VCC.n12578 VCC.n12291 0.914786
R47284 VCC.n12627 VCC.n12272 0.914786
R47285 VCC.n12626 VCC.n12625 0.914786
R47286 VCC.n12443 VCC.n12442 0.914786
R47287 VCC.n12458 VCC.n12351 0.914786
R47288 VCC.n12492 VCC.n12334 0.914786
R47289 VCC.n12491 VCC.n12490 0.914786
R47290 VCC.n12993 VCC.n12992 0.914786
R47291 VCC.n13008 VCC.n12901 0.914786
R47292 VCC.n13042 VCC.n12884 0.914786
R47293 VCC.n13041 VCC.n13040 0.914786
R47294 VCC.n13111 VCC.n13110 0.914786
R47295 VCC.n13129 VCC.n12842 0.914786
R47296 VCC.n13177 VCC.n12823 0.914786
R47297 VCC.n13176 VCC.n13175 0.914786
R47298 VCC.n13667 VCC.n13666 0.914786
R47299 VCC.n13685 VCC.n13398 0.914786
R47300 VCC.n13734 VCC.n13379 0.914786
R47301 VCC.n13733 VCC.n13732 0.914786
R47302 VCC.n13550 VCC.n13549 0.914786
R47303 VCC.n13565 VCC.n13458 0.914786
R47304 VCC.n13599 VCC.n13441 0.914786
R47305 VCC.n13598 VCC.n13597 0.914786
R47306 VCC.n14100 VCC.n14099 0.914786
R47307 VCC.n14115 VCC.n14008 0.914786
R47308 VCC.n14149 VCC.n13991 0.914786
R47309 VCC.n14148 VCC.n14147 0.914786
R47310 VCC.n14218 VCC.n14217 0.914786
R47311 VCC.n14236 VCC.n13949 0.914786
R47312 VCC.n14284 VCC.n13930 0.914786
R47313 VCC.n14283 VCC.n14282 0.914786
R47314 VCC.n14774 VCC.n14773 0.914786
R47315 VCC.n14792 VCC.n14505 0.914786
R47316 VCC.n14841 VCC.n14486 0.914786
R47317 VCC.n14840 VCC.n14839 0.914786
R47318 VCC.n14657 VCC.n14656 0.914786
R47319 VCC.n14672 VCC.n14565 0.914786
R47320 VCC.n14706 VCC.n14548 0.914786
R47321 VCC.n14705 VCC.n14704 0.914786
R47322 VCC.n15207 VCC.n15206 0.914786
R47323 VCC.n15222 VCC.n15115 0.914786
R47324 VCC.n15256 VCC.n15098 0.914786
R47325 VCC.n15255 VCC.n15254 0.914786
R47326 VCC.n15325 VCC.n15324 0.914786
R47327 VCC.n15343 VCC.n15056 0.914786
R47328 VCC.n15391 VCC.n15037 0.914786
R47329 VCC.n15390 VCC.n15389 0.914786
R47330 VCC.n15881 VCC.n15880 0.914786
R47331 VCC.n15899 VCC.n15612 0.914786
R47332 VCC.n15948 VCC.n15593 0.914786
R47333 VCC.n15947 VCC.n15946 0.914786
R47334 VCC.n15764 VCC.n15763 0.914786
R47335 VCC.n15779 VCC.n15672 0.914786
R47336 VCC.n15813 VCC.n15655 0.914786
R47337 VCC.n15812 VCC.n15811 0.914786
R47338 VCC.n16314 VCC.n16313 0.914786
R47339 VCC.n16329 VCC.n16222 0.914786
R47340 VCC.n16363 VCC.n16205 0.914786
R47341 VCC.n16362 VCC.n16361 0.914786
R47342 VCC.n16432 VCC.n16431 0.914786
R47343 VCC.n16450 VCC.n16163 0.914786
R47344 VCC.n16498 VCC.n16144 0.914786
R47345 VCC.n16497 VCC.n16496 0.914786
R47346 VCC.n16988 VCC.n16987 0.914786
R47347 VCC.n17006 VCC.n16719 0.914786
R47348 VCC.n17055 VCC.n16700 0.914786
R47349 VCC.n17054 VCC.n17053 0.914786
R47350 VCC.n16871 VCC.n16870 0.914786
R47351 VCC.n16886 VCC.n16779 0.914786
R47352 VCC.n16920 VCC.n16762 0.914786
R47353 VCC.n16919 VCC.n16918 0.914786
R47354 VCC.n17352 VCC.n17351 0.914786
R47355 VCC.n17370 VCC.n17270 0.914786
R47356 VCC.n17418 VCC.n17251 0.914786
R47357 VCC.n17417 VCC.n17416 0.914786
R47358 VCC.n223 VCC.n184 0.823357
R47359 VCC.n232 VCC.n177 0.823357
R47360 VCC.n249 VCC.n155 0.823357
R47361 VCC.n285 VCC.n144 0.823357
R47362 VCC.n341 VCC.n340 0.823357
R47363 VCC.n357 VCC.n110 0.823357
R47364 VCC.n387 VCC.n386 0.823357
R47365 VCC.n412 VCC.n84 0.823357
R47366 VCC.n775 VCC.n736 0.823357
R47367 VCC.n784 VCC.n729 0.823357
R47368 VCC.n801 VCC.n707 0.823357
R47369 VCC.n837 VCC.n696 0.823357
R47370 VCC.n893 VCC.n892 0.823357
R47371 VCC.n909 VCC.n662 0.823357
R47372 VCC.n939 VCC.n938 0.823357
R47373 VCC.n964 VCC.n636 0.823357
R47374 VCC.n1450 VCC.n1449 0.823357
R47375 VCC.n1466 VCC.n1219 0.823357
R47376 VCC.n1496 VCC.n1495 0.823357
R47377 VCC.n1521 VCC.n1193 0.823357
R47378 VCC.n1333 VCC.n1294 0.823357
R47379 VCC.n1342 VCC.n1287 0.823357
R47380 VCC.n1359 VCC.n1265 0.823357
R47381 VCC.n1395 VCC.n1254 0.823357
R47382 VCC.n1884 VCC.n1845 0.823357
R47383 VCC.n1893 VCC.n1838 0.823357
R47384 VCC.n1910 VCC.n1816 0.823357
R47385 VCC.n1946 VCC.n1805 0.823357
R47386 VCC.n2002 VCC.n2001 0.823357
R47387 VCC.n2018 VCC.n1771 0.823357
R47388 VCC.n2048 VCC.n2047 0.823357
R47389 VCC.n2073 VCC.n1745 0.823357
R47390 VCC.n2559 VCC.n2558 0.823357
R47391 VCC.n2575 VCC.n2328 0.823357
R47392 VCC.n2605 VCC.n2604 0.823357
R47393 VCC.n2630 VCC.n2302 0.823357
R47394 VCC.n2442 VCC.n2403 0.823357
R47395 VCC.n2451 VCC.n2396 0.823357
R47396 VCC.n2468 VCC.n2374 0.823357
R47397 VCC.n2504 VCC.n2363 0.823357
R47398 VCC.n2993 VCC.n2954 0.823357
R47399 VCC.n3002 VCC.n2947 0.823357
R47400 VCC.n3019 VCC.n2925 0.823357
R47401 VCC.n3055 VCC.n2914 0.823357
R47402 VCC.n3111 VCC.n3110 0.823357
R47403 VCC.n3127 VCC.n2880 0.823357
R47404 VCC.n3157 VCC.n3156 0.823357
R47405 VCC.n3182 VCC.n2854 0.823357
R47406 VCC.n3668 VCC.n3667 0.823357
R47407 VCC.n3684 VCC.n3437 0.823357
R47408 VCC.n3714 VCC.n3713 0.823357
R47409 VCC.n3739 VCC.n3411 0.823357
R47410 VCC.n3551 VCC.n3512 0.823357
R47411 VCC.n3560 VCC.n3505 0.823357
R47412 VCC.n3577 VCC.n3483 0.823357
R47413 VCC.n3613 VCC.n3472 0.823357
R47414 VCC.n4102 VCC.n4063 0.823357
R47415 VCC.n4111 VCC.n4056 0.823357
R47416 VCC.n4128 VCC.n4034 0.823357
R47417 VCC.n4164 VCC.n4023 0.823357
R47418 VCC.n4220 VCC.n4219 0.823357
R47419 VCC.n4236 VCC.n3989 0.823357
R47420 VCC.n4266 VCC.n4265 0.823357
R47421 VCC.n4291 VCC.n3963 0.823357
R47422 VCC.n4777 VCC.n4776 0.823357
R47423 VCC.n4793 VCC.n4546 0.823357
R47424 VCC.n4823 VCC.n4822 0.823357
R47425 VCC.n4848 VCC.n4520 0.823357
R47426 VCC.n4660 VCC.n4621 0.823357
R47427 VCC.n4669 VCC.n4614 0.823357
R47428 VCC.n4686 VCC.n4592 0.823357
R47429 VCC.n4722 VCC.n4581 0.823357
R47430 VCC.n5211 VCC.n5172 0.823357
R47431 VCC.n5220 VCC.n5165 0.823357
R47432 VCC.n5237 VCC.n5143 0.823357
R47433 VCC.n5273 VCC.n5132 0.823357
R47434 VCC.n5329 VCC.n5328 0.823357
R47435 VCC.n5345 VCC.n5098 0.823357
R47436 VCC.n5375 VCC.n5374 0.823357
R47437 VCC.n5400 VCC.n5072 0.823357
R47438 VCC.n5886 VCC.n5885 0.823357
R47439 VCC.n5902 VCC.n5655 0.823357
R47440 VCC.n5932 VCC.n5931 0.823357
R47441 VCC.n5957 VCC.n5629 0.823357
R47442 VCC.n5769 VCC.n5730 0.823357
R47443 VCC.n5778 VCC.n5723 0.823357
R47444 VCC.n5795 VCC.n5701 0.823357
R47445 VCC.n5831 VCC.n5690 0.823357
R47446 VCC.n6320 VCC.n6281 0.823357
R47447 VCC.n6329 VCC.n6274 0.823357
R47448 VCC.n6346 VCC.n6252 0.823357
R47449 VCC.n6382 VCC.n6241 0.823357
R47450 VCC.n6438 VCC.n6437 0.823357
R47451 VCC.n6454 VCC.n6207 0.823357
R47452 VCC.n6484 VCC.n6483 0.823357
R47453 VCC.n6509 VCC.n6181 0.823357
R47454 VCC.n6995 VCC.n6994 0.823357
R47455 VCC.n7011 VCC.n6764 0.823357
R47456 VCC.n7041 VCC.n7040 0.823357
R47457 VCC.n7066 VCC.n6738 0.823357
R47458 VCC.n6878 VCC.n6839 0.823357
R47459 VCC.n6887 VCC.n6832 0.823357
R47460 VCC.n6904 VCC.n6810 0.823357
R47461 VCC.n6940 VCC.n6799 0.823357
R47462 VCC.n7429 VCC.n7390 0.823357
R47463 VCC.n7438 VCC.n7383 0.823357
R47464 VCC.n7455 VCC.n7361 0.823357
R47465 VCC.n7491 VCC.n7350 0.823357
R47466 VCC.n7547 VCC.n7546 0.823357
R47467 VCC.n7563 VCC.n7316 0.823357
R47468 VCC.n7593 VCC.n7592 0.823357
R47469 VCC.n7618 VCC.n7290 0.823357
R47470 VCC.n8104 VCC.n8103 0.823357
R47471 VCC.n8120 VCC.n7873 0.823357
R47472 VCC.n8150 VCC.n8149 0.823357
R47473 VCC.n8175 VCC.n7847 0.823357
R47474 VCC.n7987 VCC.n7948 0.823357
R47475 VCC.n7996 VCC.n7941 0.823357
R47476 VCC.n8013 VCC.n7919 0.823357
R47477 VCC.n8049 VCC.n7908 0.823357
R47478 VCC.n8656 VCC.n8655 0.823357
R47479 VCC.n8672 VCC.n8425 0.823357
R47480 VCC.n8702 VCC.n8701 0.823357
R47481 VCC.n8727 VCC.n8399 0.823357
R47482 VCC.n8538 VCC.n8499 0.823357
R47483 VCC.n8547 VCC.n8492 0.823357
R47484 VCC.n8564 VCC.n8470 0.823357
R47485 VCC.n8600 VCC.n8459 0.823357
R47486 VCC.n9213 VCC.n9212 0.823357
R47487 VCC.n9229 VCC.n8982 0.823357
R47488 VCC.n9259 VCC.n9258 0.823357
R47489 VCC.n9284 VCC.n8956 0.823357
R47490 VCC.n9096 VCC.n9057 0.823357
R47491 VCC.n9105 VCC.n9050 0.823357
R47492 VCC.n9122 VCC.n9028 0.823357
R47493 VCC.n9158 VCC.n9017 0.823357
R47494 VCC.n9647 VCC.n9608 0.823357
R47495 VCC.n9656 VCC.n9601 0.823357
R47496 VCC.n9673 VCC.n9579 0.823357
R47497 VCC.n9709 VCC.n9568 0.823357
R47498 VCC.n9765 VCC.n9764 0.823357
R47499 VCC.n9781 VCC.n9534 0.823357
R47500 VCC.n9811 VCC.n9810 0.823357
R47501 VCC.n9836 VCC.n9508 0.823357
R47502 VCC.n10321 VCC.n10320 0.823357
R47503 VCC.n10337 VCC.n10090 0.823357
R47504 VCC.n10367 VCC.n10366 0.823357
R47505 VCC.n10392 VCC.n10064 0.823357
R47506 VCC.n10204 VCC.n10165 0.823357
R47507 VCC.n10213 VCC.n10158 0.823357
R47508 VCC.n10230 VCC.n10136 0.823357
R47509 VCC.n10266 VCC.n10125 0.823357
R47510 VCC.n10754 VCC.n10715 0.823357
R47511 VCC.n10763 VCC.n10708 0.823357
R47512 VCC.n10780 VCC.n10686 0.823357
R47513 VCC.n10816 VCC.n10675 0.823357
R47514 VCC.n10872 VCC.n10871 0.823357
R47515 VCC.n10888 VCC.n10641 0.823357
R47516 VCC.n10918 VCC.n10917 0.823357
R47517 VCC.n10943 VCC.n10615 0.823357
R47518 VCC.n11428 VCC.n11427 0.823357
R47519 VCC.n11444 VCC.n11197 0.823357
R47520 VCC.n11474 VCC.n11473 0.823357
R47521 VCC.n11499 VCC.n11171 0.823357
R47522 VCC.n11311 VCC.n11272 0.823357
R47523 VCC.n11320 VCC.n11265 0.823357
R47524 VCC.n11337 VCC.n11243 0.823357
R47525 VCC.n11373 VCC.n11232 0.823357
R47526 VCC.n11861 VCC.n11822 0.823357
R47527 VCC.n11870 VCC.n11815 0.823357
R47528 VCC.n11887 VCC.n11793 0.823357
R47529 VCC.n11923 VCC.n11782 0.823357
R47530 VCC.n11979 VCC.n11978 0.823357
R47531 VCC.n11995 VCC.n11748 0.823357
R47532 VCC.n12025 VCC.n12024 0.823357
R47533 VCC.n12050 VCC.n11722 0.823357
R47534 VCC.n12535 VCC.n12534 0.823357
R47535 VCC.n12551 VCC.n12304 0.823357
R47536 VCC.n12581 VCC.n12580 0.823357
R47537 VCC.n12606 VCC.n12278 0.823357
R47538 VCC.n12418 VCC.n12379 0.823357
R47539 VCC.n12427 VCC.n12372 0.823357
R47540 VCC.n12444 VCC.n12350 0.823357
R47541 VCC.n12480 VCC.n12339 0.823357
R47542 VCC.n12968 VCC.n12929 0.823357
R47543 VCC.n12977 VCC.n12922 0.823357
R47544 VCC.n12994 VCC.n12900 0.823357
R47545 VCC.n13030 VCC.n12889 0.823357
R47546 VCC.n13086 VCC.n13085 0.823357
R47547 VCC.n13102 VCC.n12855 0.823357
R47548 VCC.n13132 VCC.n13131 0.823357
R47549 VCC.n13157 VCC.n12829 0.823357
R47550 VCC.n13642 VCC.n13641 0.823357
R47551 VCC.n13658 VCC.n13411 0.823357
R47552 VCC.n13688 VCC.n13687 0.823357
R47553 VCC.n13713 VCC.n13385 0.823357
R47554 VCC.n13525 VCC.n13486 0.823357
R47555 VCC.n13534 VCC.n13479 0.823357
R47556 VCC.n13551 VCC.n13457 0.823357
R47557 VCC.n13587 VCC.n13446 0.823357
R47558 VCC.n14075 VCC.n14036 0.823357
R47559 VCC.n14084 VCC.n14029 0.823357
R47560 VCC.n14101 VCC.n14007 0.823357
R47561 VCC.n14137 VCC.n13996 0.823357
R47562 VCC.n14193 VCC.n14192 0.823357
R47563 VCC.n14209 VCC.n13962 0.823357
R47564 VCC.n14239 VCC.n14238 0.823357
R47565 VCC.n14264 VCC.n13936 0.823357
R47566 VCC.n14749 VCC.n14748 0.823357
R47567 VCC.n14765 VCC.n14518 0.823357
R47568 VCC.n14795 VCC.n14794 0.823357
R47569 VCC.n14820 VCC.n14492 0.823357
R47570 VCC.n14632 VCC.n14593 0.823357
R47571 VCC.n14641 VCC.n14586 0.823357
R47572 VCC.n14658 VCC.n14564 0.823357
R47573 VCC.n14694 VCC.n14553 0.823357
R47574 VCC.n15182 VCC.n15143 0.823357
R47575 VCC.n15191 VCC.n15136 0.823357
R47576 VCC.n15208 VCC.n15114 0.823357
R47577 VCC.n15244 VCC.n15103 0.823357
R47578 VCC.n15300 VCC.n15299 0.823357
R47579 VCC.n15316 VCC.n15069 0.823357
R47580 VCC.n15346 VCC.n15345 0.823357
R47581 VCC.n15371 VCC.n15043 0.823357
R47582 VCC.n15856 VCC.n15855 0.823357
R47583 VCC.n15872 VCC.n15625 0.823357
R47584 VCC.n15902 VCC.n15901 0.823357
R47585 VCC.n15927 VCC.n15599 0.823357
R47586 VCC.n15739 VCC.n15700 0.823357
R47587 VCC.n15748 VCC.n15693 0.823357
R47588 VCC.n15765 VCC.n15671 0.823357
R47589 VCC.n15801 VCC.n15660 0.823357
R47590 VCC.n16289 VCC.n16250 0.823357
R47591 VCC.n16298 VCC.n16243 0.823357
R47592 VCC.n16315 VCC.n16221 0.823357
R47593 VCC.n16351 VCC.n16210 0.823357
R47594 VCC.n16407 VCC.n16406 0.823357
R47595 VCC.n16423 VCC.n16176 0.823357
R47596 VCC.n16453 VCC.n16452 0.823357
R47597 VCC.n16478 VCC.n16150 0.823357
R47598 VCC.n16963 VCC.n16962 0.823357
R47599 VCC.n16979 VCC.n16732 0.823357
R47600 VCC.n17009 VCC.n17008 0.823357
R47601 VCC.n17034 VCC.n16706 0.823357
R47602 VCC.n16846 VCC.n16807 0.823357
R47603 VCC.n16855 VCC.n16800 0.823357
R47604 VCC.n16872 VCC.n16778 0.823357
R47605 VCC.n16908 VCC.n16767 0.823357
R47606 VCC.n17327 VCC.n17326 0.823357
R47607 VCC.n17343 VCC.n17283 0.823357
R47608 VCC.n17373 VCC.n17372 0.823357
R47609 VCC.n17398 VCC.n17257 0.823357
R47610 VCC.n184 VCC.n177 0.731929
R47611 VCC.n272 VCC.n144 0.731929
R47612 VCC.n287 VCC.n285 0.731929
R47613 VCC.n340 VCC.n110 0.731929
R47614 VCC.n399 VCC.n84 0.731929
R47615 VCC.n413 VCC.n412 0.731929
R47616 VCC.n736 VCC.n729 0.731929
R47617 VCC.n824 VCC.n696 0.731929
R47618 VCC.n839 VCC.n837 0.731929
R47619 VCC.n892 VCC.n662 0.731929
R47620 VCC.n951 VCC.n636 0.731929
R47621 VCC.n965 VCC.n964 0.731929
R47622 VCC.n1449 VCC.n1219 0.731929
R47623 VCC.n1508 VCC.n1193 0.731929
R47624 VCC.n1522 VCC.n1521 0.731929
R47625 VCC.n1294 VCC.n1287 0.731929
R47626 VCC.n1382 VCC.n1254 0.731929
R47627 VCC.n1397 VCC.n1395 0.731929
R47628 VCC.n1845 VCC.n1838 0.731929
R47629 VCC.n1933 VCC.n1805 0.731929
R47630 VCC.n1948 VCC.n1946 0.731929
R47631 VCC.n2001 VCC.n1771 0.731929
R47632 VCC.n2060 VCC.n1745 0.731929
R47633 VCC.n2074 VCC.n2073 0.731929
R47634 VCC.n2558 VCC.n2328 0.731929
R47635 VCC.n2617 VCC.n2302 0.731929
R47636 VCC.n2631 VCC.n2630 0.731929
R47637 VCC.n2403 VCC.n2396 0.731929
R47638 VCC.n2491 VCC.n2363 0.731929
R47639 VCC.n2506 VCC.n2504 0.731929
R47640 VCC.n2954 VCC.n2947 0.731929
R47641 VCC.n3042 VCC.n2914 0.731929
R47642 VCC.n3057 VCC.n3055 0.731929
R47643 VCC.n3110 VCC.n2880 0.731929
R47644 VCC.n3169 VCC.n2854 0.731929
R47645 VCC.n3183 VCC.n3182 0.731929
R47646 VCC.n3667 VCC.n3437 0.731929
R47647 VCC.n3726 VCC.n3411 0.731929
R47648 VCC.n3740 VCC.n3739 0.731929
R47649 VCC.n3512 VCC.n3505 0.731929
R47650 VCC.n3600 VCC.n3472 0.731929
R47651 VCC.n3615 VCC.n3613 0.731929
R47652 VCC.n4063 VCC.n4056 0.731929
R47653 VCC.n4151 VCC.n4023 0.731929
R47654 VCC.n4166 VCC.n4164 0.731929
R47655 VCC.n4219 VCC.n3989 0.731929
R47656 VCC.n4278 VCC.n3963 0.731929
R47657 VCC.n4292 VCC.n4291 0.731929
R47658 VCC.n4776 VCC.n4546 0.731929
R47659 VCC.n4835 VCC.n4520 0.731929
R47660 VCC.n4849 VCC.n4848 0.731929
R47661 VCC.n4621 VCC.n4614 0.731929
R47662 VCC.n4709 VCC.n4581 0.731929
R47663 VCC.n4724 VCC.n4722 0.731929
R47664 VCC.n5172 VCC.n5165 0.731929
R47665 VCC.n5260 VCC.n5132 0.731929
R47666 VCC.n5275 VCC.n5273 0.731929
R47667 VCC.n5328 VCC.n5098 0.731929
R47668 VCC.n5387 VCC.n5072 0.731929
R47669 VCC.n5401 VCC.n5400 0.731929
R47670 VCC.n5885 VCC.n5655 0.731929
R47671 VCC.n5944 VCC.n5629 0.731929
R47672 VCC.n5958 VCC.n5957 0.731929
R47673 VCC.n5730 VCC.n5723 0.731929
R47674 VCC.n5818 VCC.n5690 0.731929
R47675 VCC.n5833 VCC.n5831 0.731929
R47676 VCC.n6281 VCC.n6274 0.731929
R47677 VCC.n6369 VCC.n6241 0.731929
R47678 VCC.n6384 VCC.n6382 0.731929
R47679 VCC.n6437 VCC.n6207 0.731929
R47680 VCC.n6496 VCC.n6181 0.731929
R47681 VCC.n6510 VCC.n6509 0.731929
R47682 VCC.n6994 VCC.n6764 0.731929
R47683 VCC.n7053 VCC.n6738 0.731929
R47684 VCC.n7067 VCC.n7066 0.731929
R47685 VCC.n6839 VCC.n6832 0.731929
R47686 VCC.n6927 VCC.n6799 0.731929
R47687 VCC.n6942 VCC.n6940 0.731929
R47688 VCC.n7390 VCC.n7383 0.731929
R47689 VCC.n7478 VCC.n7350 0.731929
R47690 VCC.n7493 VCC.n7491 0.731929
R47691 VCC.n7546 VCC.n7316 0.731929
R47692 VCC.n7605 VCC.n7290 0.731929
R47693 VCC.n7619 VCC.n7618 0.731929
R47694 VCC.n8103 VCC.n7873 0.731929
R47695 VCC.n8162 VCC.n7847 0.731929
R47696 VCC.n8176 VCC.n8175 0.731929
R47697 VCC.n7948 VCC.n7941 0.731929
R47698 VCC.n8036 VCC.n7908 0.731929
R47699 VCC.n8051 VCC.n8049 0.731929
R47700 VCC.n8655 VCC.n8425 0.731929
R47701 VCC.n8714 VCC.n8399 0.731929
R47702 VCC.n8728 VCC.n8727 0.731929
R47703 VCC.n8499 VCC.n8492 0.731929
R47704 VCC.n8587 VCC.n8459 0.731929
R47705 VCC.n8602 VCC.n8600 0.731929
R47706 VCC.n9212 VCC.n8982 0.731929
R47707 VCC.n9271 VCC.n8956 0.731929
R47708 VCC.n9285 VCC.n9284 0.731929
R47709 VCC.n9057 VCC.n9050 0.731929
R47710 VCC.n9145 VCC.n9017 0.731929
R47711 VCC.n9160 VCC.n9158 0.731929
R47712 VCC.n9608 VCC.n9601 0.731929
R47713 VCC.n9696 VCC.n9568 0.731929
R47714 VCC.n9711 VCC.n9709 0.731929
R47715 VCC.n9764 VCC.n9534 0.731929
R47716 VCC.n9823 VCC.n9508 0.731929
R47717 VCC.n9837 VCC.n9836 0.731929
R47718 VCC.n10320 VCC.n10090 0.731929
R47719 VCC.n10379 VCC.n10064 0.731929
R47720 VCC.n10393 VCC.n10392 0.731929
R47721 VCC.n10165 VCC.n10158 0.731929
R47722 VCC.n10253 VCC.n10125 0.731929
R47723 VCC.n10268 VCC.n10266 0.731929
R47724 VCC.n10715 VCC.n10708 0.731929
R47725 VCC.n10803 VCC.n10675 0.731929
R47726 VCC.n10818 VCC.n10816 0.731929
R47727 VCC.n10871 VCC.n10641 0.731929
R47728 VCC.n10930 VCC.n10615 0.731929
R47729 VCC.n10944 VCC.n10943 0.731929
R47730 VCC.n11427 VCC.n11197 0.731929
R47731 VCC.n11486 VCC.n11171 0.731929
R47732 VCC.n11500 VCC.n11499 0.731929
R47733 VCC.n11272 VCC.n11265 0.731929
R47734 VCC.n11360 VCC.n11232 0.731929
R47735 VCC.n11375 VCC.n11373 0.731929
R47736 VCC.n11822 VCC.n11815 0.731929
R47737 VCC.n11910 VCC.n11782 0.731929
R47738 VCC.n11925 VCC.n11923 0.731929
R47739 VCC.n11978 VCC.n11748 0.731929
R47740 VCC.n12037 VCC.n11722 0.731929
R47741 VCC.n12051 VCC.n12050 0.731929
R47742 VCC.n12534 VCC.n12304 0.731929
R47743 VCC.n12593 VCC.n12278 0.731929
R47744 VCC.n12607 VCC.n12606 0.731929
R47745 VCC.n12379 VCC.n12372 0.731929
R47746 VCC.n12467 VCC.n12339 0.731929
R47747 VCC.n12482 VCC.n12480 0.731929
R47748 VCC.n12929 VCC.n12922 0.731929
R47749 VCC.n13017 VCC.n12889 0.731929
R47750 VCC.n13032 VCC.n13030 0.731929
R47751 VCC.n13085 VCC.n12855 0.731929
R47752 VCC.n13144 VCC.n12829 0.731929
R47753 VCC.n13158 VCC.n13157 0.731929
R47754 VCC.n13641 VCC.n13411 0.731929
R47755 VCC.n13700 VCC.n13385 0.731929
R47756 VCC.n13714 VCC.n13713 0.731929
R47757 VCC.n13486 VCC.n13479 0.731929
R47758 VCC.n13574 VCC.n13446 0.731929
R47759 VCC.n13589 VCC.n13587 0.731929
R47760 VCC.n14036 VCC.n14029 0.731929
R47761 VCC.n14124 VCC.n13996 0.731929
R47762 VCC.n14139 VCC.n14137 0.731929
R47763 VCC.n14192 VCC.n13962 0.731929
R47764 VCC.n14251 VCC.n13936 0.731929
R47765 VCC.n14265 VCC.n14264 0.731929
R47766 VCC.n14748 VCC.n14518 0.731929
R47767 VCC.n14807 VCC.n14492 0.731929
R47768 VCC.n14821 VCC.n14820 0.731929
R47769 VCC.n14593 VCC.n14586 0.731929
R47770 VCC.n14681 VCC.n14553 0.731929
R47771 VCC.n14696 VCC.n14694 0.731929
R47772 VCC.n15143 VCC.n15136 0.731929
R47773 VCC.n15231 VCC.n15103 0.731929
R47774 VCC.n15246 VCC.n15244 0.731929
R47775 VCC.n15299 VCC.n15069 0.731929
R47776 VCC.n15358 VCC.n15043 0.731929
R47777 VCC.n15372 VCC.n15371 0.731929
R47778 VCC.n15855 VCC.n15625 0.731929
R47779 VCC.n15914 VCC.n15599 0.731929
R47780 VCC.n15928 VCC.n15927 0.731929
R47781 VCC.n15700 VCC.n15693 0.731929
R47782 VCC.n15788 VCC.n15660 0.731929
R47783 VCC.n15803 VCC.n15801 0.731929
R47784 VCC.n16250 VCC.n16243 0.731929
R47785 VCC.n16338 VCC.n16210 0.731929
R47786 VCC.n16353 VCC.n16351 0.731929
R47787 VCC.n16406 VCC.n16176 0.731929
R47788 VCC.n16465 VCC.n16150 0.731929
R47789 VCC.n16479 VCC.n16478 0.731929
R47790 VCC.n16962 VCC.n16732 0.731929
R47791 VCC.n17021 VCC.n16706 0.731929
R47792 VCC.n17035 VCC.n17034 0.731929
R47793 VCC.n16807 VCC.n16800 0.731929
R47794 VCC.n16895 VCC.n16767 0.731929
R47795 VCC.n16910 VCC.n16908 0.731929
R47796 VCC.n17326 VCC.n17283 0.731929
R47797 VCC.n17385 VCC.n17257 0.731929
R47798 VCC.n17399 VCC.n17398 0.731929
R47799 VCC.n247 VCC.n169 0.6405
R47800 VCC.n297 VCC.n296 0.6405
R47801 VCC.n366 VCC.n364 0.6405
R47802 VCC.n432 VCC.n431 0.6405
R47803 VCC.n799 VCC.n721 0.6405
R47804 VCC.n849 VCC.n848 0.6405
R47805 VCC.n918 VCC.n916 0.6405
R47806 VCC.n984 VCC.n983 0.6405
R47807 VCC.n1475 VCC.n1473 0.6405
R47808 VCC.n1542 VCC.n1541 0.6405
R47809 VCC.n1357 VCC.n1279 0.6405
R47810 VCC.n1407 VCC.n1406 0.6405
R47811 VCC.n1908 VCC.n1830 0.6405
R47812 VCC.n1958 VCC.n1957 0.6405
R47813 VCC.n2027 VCC.n2025 0.6405
R47814 VCC.n2093 VCC.n2092 0.6405
R47815 VCC.n2584 VCC.n2582 0.6405
R47816 VCC.n2651 VCC.n2650 0.6405
R47817 VCC.n2466 VCC.n2388 0.6405
R47818 VCC.n2516 VCC.n2515 0.6405
R47819 VCC.n3017 VCC.n2939 0.6405
R47820 VCC.n3067 VCC.n3066 0.6405
R47821 VCC.n3136 VCC.n3134 0.6405
R47822 VCC.n3202 VCC.n3201 0.6405
R47823 VCC.n3693 VCC.n3691 0.6405
R47824 VCC.n3760 VCC.n3759 0.6405
R47825 VCC.n3575 VCC.n3497 0.6405
R47826 VCC.n3625 VCC.n3624 0.6405
R47827 VCC.n4126 VCC.n4048 0.6405
R47828 VCC.n4176 VCC.n4175 0.6405
R47829 VCC.n4245 VCC.n4243 0.6405
R47830 VCC.n4311 VCC.n4310 0.6405
R47831 VCC.n4802 VCC.n4800 0.6405
R47832 VCC.n4869 VCC.n4868 0.6405
R47833 VCC.n4684 VCC.n4606 0.6405
R47834 VCC.n4734 VCC.n4733 0.6405
R47835 VCC.n5235 VCC.n5157 0.6405
R47836 VCC.n5285 VCC.n5284 0.6405
R47837 VCC.n5354 VCC.n5352 0.6405
R47838 VCC.n5420 VCC.n5419 0.6405
R47839 VCC.n5911 VCC.n5909 0.6405
R47840 VCC.n5978 VCC.n5977 0.6405
R47841 VCC.n5793 VCC.n5715 0.6405
R47842 VCC.n5843 VCC.n5842 0.6405
R47843 VCC.n6344 VCC.n6266 0.6405
R47844 VCC.n6394 VCC.n6393 0.6405
R47845 VCC.n6463 VCC.n6461 0.6405
R47846 VCC.n6529 VCC.n6528 0.6405
R47847 VCC.n7020 VCC.n7018 0.6405
R47848 VCC.n7087 VCC.n7086 0.6405
R47849 VCC.n6902 VCC.n6824 0.6405
R47850 VCC.n6952 VCC.n6951 0.6405
R47851 VCC.n7453 VCC.n7375 0.6405
R47852 VCC.n7503 VCC.n7502 0.6405
R47853 VCC.n7572 VCC.n7570 0.6405
R47854 VCC.n7638 VCC.n7637 0.6405
R47855 VCC.n8129 VCC.n8127 0.6405
R47856 VCC.n8196 VCC.n8195 0.6405
R47857 VCC.n8011 VCC.n7933 0.6405
R47858 VCC.n8061 VCC.n8060 0.6405
R47859 VCC.n8681 VCC.n8679 0.6405
R47860 VCC.n8747 VCC.n8746 0.6405
R47861 VCC.n8562 VCC.n8484 0.6405
R47862 VCC.n8612 VCC.n8611 0.6405
R47863 VCC.n9238 VCC.n9236 0.6405
R47864 VCC.n9305 VCC.n9304 0.6405
R47865 VCC.n9120 VCC.n9042 0.6405
R47866 VCC.n9170 VCC.n9169 0.6405
R47867 VCC.n9671 VCC.n9593 0.6405
R47868 VCC.n9721 VCC.n9720 0.6405
R47869 VCC.n9790 VCC.n9788 0.6405
R47870 VCC.n9856 VCC.n9855 0.6405
R47871 VCC.n10346 VCC.n10344 0.6405
R47872 VCC.n10413 VCC.n10412 0.6405
R47873 VCC.n10228 VCC.n10150 0.6405
R47874 VCC.n10278 VCC.n10277 0.6405
R47875 VCC.n10778 VCC.n10700 0.6405
R47876 VCC.n10828 VCC.n10827 0.6405
R47877 VCC.n10897 VCC.n10895 0.6405
R47878 VCC.n10963 VCC.n10962 0.6405
R47879 VCC.n11453 VCC.n11451 0.6405
R47880 VCC.n11520 VCC.n11519 0.6405
R47881 VCC.n11335 VCC.n11257 0.6405
R47882 VCC.n11385 VCC.n11384 0.6405
R47883 VCC.n11885 VCC.n11807 0.6405
R47884 VCC.n11935 VCC.n11934 0.6405
R47885 VCC.n12004 VCC.n12002 0.6405
R47886 VCC.n12070 VCC.n12069 0.6405
R47887 VCC.n12560 VCC.n12558 0.6405
R47888 VCC.n12627 VCC.n12626 0.6405
R47889 VCC.n12442 VCC.n12364 0.6405
R47890 VCC.n12492 VCC.n12491 0.6405
R47891 VCC.n12992 VCC.n12914 0.6405
R47892 VCC.n13042 VCC.n13041 0.6405
R47893 VCC.n13111 VCC.n13109 0.6405
R47894 VCC.n13177 VCC.n13176 0.6405
R47895 VCC.n13667 VCC.n13665 0.6405
R47896 VCC.n13734 VCC.n13733 0.6405
R47897 VCC.n13549 VCC.n13471 0.6405
R47898 VCC.n13599 VCC.n13598 0.6405
R47899 VCC.n14099 VCC.n14021 0.6405
R47900 VCC.n14149 VCC.n14148 0.6405
R47901 VCC.n14218 VCC.n14216 0.6405
R47902 VCC.n14284 VCC.n14283 0.6405
R47903 VCC.n14774 VCC.n14772 0.6405
R47904 VCC.n14841 VCC.n14840 0.6405
R47905 VCC.n14656 VCC.n14578 0.6405
R47906 VCC.n14706 VCC.n14705 0.6405
R47907 VCC.n15206 VCC.n15128 0.6405
R47908 VCC.n15256 VCC.n15255 0.6405
R47909 VCC.n15325 VCC.n15323 0.6405
R47910 VCC.n15391 VCC.n15390 0.6405
R47911 VCC.n15881 VCC.n15879 0.6405
R47912 VCC.n15948 VCC.n15947 0.6405
R47913 VCC.n15763 VCC.n15685 0.6405
R47914 VCC.n15813 VCC.n15812 0.6405
R47915 VCC.n16313 VCC.n16235 0.6405
R47916 VCC.n16363 VCC.n16362 0.6405
R47917 VCC.n16432 VCC.n16430 0.6405
R47918 VCC.n16498 VCC.n16497 0.6405
R47919 VCC.n16988 VCC.n16986 0.6405
R47920 VCC.n17055 VCC.n17054 0.6405
R47921 VCC.n16870 VCC.n16792 0.6405
R47922 VCC.n16920 VCC.n16919 0.6405
R47923 VCC.n17352 VCC.n17350 0.6405
R47924 VCC.n17418 VCC.n17417 0.6405
R47925 VCC.n4989 VCC 0.621824
R47926 VCC VCC.n17547 0.621824
R47927 VCC.n207 VCC.n195 0.549071
R47928 VCC.n159 VCC.n151 0.549071
R47929 VCC.n325 VCC.n124 0.549071
R47930 VCC.n392 VCC.n391 0.549071
R47931 VCC.n759 VCC.n747 0.549071
R47932 VCC.n711 VCC.n703 0.549071
R47933 VCC.n877 VCC.n676 0.549071
R47934 VCC.n944 VCC.n943 0.549071
R47935 VCC.n1434 VCC.n1233 0.549071
R47936 VCC.n1501 VCC.n1500 0.549071
R47937 VCC.n1317 VCC.n1305 0.549071
R47938 VCC.n1269 VCC.n1261 0.549071
R47939 VCC.n1868 VCC.n1856 0.549071
R47940 VCC.n1820 VCC.n1812 0.549071
R47941 VCC.n1986 VCC.n1785 0.549071
R47942 VCC.n2053 VCC.n2052 0.549071
R47943 VCC.n2543 VCC.n2342 0.549071
R47944 VCC.n2610 VCC.n2609 0.549071
R47945 VCC.n2426 VCC.n2414 0.549071
R47946 VCC.n2378 VCC.n2370 0.549071
R47947 VCC.n2977 VCC.n2965 0.549071
R47948 VCC.n2929 VCC.n2921 0.549071
R47949 VCC.n3095 VCC.n2894 0.549071
R47950 VCC.n3162 VCC.n3161 0.549071
R47951 VCC.n3652 VCC.n3451 0.549071
R47952 VCC.n3719 VCC.n3718 0.549071
R47953 VCC.n3535 VCC.n3523 0.549071
R47954 VCC.n3487 VCC.n3479 0.549071
R47955 VCC.n4086 VCC.n4074 0.549071
R47956 VCC.n4038 VCC.n4030 0.549071
R47957 VCC.n4204 VCC.n4003 0.549071
R47958 VCC.n4271 VCC.n4270 0.549071
R47959 VCC.n4761 VCC.n4560 0.549071
R47960 VCC.n4828 VCC.n4827 0.549071
R47961 VCC.n4644 VCC.n4632 0.549071
R47962 VCC.n4596 VCC.n4588 0.549071
R47963 VCC.n5195 VCC.n5183 0.549071
R47964 VCC.n5147 VCC.n5139 0.549071
R47965 VCC.n5313 VCC.n5112 0.549071
R47966 VCC.n5380 VCC.n5379 0.549071
R47967 VCC.n5870 VCC.n5669 0.549071
R47968 VCC.n5937 VCC.n5936 0.549071
R47969 VCC.n5753 VCC.n5741 0.549071
R47970 VCC.n5705 VCC.n5697 0.549071
R47971 VCC.n6304 VCC.n6292 0.549071
R47972 VCC.n6256 VCC.n6248 0.549071
R47973 VCC.n6422 VCC.n6221 0.549071
R47974 VCC.n6489 VCC.n6488 0.549071
R47975 VCC.n6979 VCC.n6778 0.549071
R47976 VCC.n7046 VCC.n7045 0.549071
R47977 VCC.n6862 VCC.n6850 0.549071
R47978 VCC.n6814 VCC.n6806 0.549071
R47979 VCC.n7413 VCC.n7401 0.549071
R47980 VCC.n7365 VCC.n7357 0.549071
R47981 VCC.n7531 VCC.n7330 0.549071
R47982 VCC.n7598 VCC.n7597 0.549071
R47983 VCC.n8088 VCC.n7887 0.549071
R47984 VCC.n8155 VCC.n8154 0.549071
R47985 VCC.n7971 VCC.n7959 0.549071
R47986 VCC.n7923 VCC.n7915 0.549071
R47987 VCC.n8640 VCC.n8439 0.549071
R47988 VCC.n8707 VCC.n8706 0.549071
R47989 VCC.n8522 VCC.n8510 0.549071
R47990 VCC.n8474 VCC.n8466 0.549071
R47991 VCC.n9197 VCC.n8996 0.549071
R47992 VCC.n9264 VCC.n9263 0.549071
R47993 VCC.n9080 VCC.n9068 0.549071
R47994 VCC.n9032 VCC.n9024 0.549071
R47995 VCC.n9631 VCC.n9619 0.549071
R47996 VCC.n9583 VCC.n9575 0.549071
R47997 VCC.n9749 VCC.n9548 0.549071
R47998 VCC.n9816 VCC.n9815 0.549071
R47999 VCC.n10305 VCC.n10104 0.549071
R48000 VCC.n10372 VCC.n10371 0.549071
R48001 VCC.n10188 VCC.n10176 0.549071
R48002 VCC.n10140 VCC.n10132 0.549071
R48003 VCC.n10738 VCC.n10726 0.549071
R48004 VCC.n10690 VCC.n10682 0.549071
R48005 VCC.n10856 VCC.n10655 0.549071
R48006 VCC.n10923 VCC.n10922 0.549071
R48007 VCC.n11412 VCC.n11211 0.549071
R48008 VCC.n11479 VCC.n11478 0.549071
R48009 VCC.n11295 VCC.n11283 0.549071
R48010 VCC.n11247 VCC.n11239 0.549071
R48011 VCC.n11845 VCC.n11833 0.549071
R48012 VCC.n11797 VCC.n11789 0.549071
R48013 VCC.n11963 VCC.n11762 0.549071
R48014 VCC.n12030 VCC.n12029 0.549071
R48015 VCC.n12519 VCC.n12318 0.549071
R48016 VCC.n12586 VCC.n12585 0.549071
R48017 VCC.n12402 VCC.n12390 0.549071
R48018 VCC.n12354 VCC.n12346 0.549071
R48019 VCC.n12952 VCC.n12940 0.549071
R48020 VCC.n12904 VCC.n12896 0.549071
R48021 VCC.n13070 VCC.n12869 0.549071
R48022 VCC.n13137 VCC.n13136 0.549071
R48023 VCC.n13626 VCC.n13425 0.549071
R48024 VCC.n13693 VCC.n13692 0.549071
R48025 VCC.n13509 VCC.n13497 0.549071
R48026 VCC.n13461 VCC.n13453 0.549071
R48027 VCC.n14059 VCC.n14047 0.549071
R48028 VCC.n14011 VCC.n14003 0.549071
R48029 VCC.n14177 VCC.n13976 0.549071
R48030 VCC.n14244 VCC.n14243 0.549071
R48031 VCC.n14733 VCC.n14532 0.549071
R48032 VCC.n14800 VCC.n14799 0.549071
R48033 VCC.n14616 VCC.n14604 0.549071
R48034 VCC.n14568 VCC.n14560 0.549071
R48035 VCC.n15166 VCC.n15154 0.549071
R48036 VCC.n15118 VCC.n15110 0.549071
R48037 VCC.n15284 VCC.n15083 0.549071
R48038 VCC.n15351 VCC.n15350 0.549071
R48039 VCC.n15840 VCC.n15639 0.549071
R48040 VCC.n15907 VCC.n15906 0.549071
R48041 VCC.n15723 VCC.n15711 0.549071
R48042 VCC.n15675 VCC.n15667 0.549071
R48043 VCC.n16273 VCC.n16261 0.549071
R48044 VCC.n16225 VCC.n16217 0.549071
R48045 VCC.n16391 VCC.n16190 0.549071
R48046 VCC.n16458 VCC.n16457 0.549071
R48047 VCC.n16947 VCC.n16746 0.549071
R48048 VCC.n17014 VCC.n17013 0.549071
R48049 VCC.n16830 VCC.n16818 0.549071
R48050 VCC.n16782 VCC.n16774 0.549071
R48051 VCC.n17311 VCC.n17297 0.549071
R48052 VCC.n17378 VCC.n17377 0.549071
R48053 VCC.n449 VCC 0.535293
R48054 VCC.n1001 VCC 0.535293
R48055 VCC.n1559 VCC 0.535293
R48056 VCC.n2110 VCC 0.535293
R48057 VCC.n2668 VCC 0.535293
R48058 VCC.n3219 VCC 0.535293
R48059 VCC.n3777 VCC 0.535293
R48060 VCC.n4328 VCC 0.535293
R48061 VCC.n4886 VCC 0.535293
R48062 VCC.n5437 VCC 0.535293
R48063 VCC.n5995 VCC 0.535293
R48064 VCC.n6546 VCC 0.535293
R48065 VCC.n7104 VCC 0.535293
R48066 VCC.n7655 VCC 0.535293
R48067 VCC.n8213 VCC 0.535293
R48068 VCC.n8764 VCC 0.535293
R48069 VCC.n9322 VCC 0.535293
R48070 VCC.n9873 VCC 0.535293
R48071 VCC.n10430 VCC 0.535293
R48072 VCC.n10980 VCC 0.535293
R48073 VCC.n11537 VCC 0.535293
R48074 VCC.n12087 VCC 0.535293
R48075 VCC.n12644 VCC 0.535293
R48076 VCC.n13194 VCC 0.535293
R48077 VCC.n13751 VCC 0.535293
R48078 VCC.n14301 VCC 0.535293
R48079 VCC.n14858 VCC 0.535293
R48080 VCC.n15408 VCC 0.535293
R48081 VCC.n15965 VCC 0.535293
R48082 VCC.n16515 VCC 0.535293
R48083 VCC.n17072 VCC 0.535293
R48084 VCC.n17435 VCC 0.535293
R48085 VCC.n549 VCC.n3 0.507747
R48086 VCC.n1103 VCC.n557 0.507747
R48087 VCC.n1657 VCC.n1656 0.507747
R48088 VCC.n2212 VCC.n1666 0.507747
R48089 VCC.n2766 VCC.n2765 0.507747
R48090 VCC.n3321 VCC.n2775 0.507747
R48091 VCC.n3875 VCC.n3874 0.507747
R48092 VCC.n4430 VCC.n3884 0.507747
R48093 VCC.n4984 VCC.n4983 0.507747
R48094 VCC.n5539 VCC.n4993 0.507747
R48095 VCC.n6093 VCC.n6092 0.507747
R48096 VCC.n6648 VCC.n6102 0.507747
R48097 VCC.n7202 VCC.n7201 0.507747
R48098 VCC.n7757 VCC.n7211 0.507747
R48099 VCC.n8311 VCC.n8310 0.507747
R48100 VCC.n8866 VCC.n8320 0.507747
R48101 VCC.n9420 VCC.n9419 0.507747
R48102 VCC.n9975 VCC.n9429 0.507747
R48103 VCC.n10528 VCC.n10527 0.507747
R48104 VCC.n11082 VCC.n10536 0.507747
R48105 VCC.n11635 VCC.n11634 0.507747
R48106 VCC.n12189 VCC.n11643 0.507747
R48107 VCC.n12742 VCC.n12741 0.507747
R48108 VCC.n13296 VCC.n12750 0.507747
R48109 VCC.n13849 VCC.n13848 0.507747
R48110 VCC.n14403 VCC.n13857 0.507747
R48111 VCC.n14956 VCC.n14955 0.507747
R48112 VCC.n15510 VCC.n14964 0.507747
R48113 VCC.n16063 VCC.n16062 0.507747
R48114 VCC.n16617 VCC.n16071 0.507747
R48115 VCC.n17170 VCC.n17169 0.507747
R48116 VCC.n17537 VCC.n17178 0.507747
R48117 VCC.n9425 VCC 0.474765
R48118 VCC.n1532 VCC.n1174 0.465127
R48119 VCC.n2641 VCC.n2283 0.465127
R48120 VCC.n3750 VCC.n3392 0.465127
R48121 VCC.n4859 VCC.n4501 0.465127
R48122 VCC.n5968 VCC.n5610 0.465127
R48123 VCC.n7077 VCC.n6719 0.465127
R48124 VCC.n8186 VCC.n7828 0.465127
R48125 VCC.n9295 VCC.n8937 0.465127
R48126 VCC.n10403 VCC.n10045 0.465127
R48127 VCC.n11510 VCC.n11152 0.465127
R48128 VCC.n12617 VCC.n12259 0.465127
R48129 VCC.n13724 VCC.n13366 0.465127
R48130 VCC.n14831 VCC.n14473 0.465127
R48131 VCC.n15938 VCC.n15580 0.465127
R48132 VCC.n17045 VCC.n16687 0.465127
R48133 VCC.n422 VCC.n65 0.465115
R48134 VCC.n974 VCC.n617 0.465115
R48135 VCC.n2083 VCC.n1726 0.465115
R48136 VCC.n3192 VCC.n2835 0.465115
R48137 VCC.n4301 VCC.n3944 0.465115
R48138 VCC.n5410 VCC.n5053 0.465115
R48139 VCC.n6519 VCC.n6162 0.465115
R48140 VCC.n7628 VCC.n7271 0.465115
R48141 VCC.n8737 VCC.n8380 0.465115
R48142 VCC.n9846 VCC.n9489 0.465115
R48143 VCC.n10953 VCC.n10596 0.465115
R48144 VCC.n12060 VCC.n11703 0.465115
R48145 VCC.n13167 VCC.n12810 0.465115
R48146 VCC.n14274 VCC.n13917 0.465115
R48147 VCC.n15381 VCC.n15024 0.465115
R48148 VCC.n16488 VCC.n16131 0.465115
R48149 VCC.n17408 VCC.n17238 0.465115
R48150 VCC.n249 VCC.n248 0.366214
R48151 VCC.n468 VCC.n54 0.366214
R48152 VCC.n531 VCC.n529 0.366214
R48153 VCC.n801 VCC.n800 0.366214
R48154 VCC.n1020 VCC.n606 0.366214
R48155 VCC.n1083 VCC.n1081 0.366214
R48156 VCC.n1578 VCC.n1577 0.366214
R48157 VCC.n1649 VCC.n1648 0.366214
R48158 VCC.n1359 VCC.n1358 0.366214
R48159 VCC.n1910 VCC.n1909 0.366214
R48160 VCC.n2129 VCC.n1715 0.366214
R48161 VCC.n2192 VCC.n2190 0.366214
R48162 VCC.n2687 VCC.n2686 0.366214
R48163 VCC.n2758 VCC.n2757 0.366214
R48164 VCC.n2468 VCC.n2467 0.366214
R48165 VCC.n3019 VCC.n3018 0.366214
R48166 VCC.n3238 VCC.n2824 0.366214
R48167 VCC.n3301 VCC.n3299 0.366214
R48168 VCC.n3796 VCC.n3795 0.366214
R48169 VCC.n3867 VCC.n3866 0.366214
R48170 VCC.n3577 VCC.n3576 0.366214
R48171 VCC.n4128 VCC.n4127 0.366214
R48172 VCC.n4347 VCC.n3933 0.366214
R48173 VCC.n4410 VCC.n4408 0.366214
R48174 VCC.n4905 VCC.n4904 0.366214
R48175 VCC.n4976 VCC.n4975 0.366214
R48176 VCC.n4686 VCC.n4685 0.366214
R48177 VCC.n5237 VCC.n5236 0.366214
R48178 VCC.n5456 VCC.n5042 0.366214
R48179 VCC.n5519 VCC.n5517 0.366214
R48180 VCC.n6014 VCC.n6013 0.366214
R48181 VCC.n6085 VCC.n6084 0.366214
R48182 VCC.n5795 VCC.n5794 0.366214
R48183 VCC.n6346 VCC.n6345 0.366214
R48184 VCC.n6565 VCC.n6151 0.366214
R48185 VCC.n6628 VCC.n6626 0.366214
R48186 VCC.n7123 VCC.n7122 0.366214
R48187 VCC.n7194 VCC.n7193 0.366214
R48188 VCC.n6904 VCC.n6903 0.366214
R48189 VCC.n7455 VCC.n7454 0.366214
R48190 VCC.n7674 VCC.n7260 0.366214
R48191 VCC.n7737 VCC.n7735 0.366214
R48192 VCC.n8232 VCC.n8231 0.366214
R48193 VCC.n8303 VCC.n8302 0.366214
R48194 VCC.n8013 VCC.n8012 0.366214
R48195 VCC.n8783 VCC.n8369 0.366214
R48196 VCC.n8846 VCC.n8844 0.366214
R48197 VCC.n8564 VCC.n8563 0.366214
R48198 VCC.n9341 VCC.n9340 0.366214
R48199 VCC.n9412 VCC.n9411 0.366214
R48200 VCC.n9122 VCC.n9121 0.366214
R48201 VCC.n9673 VCC.n9672 0.366214
R48202 VCC.n9892 VCC.n9478 0.366214
R48203 VCC.n9955 VCC.n9953 0.366214
R48204 VCC.n10449 VCC.n10448 0.366214
R48205 VCC.n10520 VCC.n10519 0.366214
R48206 VCC.n10230 VCC.n10229 0.366214
R48207 VCC.n10780 VCC.n10779 0.366214
R48208 VCC.n10999 VCC.n10585 0.366214
R48209 VCC.n11062 VCC.n11060 0.366214
R48210 VCC.n11556 VCC.n11555 0.366214
R48211 VCC.n11627 VCC.n11626 0.366214
R48212 VCC.n11337 VCC.n11336 0.366214
R48213 VCC.n11887 VCC.n11886 0.366214
R48214 VCC.n12106 VCC.n11692 0.366214
R48215 VCC.n12169 VCC.n12167 0.366214
R48216 VCC.n12663 VCC.n12662 0.366214
R48217 VCC.n12734 VCC.n12733 0.366214
R48218 VCC.n12444 VCC.n12443 0.366214
R48219 VCC.n12994 VCC.n12993 0.366214
R48220 VCC.n13213 VCC.n12799 0.366214
R48221 VCC.n13276 VCC.n13274 0.366214
R48222 VCC.n13770 VCC.n13769 0.366214
R48223 VCC.n13841 VCC.n13840 0.366214
R48224 VCC.n13551 VCC.n13550 0.366214
R48225 VCC.n14101 VCC.n14100 0.366214
R48226 VCC.n14320 VCC.n13906 0.366214
R48227 VCC.n14383 VCC.n14381 0.366214
R48228 VCC.n14877 VCC.n14876 0.366214
R48229 VCC.n14948 VCC.n14947 0.366214
R48230 VCC.n14658 VCC.n14657 0.366214
R48231 VCC.n15208 VCC.n15207 0.366214
R48232 VCC.n15427 VCC.n15013 0.366214
R48233 VCC.n15490 VCC.n15488 0.366214
R48234 VCC.n15984 VCC.n15983 0.366214
R48235 VCC.n16055 VCC.n16054 0.366214
R48236 VCC.n15765 VCC.n15764 0.366214
R48237 VCC.n16315 VCC.n16314 0.366214
R48238 VCC.n16534 VCC.n16120 0.366214
R48239 VCC.n16597 VCC.n16595 0.366214
R48240 VCC.n17091 VCC.n17090 0.366214
R48241 VCC.n17162 VCC.n17161 0.366214
R48242 VCC.n16872 VCC.n16871 0.366214
R48243 VCC.n17454 VCC.n17227 0.366214
R48244 VCC.n17517 VCC.n17515 0.366214
R48245 VCC VCC.n553 0.338784
R48246 VCC VCC.n2771 0.338735
R48247 VCC VCC.n4989 0.338735
R48248 VCC VCC.n7207 0.338735
R48249 VCC VCC.n9425 0.338735
R48250 VCC.n17551 VCC 0.338735
R48251 VCC.n17547 VCC 0.338735
R48252 VCC.n17543 VCC 0.338735
R48253 VCC.n2771 VCC 0.309324
R48254 VCC.n7207 VCC 0.309324
R48255 VCC VCC.n17551 0.309324
R48256 VCC VCC.n17543 0.309324
R48257 VCC VCC.n552 0.300964
R48258 VCC VCC.n1106 0.300964
R48259 VCC VCC.n1660 0.300964
R48260 VCC VCC.n2215 0.300964
R48261 VCC VCC.n2769 0.300964
R48262 VCC VCC.n3324 0.300964
R48263 VCC VCC.n3878 0.300964
R48264 VCC VCC.n4433 0.300964
R48265 VCC VCC.n4987 0.300964
R48266 VCC VCC.n5542 0.300964
R48267 VCC VCC.n6096 0.300964
R48268 VCC VCC.n6651 0.300964
R48269 VCC VCC.n7205 0.300964
R48270 VCC VCC.n7760 0.300964
R48271 VCC VCC.n8314 0.300964
R48272 VCC VCC.n8869 0.300964
R48273 VCC VCC.n9423 0.300964
R48274 VCC VCC.n9978 0.300964
R48275 VCC VCC.n10531 0.300964
R48276 VCC VCC.n11085 0.300964
R48277 VCC VCC.n11638 0.300964
R48278 VCC VCC.n12192 0.300964
R48279 VCC VCC.n12745 0.300964
R48280 VCC VCC.n13299 0.300964
R48281 VCC VCC.n13852 0.300964
R48282 VCC VCC.n14406 0.300964
R48283 VCC VCC.n14959 0.300964
R48284 VCC VCC.n15513 0.300964
R48285 VCC VCC.n16066 0.300964
R48286 VCC VCC.n16620 0.300964
R48287 VCC VCC.n17173 0.300964
R48288 VCC VCC.n17540 0.300964
R48289 VCC.n191 VCC 0.294921
R48290 VCC.n743 VCC 0.294921
R48291 VCC.n1301 VCC 0.294921
R48292 VCC.n1852 VCC 0.294921
R48293 VCC.n2410 VCC 0.294921
R48294 VCC.n2961 VCC 0.294921
R48295 VCC.n3519 VCC 0.294921
R48296 VCC.n4070 VCC 0.294921
R48297 VCC.n4628 VCC 0.294921
R48298 VCC.n5179 VCC 0.294921
R48299 VCC.n5737 VCC 0.294921
R48300 VCC.n6288 VCC 0.294921
R48301 VCC.n6846 VCC 0.294921
R48302 VCC.n7397 VCC 0.294921
R48303 VCC.n7955 VCC 0.294921
R48304 VCC.n9064 VCC 0.294921
R48305 VCC.n9615 VCC 0.294921
R48306 VCC.n10172 VCC 0.294921
R48307 VCC.n10722 VCC 0.294921
R48308 VCC.n11279 VCC 0.294921
R48309 VCC.n11829 VCC 0.294921
R48310 VCC.n12386 VCC 0.294921
R48311 VCC.n12936 VCC 0.294921
R48312 VCC.n13493 VCC 0.294921
R48313 VCC.n14043 VCC 0.294921
R48314 VCC.n14600 VCC 0.294921
R48315 VCC.n15150 VCC 0.294921
R48316 VCC.n15707 VCC 0.294921
R48317 VCC.n16257 VCC 0.294921
R48318 VCC.n16814 VCC 0.294921
R48319 VCC.n17301 VCC 0.294921
R48320 VCC.n8506 VCC 0.292833
R48321 VCC.n315 VCC 0.287536
R48322 VCC.n867 VCC 0.287536
R48323 VCC.n1425 VCC 0.287536
R48324 VCC.n1976 VCC 0.287536
R48325 VCC.n2534 VCC 0.287536
R48326 VCC.n3085 VCC 0.287536
R48327 VCC.n3643 VCC 0.287536
R48328 VCC.n4194 VCC 0.287536
R48329 VCC.n4752 VCC 0.287536
R48330 VCC.n5303 VCC 0.287536
R48331 VCC.n5861 VCC 0.287536
R48332 VCC.n6412 VCC 0.287536
R48333 VCC.n6970 VCC 0.287536
R48334 VCC.n7521 VCC 0.287536
R48335 VCC.n8079 VCC 0.287536
R48336 VCC.n8630 VCC 0.287536
R48337 VCC.n9188 VCC 0.287536
R48338 VCC.n9739 VCC 0.287536
R48339 VCC.n10296 VCC 0.287536
R48340 VCC.n10846 VCC 0.287536
R48341 VCC.n11403 VCC 0.287536
R48342 VCC.n11953 VCC 0.287536
R48343 VCC.n12510 VCC 0.287536
R48344 VCC.n13060 VCC 0.287536
R48345 VCC.n13617 VCC 0.287536
R48346 VCC.n14167 VCC 0.287536
R48347 VCC.n14724 VCC 0.287536
R48348 VCC.n15274 VCC 0.287536
R48349 VCC.n15831 VCC 0.287536
R48350 VCC.n16381 VCC 0.287536
R48351 VCC.n16938 VCC 0.287536
R48352 VCC.n224 VCC.n183 0.274786
R48353 VCC.n286 VCC.n141 0.274786
R48354 VCC.n339 VCC.n118 0.274786
R48355 VCC.n365 VCC.n97 0.274786
R48356 VCC.n387 VCC.n95 0.274786
R48357 VCC.n415 VCC.n414 0.274786
R48358 VCC.n776 VCC.n735 0.274786
R48359 VCC.n838 VCC.n693 0.274786
R48360 VCC.n891 VCC.n670 0.274786
R48361 VCC.n917 VCC.n649 0.274786
R48362 VCC.n939 VCC.n647 0.274786
R48363 VCC.n967 VCC.n966 0.274786
R48364 VCC.n1448 VCC.n1227 0.274786
R48365 VCC.n1474 VCC.n1206 0.274786
R48366 VCC.n1496 VCC.n1204 0.274786
R48367 VCC.n1524 VCC.n1523 0.274786
R48368 VCC.n1334 VCC.n1293 0.274786
R48369 VCC.n1396 VCC.n1251 0.274786
R48370 VCC.n1885 VCC.n1844 0.274786
R48371 VCC.n1947 VCC.n1802 0.274786
R48372 VCC.n2000 VCC.n1779 0.274786
R48373 VCC.n2026 VCC.n1758 0.274786
R48374 VCC.n2048 VCC.n1756 0.274786
R48375 VCC.n2076 VCC.n2075 0.274786
R48376 VCC.n2557 VCC.n2336 0.274786
R48377 VCC.n2583 VCC.n2315 0.274786
R48378 VCC.n2605 VCC.n2313 0.274786
R48379 VCC.n2633 VCC.n2632 0.274786
R48380 VCC.n2443 VCC.n2402 0.274786
R48381 VCC.n2505 VCC.n2360 0.274786
R48382 VCC.n2994 VCC.n2953 0.274786
R48383 VCC.n3056 VCC.n2911 0.274786
R48384 VCC.n3109 VCC.n2888 0.274786
R48385 VCC.n3135 VCC.n2867 0.274786
R48386 VCC.n3157 VCC.n2865 0.274786
R48387 VCC.n3185 VCC.n3184 0.274786
R48388 VCC.n3666 VCC.n3445 0.274786
R48389 VCC.n3692 VCC.n3424 0.274786
R48390 VCC.n3714 VCC.n3422 0.274786
R48391 VCC.n3742 VCC.n3741 0.274786
R48392 VCC.n3552 VCC.n3511 0.274786
R48393 VCC.n3614 VCC.n3469 0.274786
R48394 VCC.n4103 VCC.n4062 0.274786
R48395 VCC.n4165 VCC.n4020 0.274786
R48396 VCC.n4218 VCC.n3997 0.274786
R48397 VCC.n4244 VCC.n3976 0.274786
R48398 VCC.n4266 VCC.n3974 0.274786
R48399 VCC.n4294 VCC.n4293 0.274786
R48400 VCC.n4775 VCC.n4554 0.274786
R48401 VCC.n4801 VCC.n4533 0.274786
R48402 VCC.n4823 VCC.n4531 0.274786
R48403 VCC.n4851 VCC.n4850 0.274786
R48404 VCC.n4661 VCC.n4620 0.274786
R48405 VCC.n4723 VCC.n4578 0.274786
R48406 VCC.n5212 VCC.n5171 0.274786
R48407 VCC.n5274 VCC.n5129 0.274786
R48408 VCC.n5327 VCC.n5106 0.274786
R48409 VCC.n5353 VCC.n5085 0.274786
R48410 VCC.n5375 VCC.n5083 0.274786
R48411 VCC.n5403 VCC.n5402 0.274786
R48412 VCC.n5884 VCC.n5663 0.274786
R48413 VCC.n5910 VCC.n5642 0.274786
R48414 VCC.n5932 VCC.n5640 0.274786
R48415 VCC.n5960 VCC.n5959 0.274786
R48416 VCC.n5770 VCC.n5729 0.274786
R48417 VCC.n5832 VCC.n5687 0.274786
R48418 VCC.n6321 VCC.n6280 0.274786
R48419 VCC.n6383 VCC.n6238 0.274786
R48420 VCC.n6436 VCC.n6215 0.274786
R48421 VCC.n6462 VCC.n6194 0.274786
R48422 VCC.n6484 VCC.n6192 0.274786
R48423 VCC.n6512 VCC.n6511 0.274786
R48424 VCC.n6993 VCC.n6772 0.274786
R48425 VCC.n7019 VCC.n6751 0.274786
R48426 VCC.n7041 VCC.n6749 0.274786
R48427 VCC.n7069 VCC.n7068 0.274786
R48428 VCC.n6879 VCC.n6838 0.274786
R48429 VCC.n6941 VCC.n6796 0.274786
R48430 VCC.n7430 VCC.n7389 0.274786
R48431 VCC.n7492 VCC.n7347 0.274786
R48432 VCC.n7545 VCC.n7324 0.274786
R48433 VCC.n7571 VCC.n7303 0.274786
R48434 VCC.n7593 VCC.n7301 0.274786
R48435 VCC.n7621 VCC.n7620 0.274786
R48436 VCC.n8102 VCC.n7881 0.274786
R48437 VCC.n8128 VCC.n7860 0.274786
R48438 VCC.n8150 VCC.n7858 0.274786
R48439 VCC.n8178 VCC.n8177 0.274786
R48440 VCC.n7988 VCC.n7947 0.274786
R48441 VCC.n8050 VCC.n7905 0.274786
R48442 VCC.n8654 VCC.n8433 0.274786
R48443 VCC.n8680 VCC.n8412 0.274786
R48444 VCC.n8702 VCC.n8410 0.274786
R48445 VCC.n8730 VCC.n8729 0.274786
R48446 VCC.n8539 VCC.n8498 0.274786
R48447 VCC.n8601 VCC.n8456 0.274786
R48448 VCC.n9211 VCC.n8990 0.274786
R48449 VCC.n9237 VCC.n8969 0.274786
R48450 VCC.n9259 VCC.n8967 0.274786
R48451 VCC.n9287 VCC.n9286 0.274786
R48452 VCC.n9097 VCC.n9056 0.274786
R48453 VCC.n9159 VCC.n9014 0.274786
R48454 VCC.n9648 VCC.n9607 0.274786
R48455 VCC.n9710 VCC.n9565 0.274786
R48456 VCC.n9763 VCC.n9542 0.274786
R48457 VCC.n9789 VCC.n9521 0.274786
R48458 VCC.n9811 VCC.n9519 0.274786
R48459 VCC.n9839 VCC.n9838 0.274786
R48460 VCC.n10319 VCC.n10098 0.274786
R48461 VCC.n10345 VCC.n10077 0.274786
R48462 VCC.n10367 VCC.n10075 0.274786
R48463 VCC.n10395 VCC.n10394 0.274786
R48464 VCC.n10205 VCC.n10164 0.274786
R48465 VCC.n10267 VCC.n10122 0.274786
R48466 VCC.n10755 VCC.n10714 0.274786
R48467 VCC.n10817 VCC.n10672 0.274786
R48468 VCC.n10870 VCC.n10649 0.274786
R48469 VCC.n10896 VCC.n10628 0.274786
R48470 VCC.n10918 VCC.n10626 0.274786
R48471 VCC.n10946 VCC.n10945 0.274786
R48472 VCC.n11426 VCC.n11205 0.274786
R48473 VCC.n11452 VCC.n11184 0.274786
R48474 VCC.n11474 VCC.n11182 0.274786
R48475 VCC.n11502 VCC.n11501 0.274786
R48476 VCC.n11312 VCC.n11271 0.274786
R48477 VCC.n11374 VCC.n11229 0.274786
R48478 VCC.n11862 VCC.n11821 0.274786
R48479 VCC.n11924 VCC.n11779 0.274786
R48480 VCC.n11977 VCC.n11756 0.274786
R48481 VCC.n12003 VCC.n11735 0.274786
R48482 VCC.n12025 VCC.n11733 0.274786
R48483 VCC.n12053 VCC.n12052 0.274786
R48484 VCC.n12533 VCC.n12312 0.274786
R48485 VCC.n12559 VCC.n12291 0.274786
R48486 VCC.n12581 VCC.n12289 0.274786
R48487 VCC.n12609 VCC.n12608 0.274786
R48488 VCC.n12419 VCC.n12378 0.274786
R48489 VCC.n12481 VCC.n12336 0.274786
R48490 VCC.n12969 VCC.n12928 0.274786
R48491 VCC.n13031 VCC.n12886 0.274786
R48492 VCC.n13084 VCC.n12863 0.274786
R48493 VCC.n13110 VCC.n12842 0.274786
R48494 VCC.n13132 VCC.n12840 0.274786
R48495 VCC.n13160 VCC.n13159 0.274786
R48496 VCC.n13640 VCC.n13419 0.274786
R48497 VCC.n13666 VCC.n13398 0.274786
R48498 VCC.n13688 VCC.n13396 0.274786
R48499 VCC.n13716 VCC.n13715 0.274786
R48500 VCC.n13526 VCC.n13485 0.274786
R48501 VCC.n13588 VCC.n13443 0.274786
R48502 VCC.n14076 VCC.n14035 0.274786
R48503 VCC.n14138 VCC.n13993 0.274786
R48504 VCC.n14191 VCC.n13970 0.274786
R48505 VCC.n14217 VCC.n13949 0.274786
R48506 VCC.n14239 VCC.n13947 0.274786
R48507 VCC.n14267 VCC.n14266 0.274786
R48508 VCC.n14747 VCC.n14526 0.274786
R48509 VCC.n14773 VCC.n14505 0.274786
R48510 VCC.n14795 VCC.n14503 0.274786
R48511 VCC.n14823 VCC.n14822 0.274786
R48512 VCC.n14633 VCC.n14592 0.274786
R48513 VCC.n14695 VCC.n14550 0.274786
R48514 VCC.n15183 VCC.n15142 0.274786
R48515 VCC.n15245 VCC.n15100 0.274786
R48516 VCC.n15298 VCC.n15077 0.274786
R48517 VCC.n15324 VCC.n15056 0.274786
R48518 VCC.n15346 VCC.n15054 0.274786
R48519 VCC.n15374 VCC.n15373 0.274786
R48520 VCC.n15854 VCC.n15633 0.274786
R48521 VCC.n15880 VCC.n15612 0.274786
R48522 VCC.n15902 VCC.n15610 0.274786
R48523 VCC.n15930 VCC.n15929 0.274786
R48524 VCC.n15740 VCC.n15699 0.274786
R48525 VCC.n15802 VCC.n15657 0.274786
R48526 VCC.n16290 VCC.n16249 0.274786
R48527 VCC.n16352 VCC.n16207 0.274786
R48528 VCC.n16405 VCC.n16184 0.274786
R48529 VCC.n16431 VCC.n16163 0.274786
R48530 VCC.n16453 VCC.n16161 0.274786
R48531 VCC.n16481 VCC.n16480 0.274786
R48532 VCC.n16961 VCC.n16740 0.274786
R48533 VCC.n16987 VCC.n16719 0.274786
R48534 VCC.n17009 VCC.n16717 0.274786
R48535 VCC.n17037 VCC.n17036 0.274786
R48536 VCC.n16847 VCC.n16806 0.274786
R48537 VCC.n16909 VCC.n16764 0.274786
R48538 VCC.n17325 VCC.n17291 0.274786
R48539 VCC.n17351 VCC.n17270 0.274786
R48540 VCC.n17373 VCC.n17268 0.274786
R48541 VCC.n17401 VCC.n17400 0.274786
R48542 VCC VCC.n313 0.213679
R48543 VCC VCC.n865 0.213679
R48544 VCC VCC.n1423 0.213679
R48545 VCC VCC.n1974 0.213679
R48546 VCC VCC.n2532 0.213679
R48547 VCC VCC.n3083 0.213679
R48548 VCC VCC.n3641 0.213679
R48549 VCC VCC.n4192 0.213679
R48550 VCC VCC.n4750 0.213679
R48551 VCC VCC.n5301 0.213679
R48552 VCC VCC.n5859 0.213679
R48553 VCC VCC.n6410 0.213679
R48554 VCC VCC.n6968 0.213679
R48555 VCC VCC.n7519 0.213679
R48556 VCC VCC.n8077 0.213679
R48557 VCC VCC.n9186 0.213679
R48558 VCC VCC.n9737 0.213679
R48559 VCC VCC.n10294 0.213679
R48560 VCC VCC.n10844 0.213679
R48561 VCC VCC.n11401 0.213679
R48562 VCC VCC.n11951 0.213679
R48563 VCC VCC.n12508 0.213679
R48564 VCC VCC.n13058 0.213679
R48565 VCC VCC.n13615 0.213679
R48566 VCC VCC.n14165 0.213679
R48567 VCC VCC.n14722 0.213679
R48568 VCC VCC.n15272 0.213679
R48569 VCC VCC.n15829 0.213679
R48570 VCC VCC.n16379 0.213679
R48571 VCC VCC.n16936 0.213679
R48572 VCC VCC.n8628 0.212167
R48573 VCC.n160 VCC.n156 0.183357
R48574 VCC.n490 VCC.n43 0.183357
R48575 VCC.n491 VCC.n490 0.183357
R48576 VCC.n523 VCC.n24 0.183357
R48577 VCC.n523 VCC.n25 0.183357
R48578 VCC.n712 VCC.n708 0.183357
R48579 VCC.n1042 VCC.n595 0.183357
R48580 VCC.n1043 VCC.n1042 0.183357
R48581 VCC.n1075 VCC.n576 0.183357
R48582 VCC.n1075 VCC.n577 0.183357
R48583 VCC.n1593 VCC.n1587 0.183357
R48584 VCC.n1587 VCC.n1160 0.183357
R48585 VCC.n1623 VCC.n1135 0.183357
R48586 VCC.n1623 VCC.n1141 0.183357
R48587 VCC.n1270 VCC.n1266 0.183357
R48588 VCC.n1821 VCC.n1817 0.183357
R48589 VCC.n2151 VCC.n1704 0.183357
R48590 VCC.n2152 VCC.n2151 0.183357
R48591 VCC.n2184 VCC.n1685 0.183357
R48592 VCC.n2184 VCC.n1686 0.183357
R48593 VCC.n2702 VCC.n2696 0.183357
R48594 VCC.n2696 VCC.n2269 0.183357
R48595 VCC.n2732 VCC.n2244 0.183357
R48596 VCC.n2732 VCC.n2250 0.183357
R48597 VCC.n2379 VCC.n2375 0.183357
R48598 VCC.n2930 VCC.n2926 0.183357
R48599 VCC.n3260 VCC.n2813 0.183357
R48600 VCC.n3261 VCC.n3260 0.183357
R48601 VCC.n3293 VCC.n2794 0.183357
R48602 VCC.n3293 VCC.n2795 0.183357
R48603 VCC.n3811 VCC.n3805 0.183357
R48604 VCC.n3805 VCC.n3378 0.183357
R48605 VCC.n3841 VCC.n3353 0.183357
R48606 VCC.n3841 VCC.n3359 0.183357
R48607 VCC.n3488 VCC.n3484 0.183357
R48608 VCC.n4039 VCC.n4035 0.183357
R48609 VCC.n4369 VCC.n3922 0.183357
R48610 VCC.n4370 VCC.n4369 0.183357
R48611 VCC.n4402 VCC.n3903 0.183357
R48612 VCC.n4402 VCC.n3904 0.183357
R48613 VCC.n4920 VCC.n4914 0.183357
R48614 VCC.n4914 VCC.n4487 0.183357
R48615 VCC.n4950 VCC.n4462 0.183357
R48616 VCC.n4950 VCC.n4468 0.183357
R48617 VCC.n4597 VCC.n4593 0.183357
R48618 VCC.n5148 VCC.n5144 0.183357
R48619 VCC.n5478 VCC.n5031 0.183357
R48620 VCC.n5479 VCC.n5478 0.183357
R48621 VCC.n5511 VCC.n5012 0.183357
R48622 VCC.n5511 VCC.n5013 0.183357
R48623 VCC.n6029 VCC.n6023 0.183357
R48624 VCC.n6023 VCC.n5596 0.183357
R48625 VCC.n6059 VCC.n5571 0.183357
R48626 VCC.n6059 VCC.n5577 0.183357
R48627 VCC.n5706 VCC.n5702 0.183357
R48628 VCC.n6257 VCC.n6253 0.183357
R48629 VCC.n6587 VCC.n6140 0.183357
R48630 VCC.n6588 VCC.n6587 0.183357
R48631 VCC.n6620 VCC.n6121 0.183357
R48632 VCC.n6620 VCC.n6122 0.183357
R48633 VCC.n7138 VCC.n7132 0.183357
R48634 VCC.n7132 VCC.n6705 0.183357
R48635 VCC.n7168 VCC.n6680 0.183357
R48636 VCC.n7168 VCC.n6686 0.183357
R48637 VCC.n6815 VCC.n6811 0.183357
R48638 VCC.n7366 VCC.n7362 0.183357
R48639 VCC.n7696 VCC.n7249 0.183357
R48640 VCC.n7697 VCC.n7696 0.183357
R48641 VCC.n7729 VCC.n7230 0.183357
R48642 VCC.n7729 VCC.n7231 0.183357
R48643 VCC.n8247 VCC.n8241 0.183357
R48644 VCC.n8241 VCC.n7814 0.183357
R48645 VCC.n8277 VCC.n7789 0.183357
R48646 VCC.n8277 VCC.n7795 0.183357
R48647 VCC.n7924 VCC.n7920 0.183357
R48648 VCC.n8805 VCC.n8358 0.183357
R48649 VCC.n8806 VCC.n8805 0.183357
R48650 VCC.n8838 VCC.n8339 0.183357
R48651 VCC.n8838 VCC.n8340 0.183357
R48652 VCC.n8475 VCC.n8471 0.183357
R48653 VCC.n9356 VCC.n9350 0.183357
R48654 VCC.n9350 VCC.n8923 0.183357
R48655 VCC.n9386 VCC.n8898 0.183357
R48656 VCC.n9386 VCC.n8904 0.183357
R48657 VCC.n9033 VCC.n9029 0.183357
R48658 VCC.n9584 VCC.n9580 0.183357
R48659 VCC.n9914 VCC.n9467 0.183357
R48660 VCC.n9915 VCC.n9914 0.183357
R48661 VCC.n9947 VCC.n9448 0.183357
R48662 VCC.n9947 VCC.n9449 0.183357
R48663 VCC.n10464 VCC.n10458 0.183357
R48664 VCC.n10458 VCC.n10031 0.183357
R48665 VCC.n10494 VCC.n10006 0.183357
R48666 VCC.n10494 VCC.n10012 0.183357
R48667 VCC.n10141 VCC.n10137 0.183357
R48668 VCC.n10691 VCC.n10687 0.183357
R48669 VCC.n11021 VCC.n10574 0.183357
R48670 VCC.n11022 VCC.n11021 0.183357
R48671 VCC.n11054 VCC.n10555 0.183357
R48672 VCC.n11054 VCC.n10556 0.183357
R48673 VCC.n11571 VCC.n11565 0.183357
R48674 VCC.n11565 VCC.n11138 0.183357
R48675 VCC.n11601 VCC.n11113 0.183357
R48676 VCC.n11601 VCC.n11119 0.183357
R48677 VCC.n11248 VCC.n11244 0.183357
R48678 VCC.n11798 VCC.n11794 0.183357
R48679 VCC.n12128 VCC.n11681 0.183357
R48680 VCC.n12129 VCC.n12128 0.183357
R48681 VCC.n12161 VCC.n11662 0.183357
R48682 VCC.n12161 VCC.n11663 0.183357
R48683 VCC.n12678 VCC.n12672 0.183357
R48684 VCC.n12672 VCC.n12245 0.183357
R48685 VCC.n12708 VCC.n12220 0.183357
R48686 VCC.n12708 VCC.n12226 0.183357
R48687 VCC.n12355 VCC.n12351 0.183357
R48688 VCC.n12905 VCC.n12901 0.183357
R48689 VCC.n13235 VCC.n12788 0.183357
R48690 VCC.n13236 VCC.n13235 0.183357
R48691 VCC.n13268 VCC.n12769 0.183357
R48692 VCC.n13268 VCC.n12770 0.183357
R48693 VCC.n13785 VCC.n13779 0.183357
R48694 VCC.n13779 VCC.n13352 0.183357
R48695 VCC.n13815 VCC.n13327 0.183357
R48696 VCC.n13815 VCC.n13333 0.183357
R48697 VCC.n13462 VCC.n13458 0.183357
R48698 VCC.n14012 VCC.n14008 0.183357
R48699 VCC.n14342 VCC.n13895 0.183357
R48700 VCC.n14343 VCC.n14342 0.183357
R48701 VCC.n14375 VCC.n13876 0.183357
R48702 VCC.n14375 VCC.n13877 0.183357
R48703 VCC.n14892 VCC.n14886 0.183357
R48704 VCC.n14886 VCC.n14459 0.183357
R48705 VCC.n14922 VCC.n14434 0.183357
R48706 VCC.n14922 VCC.n14440 0.183357
R48707 VCC.n14569 VCC.n14565 0.183357
R48708 VCC.n15119 VCC.n15115 0.183357
R48709 VCC.n15449 VCC.n15002 0.183357
R48710 VCC.n15450 VCC.n15449 0.183357
R48711 VCC.n15482 VCC.n14983 0.183357
R48712 VCC.n15482 VCC.n14984 0.183357
R48713 VCC.n15999 VCC.n15993 0.183357
R48714 VCC.n15993 VCC.n15566 0.183357
R48715 VCC.n16029 VCC.n15541 0.183357
R48716 VCC.n16029 VCC.n15547 0.183357
R48717 VCC.n15676 VCC.n15672 0.183357
R48718 VCC.n16226 VCC.n16222 0.183357
R48719 VCC.n16556 VCC.n16109 0.183357
R48720 VCC.n16557 VCC.n16556 0.183357
R48721 VCC.n16589 VCC.n16090 0.183357
R48722 VCC.n16589 VCC.n16091 0.183357
R48723 VCC.n17106 VCC.n17100 0.183357
R48724 VCC.n17100 VCC.n16673 0.183357
R48725 VCC.n17136 VCC.n16648 0.183357
R48726 VCC.n17136 VCC.n16654 0.183357
R48727 VCC.n16783 VCC.n16779 0.183357
R48728 VCC.n17476 VCC.n17216 0.183357
R48729 VCC.n17477 VCC.n17476 0.183357
R48730 VCC.n17509 VCC.n17197 0.183357
R48731 VCC.n17509 VCC.n17198 0.183357
R48732 VCC VCC.n448 0.114307
R48733 VCC VCC.n1000 0.114307
R48734 VCC VCC.n1558 0.114307
R48735 VCC VCC.n2109 0.114307
R48736 VCC VCC.n2667 0.114307
R48737 VCC VCC.n3218 0.114307
R48738 VCC VCC.n3776 0.114307
R48739 VCC VCC.n4327 0.114307
R48740 VCC VCC.n4885 0.114307
R48741 VCC VCC.n5436 0.114307
R48742 VCC VCC.n5994 0.114307
R48743 VCC VCC.n6545 0.114307
R48744 VCC VCC.n7103 0.114307
R48745 VCC VCC.n7654 0.114307
R48746 VCC VCC.n8212 0.114307
R48747 VCC VCC.n8763 0.114307
R48748 VCC VCC.n9321 0.114307
R48749 VCC VCC.n9872 0.114307
R48750 VCC VCC.n10429 0.114307
R48751 VCC VCC.n10979 0.114307
R48752 VCC VCC.n11536 0.114307
R48753 VCC VCC.n12086 0.114307
R48754 VCC VCC.n12643 0.114307
R48755 VCC VCC.n13193 0.114307
R48756 VCC VCC.n13750 0.114307
R48757 VCC VCC.n14300 0.114307
R48758 VCC VCC.n14857 0.114307
R48759 VCC VCC.n15407 0.114307
R48760 VCC VCC.n15964 0.114307
R48761 VCC VCC.n16514 0.114307
R48762 VCC VCC.n17071 0.114307
R48763 VCC VCC.n17434 0.114307
R48764 VCC.n231 VCC.n178 0.0919286
R48765 VCC.n271 VCC.n270 0.0919286
R48766 VCC.n358 VCC.n106 0.0919286
R48767 VCC.n398 VCC.n91 0.0919286
R48768 VCC.n531 VCC.n530 0.0919286
R48769 VCC.n544 VCC.n7 0.0919286
R48770 VCC.n783 VCC.n730 0.0919286
R48771 VCC.n823 VCC.n822 0.0919286
R48772 VCC.n910 VCC.n658 0.0919286
R48773 VCC.n950 VCC.n643 0.0919286
R48774 VCC.n1083 VCC.n1082 0.0919286
R48775 VCC.n1098 VCC.n561 0.0919286
R48776 VCC.n1648 VCC.n1117 0.0919286
R48777 VCC.n1124 VCC.n1123 0.0919286
R48778 VCC.n1467 VCC.n1215 0.0919286
R48779 VCC.n1507 VCC.n1200 0.0919286
R48780 VCC.n1341 VCC.n1288 0.0919286
R48781 VCC.n1381 VCC.n1380 0.0919286
R48782 VCC.n1892 VCC.n1839 0.0919286
R48783 VCC.n1932 VCC.n1931 0.0919286
R48784 VCC.n2019 VCC.n1767 0.0919286
R48785 VCC.n2059 VCC.n1752 0.0919286
R48786 VCC.n2192 VCC.n2191 0.0919286
R48787 VCC.n2207 VCC.n1670 0.0919286
R48788 VCC.n2757 VCC.n2226 0.0919286
R48789 VCC.n2233 VCC.n2232 0.0919286
R48790 VCC.n2576 VCC.n2324 0.0919286
R48791 VCC.n2616 VCC.n2309 0.0919286
R48792 VCC.n2450 VCC.n2397 0.0919286
R48793 VCC.n2490 VCC.n2489 0.0919286
R48794 VCC.n3001 VCC.n2948 0.0919286
R48795 VCC.n3041 VCC.n3040 0.0919286
R48796 VCC.n3128 VCC.n2876 0.0919286
R48797 VCC.n3168 VCC.n2861 0.0919286
R48798 VCC.n3301 VCC.n3300 0.0919286
R48799 VCC.n3316 VCC.n2779 0.0919286
R48800 VCC.n3866 VCC.n3335 0.0919286
R48801 VCC.n3342 VCC.n3341 0.0919286
R48802 VCC.n3685 VCC.n3433 0.0919286
R48803 VCC.n3725 VCC.n3418 0.0919286
R48804 VCC.n3559 VCC.n3506 0.0919286
R48805 VCC.n3599 VCC.n3598 0.0919286
R48806 VCC.n4110 VCC.n4057 0.0919286
R48807 VCC.n4150 VCC.n4149 0.0919286
R48808 VCC.n4237 VCC.n3985 0.0919286
R48809 VCC.n4277 VCC.n3970 0.0919286
R48810 VCC.n4410 VCC.n4409 0.0919286
R48811 VCC.n4425 VCC.n3888 0.0919286
R48812 VCC.n4975 VCC.n4444 0.0919286
R48813 VCC.n4451 VCC.n4450 0.0919286
R48814 VCC.n4794 VCC.n4542 0.0919286
R48815 VCC.n4834 VCC.n4527 0.0919286
R48816 VCC.n4668 VCC.n4615 0.0919286
R48817 VCC.n4708 VCC.n4707 0.0919286
R48818 VCC.n5219 VCC.n5166 0.0919286
R48819 VCC.n5259 VCC.n5258 0.0919286
R48820 VCC.n5346 VCC.n5094 0.0919286
R48821 VCC.n5386 VCC.n5079 0.0919286
R48822 VCC.n5519 VCC.n5518 0.0919286
R48823 VCC.n5534 VCC.n4997 0.0919286
R48824 VCC.n6084 VCC.n5553 0.0919286
R48825 VCC.n5560 VCC.n5559 0.0919286
R48826 VCC.n5903 VCC.n5651 0.0919286
R48827 VCC.n5943 VCC.n5636 0.0919286
R48828 VCC.n5777 VCC.n5724 0.0919286
R48829 VCC.n5817 VCC.n5816 0.0919286
R48830 VCC.n6328 VCC.n6275 0.0919286
R48831 VCC.n6368 VCC.n6367 0.0919286
R48832 VCC.n6455 VCC.n6203 0.0919286
R48833 VCC.n6495 VCC.n6188 0.0919286
R48834 VCC.n6628 VCC.n6627 0.0919286
R48835 VCC.n6643 VCC.n6106 0.0919286
R48836 VCC.n7193 VCC.n6662 0.0919286
R48837 VCC.n6669 VCC.n6668 0.0919286
R48838 VCC.n7012 VCC.n6760 0.0919286
R48839 VCC.n7052 VCC.n6745 0.0919286
R48840 VCC.n6886 VCC.n6833 0.0919286
R48841 VCC.n6926 VCC.n6925 0.0919286
R48842 VCC.n7437 VCC.n7384 0.0919286
R48843 VCC.n7477 VCC.n7476 0.0919286
R48844 VCC.n7564 VCC.n7312 0.0919286
R48845 VCC.n7604 VCC.n7297 0.0919286
R48846 VCC.n7737 VCC.n7736 0.0919286
R48847 VCC.n7752 VCC.n7215 0.0919286
R48848 VCC.n8302 VCC.n7771 0.0919286
R48849 VCC.n7778 VCC.n7777 0.0919286
R48850 VCC.n8121 VCC.n7869 0.0919286
R48851 VCC.n8161 VCC.n7854 0.0919286
R48852 VCC.n7995 VCC.n7942 0.0919286
R48853 VCC.n8035 VCC.n8034 0.0919286
R48854 VCC.n8673 VCC.n8421 0.0919286
R48855 VCC.n8713 VCC.n8406 0.0919286
R48856 VCC.n8846 VCC.n8845 0.0919286
R48857 VCC.n8861 VCC.n8324 0.0919286
R48858 VCC.n8546 VCC.n8493 0.0919286
R48859 VCC.n8586 VCC.n8585 0.0919286
R48860 VCC.n9411 VCC.n8880 0.0919286
R48861 VCC.n8887 VCC.n8886 0.0919286
R48862 VCC.n9230 VCC.n8978 0.0919286
R48863 VCC.n9270 VCC.n8963 0.0919286
R48864 VCC.n9104 VCC.n9051 0.0919286
R48865 VCC.n9144 VCC.n9143 0.0919286
R48866 VCC.n9655 VCC.n9602 0.0919286
R48867 VCC.n9695 VCC.n9694 0.0919286
R48868 VCC.n9782 VCC.n9530 0.0919286
R48869 VCC.n9822 VCC.n9515 0.0919286
R48870 VCC.n9955 VCC.n9954 0.0919286
R48871 VCC.n9970 VCC.n9433 0.0919286
R48872 VCC.n10519 VCC.n9988 0.0919286
R48873 VCC.n9995 VCC.n9994 0.0919286
R48874 VCC.n10338 VCC.n10086 0.0919286
R48875 VCC.n10378 VCC.n10071 0.0919286
R48876 VCC.n10212 VCC.n10159 0.0919286
R48877 VCC.n10252 VCC.n10251 0.0919286
R48878 VCC.n10762 VCC.n10709 0.0919286
R48879 VCC.n10802 VCC.n10801 0.0919286
R48880 VCC.n10889 VCC.n10637 0.0919286
R48881 VCC.n10929 VCC.n10622 0.0919286
R48882 VCC.n11062 VCC.n11061 0.0919286
R48883 VCC.n11077 VCC.n10540 0.0919286
R48884 VCC.n11626 VCC.n11095 0.0919286
R48885 VCC.n11102 VCC.n11101 0.0919286
R48886 VCC.n11445 VCC.n11193 0.0919286
R48887 VCC.n11485 VCC.n11178 0.0919286
R48888 VCC.n11319 VCC.n11266 0.0919286
R48889 VCC.n11359 VCC.n11358 0.0919286
R48890 VCC.n11869 VCC.n11816 0.0919286
R48891 VCC.n11909 VCC.n11908 0.0919286
R48892 VCC.n11996 VCC.n11744 0.0919286
R48893 VCC.n12036 VCC.n11729 0.0919286
R48894 VCC.n12169 VCC.n12168 0.0919286
R48895 VCC.n12184 VCC.n11647 0.0919286
R48896 VCC.n12733 VCC.n12202 0.0919286
R48897 VCC.n12209 VCC.n12208 0.0919286
R48898 VCC.n12552 VCC.n12300 0.0919286
R48899 VCC.n12592 VCC.n12285 0.0919286
R48900 VCC.n12426 VCC.n12373 0.0919286
R48901 VCC.n12466 VCC.n12465 0.0919286
R48902 VCC.n12976 VCC.n12923 0.0919286
R48903 VCC.n13016 VCC.n13015 0.0919286
R48904 VCC.n13103 VCC.n12851 0.0919286
R48905 VCC.n13143 VCC.n12836 0.0919286
R48906 VCC.n13276 VCC.n13275 0.0919286
R48907 VCC.n13291 VCC.n12754 0.0919286
R48908 VCC.n13840 VCC.n13309 0.0919286
R48909 VCC.n13316 VCC.n13315 0.0919286
R48910 VCC.n13659 VCC.n13407 0.0919286
R48911 VCC.n13699 VCC.n13392 0.0919286
R48912 VCC.n13533 VCC.n13480 0.0919286
R48913 VCC.n13573 VCC.n13572 0.0919286
R48914 VCC.n14083 VCC.n14030 0.0919286
R48915 VCC.n14123 VCC.n14122 0.0919286
R48916 VCC.n14210 VCC.n13958 0.0919286
R48917 VCC.n14250 VCC.n13943 0.0919286
R48918 VCC.n14383 VCC.n14382 0.0919286
R48919 VCC.n14398 VCC.n13861 0.0919286
R48920 VCC.n14947 VCC.n14416 0.0919286
R48921 VCC.n14423 VCC.n14422 0.0919286
R48922 VCC.n14766 VCC.n14514 0.0919286
R48923 VCC.n14806 VCC.n14499 0.0919286
R48924 VCC.n14640 VCC.n14587 0.0919286
R48925 VCC.n14680 VCC.n14679 0.0919286
R48926 VCC.n15190 VCC.n15137 0.0919286
R48927 VCC.n15230 VCC.n15229 0.0919286
R48928 VCC.n15317 VCC.n15065 0.0919286
R48929 VCC.n15357 VCC.n15050 0.0919286
R48930 VCC.n15490 VCC.n15489 0.0919286
R48931 VCC.n15505 VCC.n14968 0.0919286
R48932 VCC.n16054 VCC.n15523 0.0919286
R48933 VCC.n15530 VCC.n15529 0.0919286
R48934 VCC.n15873 VCC.n15621 0.0919286
R48935 VCC.n15913 VCC.n15606 0.0919286
R48936 VCC.n15747 VCC.n15694 0.0919286
R48937 VCC.n15787 VCC.n15786 0.0919286
R48938 VCC.n16297 VCC.n16244 0.0919286
R48939 VCC.n16337 VCC.n16336 0.0919286
R48940 VCC.n16424 VCC.n16172 0.0919286
R48941 VCC.n16464 VCC.n16157 0.0919286
R48942 VCC.n16597 VCC.n16596 0.0919286
R48943 VCC.n16612 VCC.n16075 0.0919286
R48944 VCC.n17161 VCC.n16630 0.0919286
R48945 VCC.n16637 VCC.n16636 0.0919286
R48946 VCC.n16980 VCC.n16728 0.0919286
R48947 VCC.n17020 VCC.n16713 0.0919286
R48948 VCC.n16854 VCC.n16801 0.0919286
R48949 VCC.n16894 VCC.n16893 0.0919286
R48950 VCC.n17344 VCC.n17279 0.0919286
R48951 VCC.n17384 VCC.n17264 0.0919286
R48952 VCC.n17517 VCC.n17516 0.0919286
R48953 VCC.n17532 VCC.n17182 0.0919286
R48954 VCC.n1107 VCC 0.0247197
R48955 VCC.n2216 VCC 0.0247197
R48956 VCC.n3325 VCC 0.0247197
R48957 VCC.n4434 VCC 0.0247197
R48958 VCC.n5543 VCC 0.0247197
R48959 VCC.n6652 VCC 0.0247197
R48960 VCC.n7761 VCC 0.0247197
R48961 VCC.n8870 VCC 0.0247197
R48962 VCC.n17554 VCC 0.0247197
R48963 VCC.n17552 VCC 0.0247197
R48964 VCC.n17550 VCC 0.0247197
R48965 VCC.n17548 VCC 0.0247197
R48966 VCC.n17546 VCC 0.0247197
R48967 VCC.n17544 VCC 0.0247197
R48968 VCC.n17542 VCC 0.0247197
R48969 VCC.n553 VCC 0.0246714
R48970 VCC.n1661 VCC 0.0246714
R48971 VCC.n2770 VCC 0.0246714
R48972 VCC.n3879 VCC 0.0246714
R48973 VCC.n4988 VCC 0.0246714
R48974 VCC.n6097 VCC 0.0246714
R48975 VCC.n7206 VCC 0.0246714
R48976 VCC.n8315 VCC 0.0246714
R48977 VCC.n9424 VCC 0.0246714
R48978 VCC.n10532 VCC 0.0246714
R48979 VCC.n11639 VCC 0.0246714
R48980 VCC.n12746 VCC 0.0246714
R48981 VCC.n13853 VCC 0.0246714
R48982 VCC.n14960 VCC 0.0246714
R48983 VCC.n16067 VCC 0.0246714
R48984 VCC.n17174 VCC 0.0246714
R48985 VCC.n218 VCC.n217 0.024
R48986 VCC.n308 VCC.n307 0.024
R48987 VCC.n317 VCC.n114 0.024
R48988 VCC.n443 VCC.n442 0.024
R48989 VCC.n461 VCC.n460 0.024
R48990 VCC.n537 VCC.n536 0.024
R48991 VCC.n770 VCC.n769 0.024
R48992 VCC.n860 VCC.n859 0.024
R48993 VCC.n869 VCC.n666 0.024
R48994 VCC.n995 VCC.n994 0.024
R48995 VCC.n1013 VCC.n1012 0.024
R48996 VCC.n1089 VCC.n1088 0.024
R48997 VCC.n1328 VCC.n1327 0.024
R48998 VCC.n1418 VCC.n1417 0.024
R48999 VCC.n1427 VCC.n1223 0.024
R49000 VCC.n1553 VCC.n1552 0.024
R49001 VCC.n1572 VCC.n1571 0.024
R49002 VCC.n1636 VCC.n1635 0.024
R49003 VCC.n1879 VCC.n1878 0.024
R49004 VCC.n1969 VCC.n1968 0.024
R49005 VCC.n1978 VCC.n1775 0.024
R49006 VCC.n2104 VCC.n2103 0.024
R49007 VCC.n2122 VCC.n2121 0.024
R49008 VCC.n2198 VCC.n2197 0.024
R49009 VCC.n2437 VCC.n2436 0.024
R49010 VCC.n2527 VCC.n2526 0.024
R49011 VCC.n2536 VCC.n2332 0.024
R49012 VCC.n2662 VCC.n2661 0.024
R49013 VCC.n2681 VCC.n2680 0.024
R49014 VCC.n2745 VCC.n2744 0.024
R49015 VCC.n2988 VCC.n2987 0.024
R49016 VCC.n3078 VCC.n3077 0.024
R49017 VCC.n3087 VCC.n2884 0.024
R49018 VCC.n3213 VCC.n3212 0.024
R49019 VCC.n3231 VCC.n3230 0.024
R49020 VCC.n3307 VCC.n3306 0.024
R49021 VCC.n3546 VCC.n3545 0.024
R49022 VCC.n3636 VCC.n3635 0.024
R49023 VCC.n3645 VCC.n3441 0.024
R49024 VCC.n3771 VCC.n3770 0.024
R49025 VCC.n3790 VCC.n3789 0.024
R49026 VCC.n3854 VCC.n3853 0.024
R49027 VCC.n4097 VCC.n4096 0.024
R49028 VCC.n4187 VCC.n4186 0.024
R49029 VCC.n4196 VCC.n3993 0.024
R49030 VCC.n4322 VCC.n4321 0.024
R49031 VCC.n4340 VCC.n4339 0.024
R49032 VCC.n4416 VCC.n4415 0.024
R49033 VCC.n4655 VCC.n4654 0.024
R49034 VCC.n4745 VCC.n4744 0.024
R49035 VCC.n4754 VCC.n4550 0.024
R49036 VCC.n4880 VCC.n4879 0.024
R49037 VCC.n4899 VCC.n4898 0.024
R49038 VCC.n4963 VCC.n4962 0.024
R49039 VCC.n5206 VCC.n5205 0.024
R49040 VCC.n5296 VCC.n5295 0.024
R49041 VCC.n5305 VCC.n5102 0.024
R49042 VCC.n5431 VCC.n5430 0.024
R49043 VCC.n5449 VCC.n5448 0.024
R49044 VCC.n5525 VCC.n5524 0.024
R49045 VCC.n5764 VCC.n5763 0.024
R49046 VCC.n5854 VCC.n5853 0.024
R49047 VCC.n5863 VCC.n5659 0.024
R49048 VCC.n5989 VCC.n5988 0.024
R49049 VCC.n6008 VCC.n6007 0.024
R49050 VCC.n6072 VCC.n6071 0.024
R49051 VCC.n6315 VCC.n6314 0.024
R49052 VCC.n6405 VCC.n6404 0.024
R49053 VCC.n6414 VCC.n6211 0.024
R49054 VCC.n6540 VCC.n6539 0.024
R49055 VCC.n6558 VCC.n6557 0.024
R49056 VCC.n6634 VCC.n6633 0.024
R49057 VCC.n6873 VCC.n6872 0.024
R49058 VCC.n6963 VCC.n6962 0.024
R49059 VCC.n6972 VCC.n6768 0.024
R49060 VCC.n7098 VCC.n7097 0.024
R49061 VCC.n7117 VCC.n7116 0.024
R49062 VCC.n7181 VCC.n7180 0.024
R49063 VCC.n7424 VCC.n7423 0.024
R49064 VCC.n7514 VCC.n7513 0.024
R49065 VCC.n7523 VCC.n7320 0.024
R49066 VCC.n7649 VCC.n7648 0.024
R49067 VCC.n7667 VCC.n7666 0.024
R49068 VCC.n7743 VCC.n7742 0.024
R49069 VCC.n7982 VCC.n7981 0.024
R49070 VCC.n8072 VCC.n8071 0.024
R49071 VCC.n8081 VCC.n7877 0.024
R49072 VCC.n8207 VCC.n8206 0.024
R49073 VCC.n8226 VCC.n8225 0.024
R49074 VCC.n8290 VCC.n8289 0.024
R49075 VCC.n8632 VCC.n8429 0.024
R49076 VCC.n8758 VCC.n8757 0.024
R49077 VCC.n8776 VCC.n8775 0.024
R49078 VCC.n8852 VCC.n8851 0.024
R49079 VCC.n9091 VCC.n9090 0.024
R49080 VCC.n9181 VCC.n9180 0.024
R49081 VCC.n9190 VCC.n8986 0.024
R49082 VCC.n9316 VCC.n9315 0.024
R49083 VCC.n9335 VCC.n9334 0.024
R49084 VCC.n9399 VCC.n9398 0.024
R49085 VCC.n9642 VCC.n9641 0.024
R49086 VCC.n9732 VCC.n9731 0.024
R49087 VCC.n9741 VCC.n9538 0.024
R49088 VCC.n9867 VCC.n9866 0.024
R49089 VCC.n9885 VCC.n9884 0.024
R49090 VCC.n9961 VCC.n9960 0.024
R49091 VCC.n10199 VCC.n10198 0.024
R49092 VCC.n10289 VCC.n10288 0.024
R49093 VCC.n10298 VCC.n10094 0.024
R49094 VCC.n10424 VCC.n10423 0.024
R49095 VCC.n10443 VCC.n10442 0.024
R49096 VCC.n10507 VCC.n10506 0.024
R49097 VCC.n10749 VCC.n10748 0.024
R49098 VCC.n10839 VCC.n10838 0.024
R49099 VCC.n10848 VCC.n10645 0.024
R49100 VCC.n10974 VCC.n10973 0.024
R49101 VCC.n10992 VCC.n10991 0.024
R49102 VCC.n11068 VCC.n11067 0.024
R49103 VCC.n11306 VCC.n11305 0.024
R49104 VCC.n11396 VCC.n11395 0.024
R49105 VCC.n11405 VCC.n11201 0.024
R49106 VCC.n11531 VCC.n11530 0.024
R49107 VCC.n11550 VCC.n11549 0.024
R49108 VCC.n11614 VCC.n11613 0.024
R49109 VCC.n11856 VCC.n11855 0.024
R49110 VCC.n11946 VCC.n11945 0.024
R49111 VCC.n11955 VCC.n11752 0.024
R49112 VCC.n12081 VCC.n12080 0.024
R49113 VCC.n12099 VCC.n12098 0.024
R49114 VCC.n12175 VCC.n12174 0.024
R49115 VCC.n12413 VCC.n12412 0.024
R49116 VCC.n12503 VCC.n12502 0.024
R49117 VCC.n12512 VCC.n12308 0.024
R49118 VCC.n12638 VCC.n12637 0.024
R49119 VCC.n12657 VCC.n12656 0.024
R49120 VCC.n12721 VCC.n12720 0.024
R49121 VCC.n12963 VCC.n12962 0.024
R49122 VCC.n13053 VCC.n13052 0.024
R49123 VCC.n13062 VCC.n12859 0.024
R49124 VCC.n13188 VCC.n13187 0.024
R49125 VCC.n13206 VCC.n13205 0.024
R49126 VCC.n13282 VCC.n13281 0.024
R49127 VCC.n13520 VCC.n13519 0.024
R49128 VCC.n13610 VCC.n13609 0.024
R49129 VCC.n13619 VCC.n13415 0.024
R49130 VCC.n13745 VCC.n13744 0.024
R49131 VCC.n13764 VCC.n13763 0.024
R49132 VCC.n13828 VCC.n13827 0.024
R49133 VCC.n14070 VCC.n14069 0.024
R49134 VCC.n14160 VCC.n14159 0.024
R49135 VCC.n14169 VCC.n13966 0.024
R49136 VCC.n14295 VCC.n14294 0.024
R49137 VCC.n14313 VCC.n14312 0.024
R49138 VCC.n14389 VCC.n14388 0.024
R49139 VCC.n14627 VCC.n14626 0.024
R49140 VCC.n14717 VCC.n14716 0.024
R49141 VCC.n14726 VCC.n14522 0.024
R49142 VCC.n14852 VCC.n14851 0.024
R49143 VCC.n14871 VCC.n14870 0.024
R49144 VCC.n14935 VCC.n14934 0.024
R49145 VCC.n15177 VCC.n15176 0.024
R49146 VCC.n15267 VCC.n15266 0.024
R49147 VCC.n15276 VCC.n15073 0.024
R49148 VCC.n15402 VCC.n15401 0.024
R49149 VCC.n15420 VCC.n15419 0.024
R49150 VCC.n15496 VCC.n15495 0.024
R49151 VCC.n15734 VCC.n15733 0.024
R49152 VCC.n15824 VCC.n15823 0.024
R49153 VCC.n15833 VCC.n15629 0.024
R49154 VCC.n15959 VCC.n15958 0.024
R49155 VCC.n15978 VCC.n15977 0.024
R49156 VCC.n16042 VCC.n16041 0.024
R49157 VCC.n16284 VCC.n16283 0.024
R49158 VCC.n16374 VCC.n16373 0.024
R49159 VCC.n16383 VCC.n16180 0.024
R49160 VCC.n16509 VCC.n16508 0.024
R49161 VCC.n16527 VCC.n16526 0.024
R49162 VCC.n16603 VCC.n16602 0.024
R49163 VCC.n16841 VCC.n16840 0.024
R49164 VCC.n16931 VCC.n16930 0.024
R49165 VCC.n16940 VCC.n16736 0.024
R49166 VCC.n17066 VCC.n17065 0.024
R49167 VCC.n17085 VCC.n17084 0.024
R49168 VCC.n17149 VCC.n17148 0.024
R49169 VCC.n17303 VCC.n17287 0.024
R49170 VCC.n17429 VCC.n17428 0.024
R49171 VCC.n17447 VCC.n17446 0.024
R49172 VCC.n17523 VCC.n17522 0.024
R49173 VCC.n8533 VCC.n8532 0.0238333
R49174 VCC.n8623 VCC.n8622 0.0238333
R49175 VCC.n47 VCC.n38 0.0228214
R49176 VCC.n509 VCC.n508 0.0228214
R49177 VCC.n517 VCC.n16 0.0228214
R49178 VCC.n599 VCC.n590 0.0228214
R49179 VCC.n1061 VCC.n1060 0.0228214
R49180 VCC.n1069 VCC.n568 0.0228214
R49181 VCC.n1605 VCC.n1604 0.0228214
R49182 VCC.n1148 VCC.n1133 0.0228214
R49183 VCC.n1632 VCC.n1128 0.0228214
R49184 VCC.n1708 VCC.n1699 0.0228214
R49185 VCC.n2170 VCC.n2169 0.0228214
R49186 VCC.n2178 VCC.n1677 0.0228214
R49187 VCC.n2714 VCC.n2713 0.0228214
R49188 VCC.n2257 VCC.n2242 0.0228214
R49189 VCC.n2741 VCC.n2237 0.0228214
R49190 VCC.n2817 VCC.n2808 0.0228214
R49191 VCC.n3279 VCC.n3278 0.0228214
R49192 VCC.n3287 VCC.n2786 0.0228214
R49193 VCC.n3823 VCC.n3822 0.0228214
R49194 VCC.n3366 VCC.n3351 0.0228214
R49195 VCC.n3850 VCC.n3346 0.0228214
R49196 VCC.n3926 VCC.n3917 0.0228214
R49197 VCC.n4388 VCC.n4387 0.0228214
R49198 VCC.n4396 VCC.n3895 0.0228214
R49199 VCC.n4932 VCC.n4931 0.0228214
R49200 VCC.n4475 VCC.n4460 0.0228214
R49201 VCC.n4959 VCC.n4455 0.0228214
R49202 VCC.n5035 VCC.n5026 0.0228214
R49203 VCC.n5497 VCC.n5496 0.0228214
R49204 VCC.n5505 VCC.n5004 0.0228214
R49205 VCC.n6041 VCC.n6040 0.0228214
R49206 VCC.n5584 VCC.n5569 0.0228214
R49207 VCC.n6068 VCC.n5564 0.0228214
R49208 VCC.n6144 VCC.n6135 0.0228214
R49209 VCC.n6606 VCC.n6605 0.0228214
R49210 VCC.n6614 VCC.n6113 0.0228214
R49211 VCC.n7150 VCC.n7149 0.0228214
R49212 VCC.n6693 VCC.n6678 0.0228214
R49213 VCC.n7177 VCC.n6673 0.0228214
R49214 VCC.n7253 VCC.n7244 0.0228214
R49215 VCC.n7715 VCC.n7714 0.0228214
R49216 VCC.n7723 VCC.n7222 0.0228214
R49217 VCC.n8259 VCC.n8258 0.0228214
R49218 VCC.n7802 VCC.n7787 0.0228214
R49219 VCC.n8286 VCC.n7782 0.0228214
R49220 VCC.n8362 VCC.n8353 0.0228214
R49221 VCC.n8824 VCC.n8823 0.0228214
R49222 VCC.n8832 VCC.n8331 0.0228214
R49223 VCC.n9368 VCC.n9367 0.0228214
R49224 VCC.n8911 VCC.n8896 0.0228214
R49225 VCC.n9395 VCC.n8891 0.0228214
R49226 VCC.n9471 VCC.n9462 0.0228214
R49227 VCC.n9933 VCC.n9932 0.0228214
R49228 VCC.n9941 VCC.n9440 0.0228214
R49229 VCC.n10476 VCC.n10475 0.0228214
R49230 VCC.n10019 VCC.n10004 0.0228214
R49231 VCC.n10503 VCC.n9999 0.0228214
R49232 VCC.n10578 VCC.n10569 0.0228214
R49233 VCC.n11040 VCC.n11039 0.0228214
R49234 VCC.n11048 VCC.n10547 0.0228214
R49235 VCC.n11583 VCC.n11582 0.0228214
R49236 VCC.n11126 VCC.n11111 0.0228214
R49237 VCC.n11610 VCC.n11106 0.0228214
R49238 VCC.n11685 VCC.n11676 0.0228214
R49239 VCC.n12147 VCC.n12146 0.0228214
R49240 VCC.n12155 VCC.n11654 0.0228214
R49241 VCC.n12690 VCC.n12689 0.0228214
R49242 VCC.n12233 VCC.n12218 0.0228214
R49243 VCC.n12717 VCC.n12213 0.0228214
R49244 VCC.n12792 VCC.n12783 0.0228214
R49245 VCC.n13254 VCC.n13253 0.0228214
R49246 VCC.n13262 VCC.n12761 0.0228214
R49247 VCC.n13797 VCC.n13796 0.0228214
R49248 VCC.n13340 VCC.n13325 0.0228214
R49249 VCC.n13824 VCC.n13320 0.0228214
R49250 VCC.n13899 VCC.n13890 0.0228214
R49251 VCC.n14361 VCC.n14360 0.0228214
R49252 VCC.n14369 VCC.n13868 0.0228214
R49253 VCC.n14904 VCC.n14903 0.0228214
R49254 VCC.n14447 VCC.n14432 0.0228214
R49255 VCC.n14931 VCC.n14427 0.0228214
R49256 VCC.n15006 VCC.n14997 0.0228214
R49257 VCC.n15468 VCC.n15467 0.0228214
R49258 VCC.n15476 VCC.n14975 0.0228214
R49259 VCC.n16011 VCC.n16010 0.0228214
R49260 VCC.n15554 VCC.n15539 0.0228214
R49261 VCC.n16038 VCC.n15534 0.0228214
R49262 VCC.n16113 VCC.n16104 0.0228214
R49263 VCC.n16575 VCC.n16574 0.0228214
R49264 VCC.n16583 VCC.n16082 0.0228214
R49265 VCC.n17118 VCC.n17117 0.0228214
R49266 VCC.n16661 VCC.n16646 0.0228214
R49267 VCC.n17145 VCC.n16641 0.0228214
R49268 VCC.n17220 VCC.n17211 0.0228214
R49269 VCC.n17495 VCC.n17494 0.0228214
R49270 VCC.n17503 VCC.n17189 0.0228214
R49271 VCC.n553 VCC 0.0199714
R49272 VCC.n1661 VCC 0.0199714
R49273 VCC.n2770 VCC 0.0199714
R49274 VCC.n3879 VCC 0.0199714
R49275 VCC.n4988 VCC 0.0199714
R49276 VCC.n6097 VCC 0.0199714
R49277 VCC.n7206 VCC 0.0199714
R49278 VCC.n8315 VCC 0.0199714
R49279 VCC.n9424 VCC 0.0199714
R49280 VCC.n10532 VCC 0.0199714
R49281 VCC.n11639 VCC 0.0199714
R49282 VCC.n12746 VCC 0.0199714
R49283 VCC.n13853 VCC 0.0199714
R49284 VCC.n14960 VCC 0.0199714
R49285 VCC.n16067 VCC 0.0199714
R49286 VCC.n17174 VCC 0.0199714
R49287 VCC.n253 VCC.n157 0.0174643
R49288 VCC.n252 VCC.n163 0.0174643
R49289 VCC.n376 VCC.n99 0.0174643
R49290 VCC.n377 VCC.n376 0.0174643
R49291 VCC.n381 VCC.n101 0.0174643
R49292 VCC.n378 VCC.n101 0.0174643
R49293 VCC.n501 VCC.n500 0.0174643
R49294 VCC.n500 VCC.n32 0.0174643
R49295 VCC.n502 VCC.n37 0.0174643
R49296 VCC.n37 VCC.n33 0.0174643
R49297 VCC.n805 VCC.n709 0.0174643
R49298 VCC.n804 VCC.n715 0.0174643
R49299 VCC.n928 VCC.n651 0.0174643
R49300 VCC.n929 VCC.n928 0.0174643
R49301 VCC.n933 VCC.n653 0.0174643
R49302 VCC.n930 VCC.n653 0.0174643
R49303 VCC.n1053 VCC.n1052 0.0174643
R49304 VCC.n1052 VCC.n584 0.0174643
R49305 VCC.n1054 VCC.n589 0.0174643
R49306 VCC.n589 VCC.n585 0.0174643
R49307 VCC.n1615 VCC.n1146 0.0174643
R49308 VCC.n1615 VCC.n1614 0.0174643
R49309 VCC.n1607 VCC.n1147 0.0174643
R49310 VCC.n1613 VCC.n1147 0.0174643
R49311 VCC.n1485 VCC.n1208 0.0174643
R49312 VCC.n1486 VCC.n1485 0.0174643
R49313 VCC.n1490 VCC.n1210 0.0174643
R49314 VCC.n1487 VCC.n1210 0.0174643
R49315 VCC.n1363 VCC.n1267 0.0174643
R49316 VCC.n1362 VCC.n1273 0.0174643
R49317 VCC.n1914 VCC.n1818 0.0174643
R49318 VCC.n1913 VCC.n1824 0.0174643
R49319 VCC.n2037 VCC.n1760 0.0174643
R49320 VCC.n2038 VCC.n2037 0.0174643
R49321 VCC.n2042 VCC.n1762 0.0174643
R49322 VCC.n2039 VCC.n1762 0.0174643
R49323 VCC.n2162 VCC.n2161 0.0174643
R49324 VCC.n2161 VCC.n1693 0.0174643
R49325 VCC.n2163 VCC.n1698 0.0174643
R49326 VCC.n1698 VCC.n1694 0.0174643
R49327 VCC.n2724 VCC.n2255 0.0174643
R49328 VCC.n2724 VCC.n2723 0.0174643
R49329 VCC.n2716 VCC.n2256 0.0174643
R49330 VCC.n2722 VCC.n2256 0.0174643
R49331 VCC.n2594 VCC.n2317 0.0174643
R49332 VCC.n2595 VCC.n2594 0.0174643
R49333 VCC.n2599 VCC.n2319 0.0174643
R49334 VCC.n2596 VCC.n2319 0.0174643
R49335 VCC.n2472 VCC.n2376 0.0174643
R49336 VCC.n2471 VCC.n2382 0.0174643
R49337 VCC.n3023 VCC.n2927 0.0174643
R49338 VCC.n3022 VCC.n2933 0.0174643
R49339 VCC.n3146 VCC.n2869 0.0174643
R49340 VCC.n3147 VCC.n3146 0.0174643
R49341 VCC.n3151 VCC.n2871 0.0174643
R49342 VCC.n3148 VCC.n2871 0.0174643
R49343 VCC.n3271 VCC.n3270 0.0174643
R49344 VCC.n3270 VCC.n2802 0.0174643
R49345 VCC.n3272 VCC.n2807 0.0174643
R49346 VCC.n2807 VCC.n2803 0.0174643
R49347 VCC.n3833 VCC.n3364 0.0174643
R49348 VCC.n3833 VCC.n3832 0.0174643
R49349 VCC.n3825 VCC.n3365 0.0174643
R49350 VCC.n3831 VCC.n3365 0.0174643
R49351 VCC.n3703 VCC.n3426 0.0174643
R49352 VCC.n3704 VCC.n3703 0.0174643
R49353 VCC.n3708 VCC.n3428 0.0174643
R49354 VCC.n3705 VCC.n3428 0.0174643
R49355 VCC.n3581 VCC.n3485 0.0174643
R49356 VCC.n3580 VCC.n3491 0.0174643
R49357 VCC.n4132 VCC.n4036 0.0174643
R49358 VCC.n4131 VCC.n4042 0.0174643
R49359 VCC.n4255 VCC.n3978 0.0174643
R49360 VCC.n4256 VCC.n4255 0.0174643
R49361 VCC.n4260 VCC.n3980 0.0174643
R49362 VCC.n4257 VCC.n3980 0.0174643
R49363 VCC.n4380 VCC.n4379 0.0174643
R49364 VCC.n4379 VCC.n3911 0.0174643
R49365 VCC.n4381 VCC.n3916 0.0174643
R49366 VCC.n3916 VCC.n3912 0.0174643
R49367 VCC.n4942 VCC.n4473 0.0174643
R49368 VCC.n4942 VCC.n4941 0.0174643
R49369 VCC.n4934 VCC.n4474 0.0174643
R49370 VCC.n4940 VCC.n4474 0.0174643
R49371 VCC.n4812 VCC.n4535 0.0174643
R49372 VCC.n4813 VCC.n4812 0.0174643
R49373 VCC.n4817 VCC.n4537 0.0174643
R49374 VCC.n4814 VCC.n4537 0.0174643
R49375 VCC.n4690 VCC.n4594 0.0174643
R49376 VCC.n4689 VCC.n4600 0.0174643
R49377 VCC.n5241 VCC.n5145 0.0174643
R49378 VCC.n5240 VCC.n5151 0.0174643
R49379 VCC.n5364 VCC.n5087 0.0174643
R49380 VCC.n5365 VCC.n5364 0.0174643
R49381 VCC.n5369 VCC.n5089 0.0174643
R49382 VCC.n5366 VCC.n5089 0.0174643
R49383 VCC.n5489 VCC.n5488 0.0174643
R49384 VCC.n5488 VCC.n5020 0.0174643
R49385 VCC.n5490 VCC.n5025 0.0174643
R49386 VCC.n5025 VCC.n5021 0.0174643
R49387 VCC.n6051 VCC.n5582 0.0174643
R49388 VCC.n6051 VCC.n6050 0.0174643
R49389 VCC.n6043 VCC.n5583 0.0174643
R49390 VCC.n6049 VCC.n5583 0.0174643
R49391 VCC.n5921 VCC.n5644 0.0174643
R49392 VCC.n5922 VCC.n5921 0.0174643
R49393 VCC.n5926 VCC.n5646 0.0174643
R49394 VCC.n5923 VCC.n5646 0.0174643
R49395 VCC.n5799 VCC.n5703 0.0174643
R49396 VCC.n5798 VCC.n5709 0.0174643
R49397 VCC.n6350 VCC.n6254 0.0174643
R49398 VCC.n6349 VCC.n6260 0.0174643
R49399 VCC.n6473 VCC.n6196 0.0174643
R49400 VCC.n6474 VCC.n6473 0.0174643
R49401 VCC.n6478 VCC.n6198 0.0174643
R49402 VCC.n6475 VCC.n6198 0.0174643
R49403 VCC.n6598 VCC.n6597 0.0174643
R49404 VCC.n6597 VCC.n6129 0.0174643
R49405 VCC.n6599 VCC.n6134 0.0174643
R49406 VCC.n6134 VCC.n6130 0.0174643
R49407 VCC.n7160 VCC.n6691 0.0174643
R49408 VCC.n7160 VCC.n7159 0.0174643
R49409 VCC.n7152 VCC.n6692 0.0174643
R49410 VCC.n7158 VCC.n6692 0.0174643
R49411 VCC.n7030 VCC.n6753 0.0174643
R49412 VCC.n7031 VCC.n7030 0.0174643
R49413 VCC.n7035 VCC.n6755 0.0174643
R49414 VCC.n7032 VCC.n6755 0.0174643
R49415 VCC.n6908 VCC.n6812 0.0174643
R49416 VCC.n6907 VCC.n6818 0.0174643
R49417 VCC.n7459 VCC.n7363 0.0174643
R49418 VCC.n7458 VCC.n7369 0.0174643
R49419 VCC.n7582 VCC.n7305 0.0174643
R49420 VCC.n7583 VCC.n7582 0.0174643
R49421 VCC.n7587 VCC.n7307 0.0174643
R49422 VCC.n7584 VCC.n7307 0.0174643
R49423 VCC.n7707 VCC.n7706 0.0174643
R49424 VCC.n7706 VCC.n7238 0.0174643
R49425 VCC.n7708 VCC.n7243 0.0174643
R49426 VCC.n7243 VCC.n7239 0.0174643
R49427 VCC.n8269 VCC.n7800 0.0174643
R49428 VCC.n8269 VCC.n8268 0.0174643
R49429 VCC.n8261 VCC.n7801 0.0174643
R49430 VCC.n8267 VCC.n7801 0.0174643
R49431 VCC.n8139 VCC.n7862 0.0174643
R49432 VCC.n8140 VCC.n8139 0.0174643
R49433 VCC.n8144 VCC.n7864 0.0174643
R49434 VCC.n8141 VCC.n7864 0.0174643
R49435 VCC.n8017 VCC.n7921 0.0174643
R49436 VCC.n8016 VCC.n7927 0.0174643
R49437 VCC.n8691 VCC.n8414 0.0174643
R49438 VCC.n8692 VCC.n8691 0.0174643
R49439 VCC.n8696 VCC.n8416 0.0174643
R49440 VCC.n8693 VCC.n8416 0.0174643
R49441 VCC.n8816 VCC.n8815 0.0174643
R49442 VCC.n8815 VCC.n8347 0.0174643
R49443 VCC.n8817 VCC.n8352 0.0174643
R49444 VCC.n8352 VCC.n8348 0.0174643
R49445 VCC.n8568 VCC.n8472 0.0174643
R49446 VCC.n8567 VCC.n8478 0.0174643
R49447 VCC.n9378 VCC.n8909 0.0174643
R49448 VCC.n9378 VCC.n9377 0.0174643
R49449 VCC.n9370 VCC.n8910 0.0174643
R49450 VCC.n9376 VCC.n8910 0.0174643
R49451 VCC.n9248 VCC.n8971 0.0174643
R49452 VCC.n9249 VCC.n9248 0.0174643
R49453 VCC.n9253 VCC.n8973 0.0174643
R49454 VCC.n9250 VCC.n8973 0.0174643
R49455 VCC.n9126 VCC.n9030 0.0174643
R49456 VCC.n9125 VCC.n9036 0.0174643
R49457 VCC.n9677 VCC.n9581 0.0174643
R49458 VCC.n9676 VCC.n9587 0.0174643
R49459 VCC.n9800 VCC.n9523 0.0174643
R49460 VCC.n9801 VCC.n9800 0.0174643
R49461 VCC.n9805 VCC.n9525 0.0174643
R49462 VCC.n9802 VCC.n9525 0.0174643
R49463 VCC.n9925 VCC.n9924 0.0174643
R49464 VCC.n9924 VCC.n9456 0.0174643
R49465 VCC.n9926 VCC.n9461 0.0174643
R49466 VCC.n9461 VCC.n9457 0.0174643
R49467 VCC.n10486 VCC.n10017 0.0174643
R49468 VCC.n10486 VCC.n10485 0.0174643
R49469 VCC.n10478 VCC.n10018 0.0174643
R49470 VCC.n10484 VCC.n10018 0.0174643
R49471 VCC.n10356 VCC.n10079 0.0174643
R49472 VCC.n10357 VCC.n10356 0.0174643
R49473 VCC.n10361 VCC.n10081 0.0174643
R49474 VCC.n10358 VCC.n10081 0.0174643
R49475 VCC.n10234 VCC.n10138 0.0174643
R49476 VCC.n10233 VCC.n10144 0.0174643
R49477 VCC.n10784 VCC.n10688 0.0174643
R49478 VCC.n10783 VCC.n10694 0.0174643
R49479 VCC.n10907 VCC.n10630 0.0174643
R49480 VCC.n10908 VCC.n10907 0.0174643
R49481 VCC.n10912 VCC.n10632 0.0174643
R49482 VCC.n10909 VCC.n10632 0.0174643
R49483 VCC.n11032 VCC.n11031 0.0174643
R49484 VCC.n11031 VCC.n10563 0.0174643
R49485 VCC.n11033 VCC.n10568 0.0174643
R49486 VCC.n10568 VCC.n10564 0.0174643
R49487 VCC.n11593 VCC.n11124 0.0174643
R49488 VCC.n11593 VCC.n11592 0.0174643
R49489 VCC.n11585 VCC.n11125 0.0174643
R49490 VCC.n11591 VCC.n11125 0.0174643
R49491 VCC.n11463 VCC.n11186 0.0174643
R49492 VCC.n11464 VCC.n11463 0.0174643
R49493 VCC.n11468 VCC.n11188 0.0174643
R49494 VCC.n11465 VCC.n11188 0.0174643
R49495 VCC.n11341 VCC.n11245 0.0174643
R49496 VCC.n11340 VCC.n11251 0.0174643
R49497 VCC.n11891 VCC.n11795 0.0174643
R49498 VCC.n11890 VCC.n11801 0.0174643
R49499 VCC.n12014 VCC.n11737 0.0174643
R49500 VCC.n12015 VCC.n12014 0.0174643
R49501 VCC.n12019 VCC.n11739 0.0174643
R49502 VCC.n12016 VCC.n11739 0.0174643
R49503 VCC.n12139 VCC.n12138 0.0174643
R49504 VCC.n12138 VCC.n11670 0.0174643
R49505 VCC.n12140 VCC.n11675 0.0174643
R49506 VCC.n11675 VCC.n11671 0.0174643
R49507 VCC.n12700 VCC.n12231 0.0174643
R49508 VCC.n12700 VCC.n12699 0.0174643
R49509 VCC.n12692 VCC.n12232 0.0174643
R49510 VCC.n12698 VCC.n12232 0.0174643
R49511 VCC.n12570 VCC.n12293 0.0174643
R49512 VCC.n12571 VCC.n12570 0.0174643
R49513 VCC.n12575 VCC.n12295 0.0174643
R49514 VCC.n12572 VCC.n12295 0.0174643
R49515 VCC.n12448 VCC.n12352 0.0174643
R49516 VCC.n12447 VCC.n12358 0.0174643
R49517 VCC.n12998 VCC.n12902 0.0174643
R49518 VCC.n12997 VCC.n12908 0.0174643
R49519 VCC.n13121 VCC.n12844 0.0174643
R49520 VCC.n13122 VCC.n13121 0.0174643
R49521 VCC.n13126 VCC.n12846 0.0174643
R49522 VCC.n13123 VCC.n12846 0.0174643
R49523 VCC.n13246 VCC.n13245 0.0174643
R49524 VCC.n13245 VCC.n12777 0.0174643
R49525 VCC.n13247 VCC.n12782 0.0174643
R49526 VCC.n12782 VCC.n12778 0.0174643
R49527 VCC.n13807 VCC.n13338 0.0174643
R49528 VCC.n13807 VCC.n13806 0.0174643
R49529 VCC.n13799 VCC.n13339 0.0174643
R49530 VCC.n13805 VCC.n13339 0.0174643
R49531 VCC.n13677 VCC.n13400 0.0174643
R49532 VCC.n13678 VCC.n13677 0.0174643
R49533 VCC.n13682 VCC.n13402 0.0174643
R49534 VCC.n13679 VCC.n13402 0.0174643
R49535 VCC.n13555 VCC.n13459 0.0174643
R49536 VCC.n13554 VCC.n13465 0.0174643
R49537 VCC.n14105 VCC.n14009 0.0174643
R49538 VCC.n14104 VCC.n14015 0.0174643
R49539 VCC.n14228 VCC.n13951 0.0174643
R49540 VCC.n14229 VCC.n14228 0.0174643
R49541 VCC.n14233 VCC.n13953 0.0174643
R49542 VCC.n14230 VCC.n13953 0.0174643
R49543 VCC.n14353 VCC.n14352 0.0174643
R49544 VCC.n14352 VCC.n13884 0.0174643
R49545 VCC.n14354 VCC.n13889 0.0174643
R49546 VCC.n13889 VCC.n13885 0.0174643
R49547 VCC.n14914 VCC.n14445 0.0174643
R49548 VCC.n14914 VCC.n14913 0.0174643
R49549 VCC.n14906 VCC.n14446 0.0174643
R49550 VCC.n14912 VCC.n14446 0.0174643
R49551 VCC.n14784 VCC.n14507 0.0174643
R49552 VCC.n14785 VCC.n14784 0.0174643
R49553 VCC.n14789 VCC.n14509 0.0174643
R49554 VCC.n14786 VCC.n14509 0.0174643
R49555 VCC.n14662 VCC.n14566 0.0174643
R49556 VCC.n14661 VCC.n14572 0.0174643
R49557 VCC.n15212 VCC.n15116 0.0174643
R49558 VCC.n15211 VCC.n15122 0.0174643
R49559 VCC.n15335 VCC.n15058 0.0174643
R49560 VCC.n15336 VCC.n15335 0.0174643
R49561 VCC.n15340 VCC.n15060 0.0174643
R49562 VCC.n15337 VCC.n15060 0.0174643
R49563 VCC.n15460 VCC.n15459 0.0174643
R49564 VCC.n15459 VCC.n14991 0.0174643
R49565 VCC.n15461 VCC.n14996 0.0174643
R49566 VCC.n14996 VCC.n14992 0.0174643
R49567 VCC.n16021 VCC.n15552 0.0174643
R49568 VCC.n16021 VCC.n16020 0.0174643
R49569 VCC.n16013 VCC.n15553 0.0174643
R49570 VCC.n16019 VCC.n15553 0.0174643
R49571 VCC.n15891 VCC.n15614 0.0174643
R49572 VCC.n15892 VCC.n15891 0.0174643
R49573 VCC.n15896 VCC.n15616 0.0174643
R49574 VCC.n15893 VCC.n15616 0.0174643
R49575 VCC.n15769 VCC.n15673 0.0174643
R49576 VCC.n15768 VCC.n15679 0.0174643
R49577 VCC.n16319 VCC.n16223 0.0174643
R49578 VCC.n16318 VCC.n16229 0.0174643
R49579 VCC.n16442 VCC.n16165 0.0174643
R49580 VCC.n16443 VCC.n16442 0.0174643
R49581 VCC.n16447 VCC.n16167 0.0174643
R49582 VCC.n16444 VCC.n16167 0.0174643
R49583 VCC.n16567 VCC.n16566 0.0174643
R49584 VCC.n16566 VCC.n16098 0.0174643
R49585 VCC.n16568 VCC.n16103 0.0174643
R49586 VCC.n16103 VCC.n16099 0.0174643
R49587 VCC.n17128 VCC.n16659 0.0174643
R49588 VCC.n17128 VCC.n17127 0.0174643
R49589 VCC.n17120 VCC.n16660 0.0174643
R49590 VCC.n17126 VCC.n16660 0.0174643
R49591 VCC.n16998 VCC.n16721 0.0174643
R49592 VCC.n16999 VCC.n16998 0.0174643
R49593 VCC.n17003 VCC.n16723 0.0174643
R49594 VCC.n17000 VCC.n16723 0.0174643
R49595 VCC.n16876 VCC.n16780 0.0174643
R49596 VCC.n16875 VCC.n16786 0.0174643
R49597 VCC.n17362 VCC.n17272 0.0174643
R49598 VCC.n17363 VCC.n17362 0.0174643
R49599 VCC.n17367 VCC.n17274 0.0174643
R49600 VCC.n17364 VCC.n17274 0.0174643
R49601 VCC.n17487 VCC.n17486 0.0174643
R49602 VCC.n17486 VCC.n17205 0.0174643
R49603 VCC.n17488 VCC.n17210 0.0174643
R49604 VCC.n17210 VCC.n17206 0.0174643
R49605 VCC.n238 VCC.n233 0.0165714
R49606 VCC.n255 VCC.n254 0.0165714
R49607 VCC.n204 VCC.n197 0.0165714
R49608 VCC.n240 VCC.n239 0.0165714
R49609 VCC.n256 VCC.n167 0.0165714
R49610 VCC.n282 VCC.n146 0.0165714
R49611 VCC.n301 VCC.n300 0.0165714
R49612 VCC.n401 VCC.n400 0.0165714
R49613 VCC.n329 VCC.n321 0.0165714
R49614 VCC.n354 VCC.n348 0.0165714
R49615 VCC.n409 VCC.n86 0.0165714
R49616 VCC.n436 VCC.n435 0.0165714
R49617 VCC.n454 VCC.n60 0.0165714
R49618 VCC.n514 VCC.n29 0.0165714
R49619 VCC.n541 VCC.n10 0.0165714
R49620 VCC.n790 VCC.n785 0.0165714
R49621 VCC.n807 VCC.n806 0.0165714
R49622 VCC.n756 VCC.n749 0.0165714
R49623 VCC.n792 VCC.n791 0.0165714
R49624 VCC.n808 VCC.n719 0.0165714
R49625 VCC.n834 VCC.n698 0.0165714
R49626 VCC.n853 VCC.n852 0.0165714
R49627 VCC.n953 VCC.n952 0.0165714
R49628 VCC.n881 VCC.n873 0.0165714
R49629 VCC.n906 VCC.n900 0.0165714
R49630 VCC.n961 VCC.n638 0.0165714
R49631 VCC.n988 VCC.n987 0.0165714
R49632 VCC.n1006 VCC.n612 0.0165714
R49633 VCC.n1066 VCC.n581 0.0165714
R49634 VCC.n1095 VCC.n564 0.0165714
R49635 VCC.n1565 VCC.n1564 0.0165714
R49636 VCC.n1631 VCC.n1630 0.0165714
R49637 VCC.n1644 VCC.n1643 0.0165714
R49638 VCC.n1510 VCC.n1509 0.0165714
R49639 VCC.n1438 VCC.n1429 0.0165714
R49640 VCC.n1463 VCC.n1457 0.0165714
R49641 VCC.n1518 VCC.n1195 0.0165714
R49642 VCC.n1546 VCC.n1545 0.0165714
R49643 VCC.n1348 VCC.n1343 0.0165714
R49644 VCC.n1365 VCC.n1364 0.0165714
R49645 VCC.n1314 VCC.n1307 0.0165714
R49646 VCC.n1350 VCC.n1349 0.0165714
R49647 VCC.n1366 VCC.n1277 0.0165714
R49648 VCC.n1392 VCC.n1256 0.0165714
R49649 VCC.n1411 VCC.n1410 0.0165714
R49650 VCC.n1899 VCC.n1894 0.0165714
R49651 VCC.n1916 VCC.n1915 0.0165714
R49652 VCC.n1865 VCC.n1858 0.0165714
R49653 VCC.n1901 VCC.n1900 0.0165714
R49654 VCC.n1917 VCC.n1828 0.0165714
R49655 VCC.n1943 VCC.n1807 0.0165714
R49656 VCC.n1962 VCC.n1961 0.0165714
R49657 VCC.n2062 VCC.n2061 0.0165714
R49658 VCC.n1990 VCC.n1982 0.0165714
R49659 VCC.n2015 VCC.n2009 0.0165714
R49660 VCC.n2070 VCC.n1747 0.0165714
R49661 VCC.n2097 VCC.n2096 0.0165714
R49662 VCC.n2115 VCC.n1721 0.0165714
R49663 VCC.n2175 VCC.n1690 0.0165714
R49664 VCC.n2204 VCC.n1673 0.0165714
R49665 VCC.n2674 VCC.n2673 0.0165714
R49666 VCC.n2740 VCC.n2739 0.0165714
R49667 VCC.n2753 VCC.n2752 0.0165714
R49668 VCC.n2619 VCC.n2618 0.0165714
R49669 VCC.n2547 VCC.n2538 0.0165714
R49670 VCC.n2572 VCC.n2566 0.0165714
R49671 VCC.n2627 VCC.n2304 0.0165714
R49672 VCC.n2655 VCC.n2654 0.0165714
R49673 VCC.n2457 VCC.n2452 0.0165714
R49674 VCC.n2474 VCC.n2473 0.0165714
R49675 VCC.n2423 VCC.n2416 0.0165714
R49676 VCC.n2459 VCC.n2458 0.0165714
R49677 VCC.n2475 VCC.n2386 0.0165714
R49678 VCC.n2501 VCC.n2365 0.0165714
R49679 VCC.n2520 VCC.n2519 0.0165714
R49680 VCC.n3008 VCC.n3003 0.0165714
R49681 VCC.n3025 VCC.n3024 0.0165714
R49682 VCC.n2974 VCC.n2967 0.0165714
R49683 VCC.n3010 VCC.n3009 0.0165714
R49684 VCC.n3026 VCC.n2937 0.0165714
R49685 VCC.n3052 VCC.n2916 0.0165714
R49686 VCC.n3071 VCC.n3070 0.0165714
R49687 VCC.n3171 VCC.n3170 0.0165714
R49688 VCC.n3099 VCC.n3091 0.0165714
R49689 VCC.n3124 VCC.n3118 0.0165714
R49690 VCC.n3179 VCC.n2856 0.0165714
R49691 VCC.n3206 VCC.n3205 0.0165714
R49692 VCC.n3224 VCC.n2830 0.0165714
R49693 VCC.n3284 VCC.n2799 0.0165714
R49694 VCC.n3313 VCC.n2782 0.0165714
R49695 VCC.n3783 VCC.n3782 0.0165714
R49696 VCC.n3849 VCC.n3848 0.0165714
R49697 VCC.n3862 VCC.n3861 0.0165714
R49698 VCC.n3728 VCC.n3727 0.0165714
R49699 VCC.n3656 VCC.n3647 0.0165714
R49700 VCC.n3681 VCC.n3675 0.0165714
R49701 VCC.n3736 VCC.n3413 0.0165714
R49702 VCC.n3764 VCC.n3763 0.0165714
R49703 VCC.n3566 VCC.n3561 0.0165714
R49704 VCC.n3583 VCC.n3582 0.0165714
R49705 VCC.n3532 VCC.n3525 0.0165714
R49706 VCC.n3568 VCC.n3567 0.0165714
R49707 VCC.n3584 VCC.n3495 0.0165714
R49708 VCC.n3610 VCC.n3474 0.0165714
R49709 VCC.n3629 VCC.n3628 0.0165714
R49710 VCC.n4117 VCC.n4112 0.0165714
R49711 VCC.n4134 VCC.n4133 0.0165714
R49712 VCC.n4083 VCC.n4076 0.0165714
R49713 VCC.n4119 VCC.n4118 0.0165714
R49714 VCC.n4135 VCC.n4046 0.0165714
R49715 VCC.n4161 VCC.n4025 0.0165714
R49716 VCC.n4180 VCC.n4179 0.0165714
R49717 VCC.n4280 VCC.n4279 0.0165714
R49718 VCC.n4208 VCC.n4200 0.0165714
R49719 VCC.n4233 VCC.n4227 0.0165714
R49720 VCC.n4288 VCC.n3965 0.0165714
R49721 VCC.n4315 VCC.n4314 0.0165714
R49722 VCC.n4333 VCC.n3939 0.0165714
R49723 VCC.n4393 VCC.n3908 0.0165714
R49724 VCC.n4422 VCC.n3891 0.0165714
R49725 VCC.n4892 VCC.n4891 0.0165714
R49726 VCC.n4958 VCC.n4957 0.0165714
R49727 VCC.n4971 VCC.n4970 0.0165714
R49728 VCC.n4837 VCC.n4836 0.0165714
R49729 VCC.n4765 VCC.n4756 0.0165714
R49730 VCC.n4790 VCC.n4784 0.0165714
R49731 VCC.n4845 VCC.n4522 0.0165714
R49732 VCC.n4873 VCC.n4872 0.0165714
R49733 VCC.n4675 VCC.n4670 0.0165714
R49734 VCC.n4692 VCC.n4691 0.0165714
R49735 VCC.n4641 VCC.n4634 0.0165714
R49736 VCC.n4677 VCC.n4676 0.0165714
R49737 VCC.n4693 VCC.n4604 0.0165714
R49738 VCC.n4719 VCC.n4583 0.0165714
R49739 VCC.n4738 VCC.n4737 0.0165714
R49740 VCC.n5226 VCC.n5221 0.0165714
R49741 VCC.n5243 VCC.n5242 0.0165714
R49742 VCC.n5192 VCC.n5185 0.0165714
R49743 VCC.n5228 VCC.n5227 0.0165714
R49744 VCC.n5244 VCC.n5155 0.0165714
R49745 VCC.n5270 VCC.n5134 0.0165714
R49746 VCC.n5289 VCC.n5288 0.0165714
R49747 VCC.n5389 VCC.n5388 0.0165714
R49748 VCC.n5317 VCC.n5309 0.0165714
R49749 VCC.n5342 VCC.n5336 0.0165714
R49750 VCC.n5397 VCC.n5074 0.0165714
R49751 VCC.n5424 VCC.n5423 0.0165714
R49752 VCC.n5442 VCC.n5048 0.0165714
R49753 VCC.n5502 VCC.n5017 0.0165714
R49754 VCC.n5531 VCC.n5000 0.0165714
R49755 VCC.n6001 VCC.n6000 0.0165714
R49756 VCC.n6067 VCC.n6066 0.0165714
R49757 VCC.n6080 VCC.n6079 0.0165714
R49758 VCC.n5946 VCC.n5945 0.0165714
R49759 VCC.n5874 VCC.n5865 0.0165714
R49760 VCC.n5899 VCC.n5893 0.0165714
R49761 VCC.n5954 VCC.n5631 0.0165714
R49762 VCC.n5982 VCC.n5981 0.0165714
R49763 VCC.n5784 VCC.n5779 0.0165714
R49764 VCC.n5801 VCC.n5800 0.0165714
R49765 VCC.n5750 VCC.n5743 0.0165714
R49766 VCC.n5786 VCC.n5785 0.0165714
R49767 VCC.n5802 VCC.n5713 0.0165714
R49768 VCC.n5828 VCC.n5692 0.0165714
R49769 VCC.n5847 VCC.n5846 0.0165714
R49770 VCC.n6335 VCC.n6330 0.0165714
R49771 VCC.n6352 VCC.n6351 0.0165714
R49772 VCC.n6301 VCC.n6294 0.0165714
R49773 VCC.n6337 VCC.n6336 0.0165714
R49774 VCC.n6353 VCC.n6264 0.0165714
R49775 VCC.n6379 VCC.n6243 0.0165714
R49776 VCC.n6398 VCC.n6397 0.0165714
R49777 VCC.n6498 VCC.n6497 0.0165714
R49778 VCC.n6426 VCC.n6418 0.0165714
R49779 VCC.n6451 VCC.n6445 0.0165714
R49780 VCC.n6506 VCC.n6183 0.0165714
R49781 VCC.n6533 VCC.n6532 0.0165714
R49782 VCC.n6551 VCC.n6157 0.0165714
R49783 VCC.n6611 VCC.n6126 0.0165714
R49784 VCC.n6640 VCC.n6109 0.0165714
R49785 VCC.n7110 VCC.n7109 0.0165714
R49786 VCC.n7176 VCC.n7175 0.0165714
R49787 VCC.n7189 VCC.n7188 0.0165714
R49788 VCC.n7055 VCC.n7054 0.0165714
R49789 VCC.n6983 VCC.n6974 0.0165714
R49790 VCC.n7008 VCC.n7002 0.0165714
R49791 VCC.n7063 VCC.n6740 0.0165714
R49792 VCC.n7091 VCC.n7090 0.0165714
R49793 VCC.n6893 VCC.n6888 0.0165714
R49794 VCC.n6910 VCC.n6909 0.0165714
R49795 VCC.n6859 VCC.n6852 0.0165714
R49796 VCC.n6895 VCC.n6894 0.0165714
R49797 VCC.n6911 VCC.n6822 0.0165714
R49798 VCC.n6937 VCC.n6801 0.0165714
R49799 VCC.n6956 VCC.n6955 0.0165714
R49800 VCC.n7444 VCC.n7439 0.0165714
R49801 VCC.n7461 VCC.n7460 0.0165714
R49802 VCC.n7410 VCC.n7403 0.0165714
R49803 VCC.n7446 VCC.n7445 0.0165714
R49804 VCC.n7462 VCC.n7373 0.0165714
R49805 VCC.n7488 VCC.n7352 0.0165714
R49806 VCC.n7507 VCC.n7506 0.0165714
R49807 VCC.n7607 VCC.n7606 0.0165714
R49808 VCC.n7535 VCC.n7527 0.0165714
R49809 VCC.n7560 VCC.n7554 0.0165714
R49810 VCC.n7615 VCC.n7292 0.0165714
R49811 VCC.n7642 VCC.n7641 0.0165714
R49812 VCC.n7660 VCC.n7266 0.0165714
R49813 VCC.n7720 VCC.n7235 0.0165714
R49814 VCC.n7749 VCC.n7218 0.0165714
R49815 VCC.n8219 VCC.n8218 0.0165714
R49816 VCC.n8285 VCC.n8284 0.0165714
R49817 VCC.n8298 VCC.n8297 0.0165714
R49818 VCC.n8164 VCC.n8163 0.0165714
R49819 VCC.n8092 VCC.n8083 0.0165714
R49820 VCC.n8117 VCC.n8111 0.0165714
R49821 VCC.n8172 VCC.n7849 0.0165714
R49822 VCC.n8200 VCC.n8199 0.0165714
R49823 VCC.n8002 VCC.n7997 0.0165714
R49824 VCC.n8019 VCC.n8018 0.0165714
R49825 VCC.n7968 VCC.n7961 0.0165714
R49826 VCC.n8004 VCC.n8003 0.0165714
R49827 VCC.n8020 VCC.n7931 0.0165714
R49828 VCC.n8046 VCC.n7910 0.0165714
R49829 VCC.n8065 VCC.n8064 0.0165714
R49830 VCC.n8716 VCC.n8715 0.0165714
R49831 VCC.n8644 VCC.n8636 0.0165714
R49832 VCC.n8669 VCC.n8663 0.0165714
R49833 VCC.n8724 VCC.n8401 0.0165714
R49834 VCC.n8751 VCC.n8750 0.0165714
R49835 VCC.n8769 VCC.n8375 0.0165714
R49836 VCC.n8829 VCC.n8344 0.0165714
R49837 VCC.n8858 VCC.n8327 0.0165714
R49838 VCC.n8553 VCC.n8548 0.0165714
R49839 VCC.n8570 VCC.n8569 0.0165714
R49840 VCC.n8519 VCC.n8512 0.0165714
R49841 VCC.n8555 VCC.n8554 0.0165714
R49842 VCC.n8571 VCC.n8482 0.0165714
R49843 VCC.n8597 VCC.n8461 0.0165714
R49844 VCC.n8616 VCC.n8615 0.0165714
R49845 VCC.n9328 VCC.n9327 0.0165714
R49846 VCC.n9394 VCC.n9393 0.0165714
R49847 VCC.n9407 VCC.n9406 0.0165714
R49848 VCC.n9273 VCC.n9272 0.0165714
R49849 VCC.n9201 VCC.n9192 0.0165714
R49850 VCC.n9226 VCC.n9220 0.0165714
R49851 VCC.n9281 VCC.n8958 0.0165714
R49852 VCC.n9309 VCC.n9308 0.0165714
R49853 VCC.n9111 VCC.n9106 0.0165714
R49854 VCC.n9128 VCC.n9127 0.0165714
R49855 VCC.n9077 VCC.n9070 0.0165714
R49856 VCC.n9113 VCC.n9112 0.0165714
R49857 VCC.n9129 VCC.n9040 0.0165714
R49858 VCC.n9155 VCC.n9019 0.0165714
R49859 VCC.n9174 VCC.n9173 0.0165714
R49860 VCC.n9662 VCC.n9657 0.0165714
R49861 VCC.n9679 VCC.n9678 0.0165714
R49862 VCC.n9628 VCC.n9621 0.0165714
R49863 VCC.n9664 VCC.n9663 0.0165714
R49864 VCC.n9680 VCC.n9591 0.0165714
R49865 VCC.n9706 VCC.n9570 0.0165714
R49866 VCC.n9725 VCC.n9724 0.0165714
R49867 VCC.n9825 VCC.n9824 0.0165714
R49868 VCC.n9753 VCC.n9745 0.0165714
R49869 VCC.n9778 VCC.n9772 0.0165714
R49870 VCC.n9833 VCC.n9510 0.0165714
R49871 VCC.n9860 VCC.n9859 0.0165714
R49872 VCC.n9878 VCC.n9484 0.0165714
R49873 VCC.n9938 VCC.n9453 0.0165714
R49874 VCC.n9967 VCC.n9436 0.0165714
R49875 VCC.n10436 VCC.n10435 0.0165714
R49876 VCC.n10502 VCC.n10501 0.0165714
R49877 VCC.n10515 VCC.n10514 0.0165714
R49878 VCC.n10381 VCC.n10380 0.0165714
R49879 VCC.n10309 VCC.n10300 0.0165714
R49880 VCC.n10334 VCC.n10328 0.0165714
R49881 VCC.n10389 VCC.n10066 0.0165714
R49882 VCC.n10417 VCC.n10416 0.0165714
R49883 VCC.n10219 VCC.n10214 0.0165714
R49884 VCC.n10236 VCC.n10235 0.0165714
R49885 VCC.n10185 VCC.n10178 0.0165714
R49886 VCC.n10221 VCC.n10220 0.0165714
R49887 VCC.n10237 VCC.n10148 0.0165714
R49888 VCC.n10263 VCC.n10127 0.0165714
R49889 VCC.n10282 VCC.n10281 0.0165714
R49890 VCC.n10769 VCC.n10764 0.0165714
R49891 VCC.n10786 VCC.n10785 0.0165714
R49892 VCC.n10735 VCC.n10728 0.0165714
R49893 VCC.n10771 VCC.n10770 0.0165714
R49894 VCC.n10787 VCC.n10698 0.0165714
R49895 VCC.n10813 VCC.n10677 0.0165714
R49896 VCC.n10832 VCC.n10831 0.0165714
R49897 VCC.n10932 VCC.n10931 0.0165714
R49898 VCC.n10860 VCC.n10852 0.0165714
R49899 VCC.n10885 VCC.n10879 0.0165714
R49900 VCC.n10940 VCC.n10617 0.0165714
R49901 VCC.n10967 VCC.n10966 0.0165714
R49902 VCC.n10985 VCC.n10591 0.0165714
R49903 VCC.n11045 VCC.n10560 0.0165714
R49904 VCC.n11074 VCC.n10543 0.0165714
R49905 VCC.n11543 VCC.n11542 0.0165714
R49906 VCC.n11609 VCC.n11608 0.0165714
R49907 VCC.n11622 VCC.n11621 0.0165714
R49908 VCC.n11488 VCC.n11487 0.0165714
R49909 VCC.n11416 VCC.n11407 0.0165714
R49910 VCC.n11441 VCC.n11435 0.0165714
R49911 VCC.n11496 VCC.n11173 0.0165714
R49912 VCC.n11524 VCC.n11523 0.0165714
R49913 VCC.n11326 VCC.n11321 0.0165714
R49914 VCC.n11343 VCC.n11342 0.0165714
R49915 VCC.n11292 VCC.n11285 0.0165714
R49916 VCC.n11328 VCC.n11327 0.0165714
R49917 VCC.n11344 VCC.n11255 0.0165714
R49918 VCC.n11370 VCC.n11234 0.0165714
R49919 VCC.n11389 VCC.n11388 0.0165714
R49920 VCC.n11876 VCC.n11871 0.0165714
R49921 VCC.n11893 VCC.n11892 0.0165714
R49922 VCC.n11842 VCC.n11835 0.0165714
R49923 VCC.n11878 VCC.n11877 0.0165714
R49924 VCC.n11894 VCC.n11805 0.0165714
R49925 VCC.n11920 VCC.n11784 0.0165714
R49926 VCC.n11939 VCC.n11938 0.0165714
R49927 VCC.n12039 VCC.n12038 0.0165714
R49928 VCC.n11967 VCC.n11959 0.0165714
R49929 VCC.n11992 VCC.n11986 0.0165714
R49930 VCC.n12047 VCC.n11724 0.0165714
R49931 VCC.n12074 VCC.n12073 0.0165714
R49932 VCC.n12092 VCC.n11698 0.0165714
R49933 VCC.n12152 VCC.n11667 0.0165714
R49934 VCC.n12181 VCC.n11650 0.0165714
R49935 VCC.n12650 VCC.n12649 0.0165714
R49936 VCC.n12716 VCC.n12715 0.0165714
R49937 VCC.n12729 VCC.n12728 0.0165714
R49938 VCC.n12595 VCC.n12594 0.0165714
R49939 VCC.n12523 VCC.n12514 0.0165714
R49940 VCC.n12548 VCC.n12542 0.0165714
R49941 VCC.n12603 VCC.n12280 0.0165714
R49942 VCC.n12631 VCC.n12630 0.0165714
R49943 VCC.n12433 VCC.n12428 0.0165714
R49944 VCC.n12450 VCC.n12449 0.0165714
R49945 VCC.n12399 VCC.n12392 0.0165714
R49946 VCC.n12435 VCC.n12434 0.0165714
R49947 VCC.n12451 VCC.n12362 0.0165714
R49948 VCC.n12477 VCC.n12341 0.0165714
R49949 VCC.n12496 VCC.n12495 0.0165714
R49950 VCC.n12983 VCC.n12978 0.0165714
R49951 VCC.n13000 VCC.n12999 0.0165714
R49952 VCC.n12949 VCC.n12942 0.0165714
R49953 VCC.n12985 VCC.n12984 0.0165714
R49954 VCC.n13001 VCC.n12912 0.0165714
R49955 VCC.n13027 VCC.n12891 0.0165714
R49956 VCC.n13046 VCC.n13045 0.0165714
R49957 VCC.n13146 VCC.n13145 0.0165714
R49958 VCC.n13074 VCC.n13066 0.0165714
R49959 VCC.n13099 VCC.n13093 0.0165714
R49960 VCC.n13154 VCC.n12831 0.0165714
R49961 VCC.n13181 VCC.n13180 0.0165714
R49962 VCC.n13199 VCC.n12805 0.0165714
R49963 VCC.n13259 VCC.n12774 0.0165714
R49964 VCC.n13288 VCC.n12757 0.0165714
R49965 VCC.n13757 VCC.n13756 0.0165714
R49966 VCC.n13823 VCC.n13822 0.0165714
R49967 VCC.n13836 VCC.n13835 0.0165714
R49968 VCC.n13702 VCC.n13701 0.0165714
R49969 VCC.n13630 VCC.n13621 0.0165714
R49970 VCC.n13655 VCC.n13649 0.0165714
R49971 VCC.n13710 VCC.n13387 0.0165714
R49972 VCC.n13738 VCC.n13737 0.0165714
R49973 VCC.n13540 VCC.n13535 0.0165714
R49974 VCC.n13557 VCC.n13556 0.0165714
R49975 VCC.n13506 VCC.n13499 0.0165714
R49976 VCC.n13542 VCC.n13541 0.0165714
R49977 VCC.n13558 VCC.n13469 0.0165714
R49978 VCC.n13584 VCC.n13448 0.0165714
R49979 VCC.n13603 VCC.n13602 0.0165714
R49980 VCC.n14090 VCC.n14085 0.0165714
R49981 VCC.n14107 VCC.n14106 0.0165714
R49982 VCC.n14056 VCC.n14049 0.0165714
R49983 VCC.n14092 VCC.n14091 0.0165714
R49984 VCC.n14108 VCC.n14019 0.0165714
R49985 VCC.n14134 VCC.n13998 0.0165714
R49986 VCC.n14153 VCC.n14152 0.0165714
R49987 VCC.n14253 VCC.n14252 0.0165714
R49988 VCC.n14181 VCC.n14173 0.0165714
R49989 VCC.n14206 VCC.n14200 0.0165714
R49990 VCC.n14261 VCC.n13938 0.0165714
R49991 VCC.n14288 VCC.n14287 0.0165714
R49992 VCC.n14306 VCC.n13912 0.0165714
R49993 VCC.n14366 VCC.n13881 0.0165714
R49994 VCC.n14395 VCC.n13864 0.0165714
R49995 VCC.n14864 VCC.n14863 0.0165714
R49996 VCC.n14930 VCC.n14929 0.0165714
R49997 VCC.n14943 VCC.n14942 0.0165714
R49998 VCC.n14809 VCC.n14808 0.0165714
R49999 VCC.n14737 VCC.n14728 0.0165714
R50000 VCC.n14762 VCC.n14756 0.0165714
R50001 VCC.n14817 VCC.n14494 0.0165714
R50002 VCC.n14845 VCC.n14844 0.0165714
R50003 VCC.n14647 VCC.n14642 0.0165714
R50004 VCC.n14664 VCC.n14663 0.0165714
R50005 VCC.n14613 VCC.n14606 0.0165714
R50006 VCC.n14649 VCC.n14648 0.0165714
R50007 VCC.n14665 VCC.n14576 0.0165714
R50008 VCC.n14691 VCC.n14555 0.0165714
R50009 VCC.n14710 VCC.n14709 0.0165714
R50010 VCC.n15197 VCC.n15192 0.0165714
R50011 VCC.n15214 VCC.n15213 0.0165714
R50012 VCC.n15163 VCC.n15156 0.0165714
R50013 VCC.n15199 VCC.n15198 0.0165714
R50014 VCC.n15215 VCC.n15126 0.0165714
R50015 VCC.n15241 VCC.n15105 0.0165714
R50016 VCC.n15260 VCC.n15259 0.0165714
R50017 VCC.n15360 VCC.n15359 0.0165714
R50018 VCC.n15288 VCC.n15280 0.0165714
R50019 VCC.n15313 VCC.n15307 0.0165714
R50020 VCC.n15368 VCC.n15045 0.0165714
R50021 VCC.n15395 VCC.n15394 0.0165714
R50022 VCC.n15413 VCC.n15019 0.0165714
R50023 VCC.n15473 VCC.n14988 0.0165714
R50024 VCC.n15502 VCC.n14971 0.0165714
R50025 VCC.n15971 VCC.n15970 0.0165714
R50026 VCC.n16037 VCC.n16036 0.0165714
R50027 VCC.n16050 VCC.n16049 0.0165714
R50028 VCC.n15916 VCC.n15915 0.0165714
R50029 VCC.n15844 VCC.n15835 0.0165714
R50030 VCC.n15869 VCC.n15863 0.0165714
R50031 VCC.n15924 VCC.n15601 0.0165714
R50032 VCC.n15952 VCC.n15951 0.0165714
R50033 VCC.n15754 VCC.n15749 0.0165714
R50034 VCC.n15771 VCC.n15770 0.0165714
R50035 VCC.n15720 VCC.n15713 0.0165714
R50036 VCC.n15756 VCC.n15755 0.0165714
R50037 VCC.n15772 VCC.n15683 0.0165714
R50038 VCC.n15798 VCC.n15662 0.0165714
R50039 VCC.n15817 VCC.n15816 0.0165714
R50040 VCC.n16304 VCC.n16299 0.0165714
R50041 VCC.n16321 VCC.n16320 0.0165714
R50042 VCC.n16270 VCC.n16263 0.0165714
R50043 VCC.n16306 VCC.n16305 0.0165714
R50044 VCC.n16322 VCC.n16233 0.0165714
R50045 VCC.n16348 VCC.n16212 0.0165714
R50046 VCC.n16367 VCC.n16366 0.0165714
R50047 VCC.n16467 VCC.n16466 0.0165714
R50048 VCC.n16395 VCC.n16387 0.0165714
R50049 VCC.n16420 VCC.n16414 0.0165714
R50050 VCC.n16475 VCC.n16152 0.0165714
R50051 VCC.n16502 VCC.n16501 0.0165714
R50052 VCC.n16520 VCC.n16126 0.0165714
R50053 VCC.n16580 VCC.n16095 0.0165714
R50054 VCC.n16609 VCC.n16078 0.0165714
R50055 VCC.n17078 VCC.n17077 0.0165714
R50056 VCC.n17144 VCC.n17143 0.0165714
R50057 VCC.n17157 VCC.n17156 0.0165714
R50058 VCC.n17023 VCC.n17022 0.0165714
R50059 VCC.n16951 VCC.n16942 0.0165714
R50060 VCC.n16976 VCC.n16970 0.0165714
R50061 VCC.n17031 VCC.n16708 0.0165714
R50062 VCC.n17059 VCC.n17058 0.0165714
R50063 VCC.n16861 VCC.n16856 0.0165714
R50064 VCC.n16878 VCC.n16877 0.0165714
R50065 VCC.n16827 VCC.n16820 0.0165714
R50066 VCC.n16863 VCC.n16862 0.0165714
R50067 VCC.n16879 VCC.n16790 0.0165714
R50068 VCC.n16905 VCC.n16769 0.0165714
R50069 VCC.n16924 VCC.n16923 0.0165714
R50070 VCC.n17387 VCC.n17386 0.0165714
R50071 VCC.n17315 VCC.n17307 0.0165714
R50072 VCC.n17340 VCC.n17334 0.0165714
R50073 VCC.n17395 VCC.n17259 0.0165714
R50074 VCC.n17422 VCC.n17421 0.0165714
R50075 VCC.n17440 VCC.n17233 0.0165714
R50076 VCC.n17500 VCC.n17202 0.0165714
R50077 VCC.n17529 VCC.n17185 0.0165714
R50078 VCC.n274 VCC.n273 0.0156786
R50079 VCC.n240 VCC.n174 0.0156786
R50080 VCC.n356 VCC.n355 0.0156786
R50081 VCC.n410 VCC.n409 0.0156786
R50082 VCC.n480 VCC.n50 0.0156786
R50083 VCC.n826 VCC.n825 0.0156786
R50084 VCC.n792 VCC.n726 0.0156786
R50085 VCC.n908 VCC.n907 0.0156786
R50086 VCC.n962 VCC.n961 0.0156786
R50087 VCC.n1032 VCC.n602 0.0156786
R50088 VCC.n1598 VCC.n1155 0.0156786
R50089 VCC.n1465 VCC.n1464 0.0156786
R50090 VCC.n1519 VCC.n1518 0.0156786
R50091 VCC.n1384 VCC.n1383 0.0156786
R50092 VCC.n1350 VCC.n1284 0.0156786
R50093 VCC.n1935 VCC.n1934 0.0156786
R50094 VCC.n1901 VCC.n1835 0.0156786
R50095 VCC.n2017 VCC.n2016 0.0156786
R50096 VCC.n2071 VCC.n2070 0.0156786
R50097 VCC.n2141 VCC.n1711 0.0156786
R50098 VCC.n2707 VCC.n2264 0.0156786
R50099 VCC.n2574 VCC.n2573 0.0156786
R50100 VCC.n2628 VCC.n2627 0.0156786
R50101 VCC.n2493 VCC.n2492 0.0156786
R50102 VCC.n2459 VCC.n2393 0.0156786
R50103 VCC.n3044 VCC.n3043 0.0156786
R50104 VCC.n3010 VCC.n2944 0.0156786
R50105 VCC.n3126 VCC.n3125 0.0156786
R50106 VCC.n3180 VCC.n3179 0.0156786
R50107 VCC.n3250 VCC.n2820 0.0156786
R50108 VCC.n3816 VCC.n3373 0.0156786
R50109 VCC.n3683 VCC.n3682 0.0156786
R50110 VCC.n3737 VCC.n3736 0.0156786
R50111 VCC.n3602 VCC.n3601 0.0156786
R50112 VCC.n3568 VCC.n3502 0.0156786
R50113 VCC.n4153 VCC.n4152 0.0156786
R50114 VCC.n4119 VCC.n4053 0.0156786
R50115 VCC.n4235 VCC.n4234 0.0156786
R50116 VCC.n4289 VCC.n4288 0.0156786
R50117 VCC.n4359 VCC.n3929 0.0156786
R50118 VCC.n4925 VCC.n4482 0.0156786
R50119 VCC.n4792 VCC.n4791 0.0156786
R50120 VCC.n4846 VCC.n4845 0.0156786
R50121 VCC.n4711 VCC.n4710 0.0156786
R50122 VCC.n4677 VCC.n4611 0.0156786
R50123 VCC.n5262 VCC.n5261 0.0156786
R50124 VCC.n5228 VCC.n5162 0.0156786
R50125 VCC.n5344 VCC.n5343 0.0156786
R50126 VCC.n5398 VCC.n5397 0.0156786
R50127 VCC.n5468 VCC.n5038 0.0156786
R50128 VCC.n6034 VCC.n5591 0.0156786
R50129 VCC.n5901 VCC.n5900 0.0156786
R50130 VCC.n5955 VCC.n5954 0.0156786
R50131 VCC.n5820 VCC.n5819 0.0156786
R50132 VCC.n5786 VCC.n5720 0.0156786
R50133 VCC.n6371 VCC.n6370 0.0156786
R50134 VCC.n6337 VCC.n6271 0.0156786
R50135 VCC.n6453 VCC.n6452 0.0156786
R50136 VCC.n6507 VCC.n6506 0.0156786
R50137 VCC.n6577 VCC.n6147 0.0156786
R50138 VCC.n7143 VCC.n6700 0.0156786
R50139 VCC.n7010 VCC.n7009 0.0156786
R50140 VCC.n7064 VCC.n7063 0.0156786
R50141 VCC.n6929 VCC.n6928 0.0156786
R50142 VCC.n6895 VCC.n6829 0.0156786
R50143 VCC.n7480 VCC.n7479 0.0156786
R50144 VCC.n7446 VCC.n7380 0.0156786
R50145 VCC.n7562 VCC.n7561 0.0156786
R50146 VCC.n7616 VCC.n7615 0.0156786
R50147 VCC.n7686 VCC.n7256 0.0156786
R50148 VCC.n8252 VCC.n7809 0.0156786
R50149 VCC.n8119 VCC.n8118 0.0156786
R50150 VCC.n8173 VCC.n8172 0.0156786
R50151 VCC.n8038 VCC.n8037 0.0156786
R50152 VCC.n8004 VCC.n7938 0.0156786
R50153 VCC.n8671 VCC.n8670 0.0156786
R50154 VCC.n8725 VCC.n8724 0.0156786
R50155 VCC.n8795 VCC.n8365 0.0156786
R50156 VCC.n8589 VCC.n8588 0.0156786
R50157 VCC.n8555 VCC.n8489 0.0156786
R50158 VCC.n9361 VCC.n8918 0.0156786
R50159 VCC.n9228 VCC.n9227 0.0156786
R50160 VCC.n9282 VCC.n9281 0.0156786
R50161 VCC.n9147 VCC.n9146 0.0156786
R50162 VCC.n9113 VCC.n9047 0.0156786
R50163 VCC.n9698 VCC.n9697 0.0156786
R50164 VCC.n9664 VCC.n9598 0.0156786
R50165 VCC.n9780 VCC.n9779 0.0156786
R50166 VCC.n9834 VCC.n9833 0.0156786
R50167 VCC.n9904 VCC.n9474 0.0156786
R50168 VCC.n10469 VCC.n10026 0.0156786
R50169 VCC.n10336 VCC.n10335 0.0156786
R50170 VCC.n10390 VCC.n10389 0.0156786
R50171 VCC.n10255 VCC.n10254 0.0156786
R50172 VCC.n10221 VCC.n10155 0.0156786
R50173 VCC.n10805 VCC.n10804 0.0156786
R50174 VCC.n10771 VCC.n10705 0.0156786
R50175 VCC.n10887 VCC.n10886 0.0156786
R50176 VCC.n10941 VCC.n10940 0.0156786
R50177 VCC.n11011 VCC.n10581 0.0156786
R50178 VCC.n11576 VCC.n11133 0.0156786
R50179 VCC.n11443 VCC.n11442 0.0156786
R50180 VCC.n11497 VCC.n11496 0.0156786
R50181 VCC.n11362 VCC.n11361 0.0156786
R50182 VCC.n11328 VCC.n11262 0.0156786
R50183 VCC.n11912 VCC.n11911 0.0156786
R50184 VCC.n11878 VCC.n11812 0.0156786
R50185 VCC.n11994 VCC.n11993 0.0156786
R50186 VCC.n12048 VCC.n12047 0.0156786
R50187 VCC.n12118 VCC.n11688 0.0156786
R50188 VCC.n12683 VCC.n12240 0.0156786
R50189 VCC.n12550 VCC.n12549 0.0156786
R50190 VCC.n12604 VCC.n12603 0.0156786
R50191 VCC.n12469 VCC.n12468 0.0156786
R50192 VCC.n12435 VCC.n12369 0.0156786
R50193 VCC.n13019 VCC.n13018 0.0156786
R50194 VCC.n12985 VCC.n12919 0.0156786
R50195 VCC.n13101 VCC.n13100 0.0156786
R50196 VCC.n13155 VCC.n13154 0.0156786
R50197 VCC.n13225 VCC.n12795 0.0156786
R50198 VCC.n13790 VCC.n13347 0.0156786
R50199 VCC.n13657 VCC.n13656 0.0156786
R50200 VCC.n13711 VCC.n13710 0.0156786
R50201 VCC.n13576 VCC.n13575 0.0156786
R50202 VCC.n13542 VCC.n13476 0.0156786
R50203 VCC.n14126 VCC.n14125 0.0156786
R50204 VCC.n14092 VCC.n14026 0.0156786
R50205 VCC.n14208 VCC.n14207 0.0156786
R50206 VCC.n14262 VCC.n14261 0.0156786
R50207 VCC.n14332 VCC.n13902 0.0156786
R50208 VCC.n14897 VCC.n14454 0.0156786
R50209 VCC.n14764 VCC.n14763 0.0156786
R50210 VCC.n14818 VCC.n14817 0.0156786
R50211 VCC.n14683 VCC.n14682 0.0156786
R50212 VCC.n14649 VCC.n14583 0.0156786
R50213 VCC.n15233 VCC.n15232 0.0156786
R50214 VCC.n15199 VCC.n15133 0.0156786
R50215 VCC.n15315 VCC.n15314 0.0156786
R50216 VCC.n15369 VCC.n15368 0.0156786
R50217 VCC.n15439 VCC.n15009 0.0156786
R50218 VCC.n16004 VCC.n15561 0.0156786
R50219 VCC.n15871 VCC.n15870 0.0156786
R50220 VCC.n15925 VCC.n15924 0.0156786
R50221 VCC.n15790 VCC.n15789 0.0156786
R50222 VCC.n15756 VCC.n15690 0.0156786
R50223 VCC.n16340 VCC.n16339 0.0156786
R50224 VCC.n16306 VCC.n16240 0.0156786
R50225 VCC.n16422 VCC.n16421 0.0156786
R50226 VCC.n16476 VCC.n16475 0.0156786
R50227 VCC.n16546 VCC.n16116 0.0156786
R50228 VCC.n17111 VCC.n16668 0.0156786
R50229 VCC.n16978 VCC.n16977 0.0156786
R50230 VCC.n17032 VCC.n17031 0.0156786
R50231 VCC.n16897 VCC.n16896 0.0156786
R50232 VCC.n16863 VCC.n16797 0.0156786
R50233 VCC.n17342 VCC.n17341 0.0156786
R50234 VCC.n17396 VCC.n17395 0.0156786
R50235 VCC.n17466 VCC.n17223 0.0156786
R50236 VCC.n242 VCC.n241 0.0152714
R50237 VCC.n281 VCC.n280 0.0152714
R50238 VCC.n347 VCC.n102 0.0152714
R50239 VCC.n408 VCC.n407 0.0152714
R50240 VCC.n485 VCC.n481 0.0152714
R50241 VCC.n513 VCC.n512 0.0152714
R50242 VCC.n794 VCC.n793 0.0152714
R50243 VCC.n833 VCC.n832 0.0152714
R50244 VCC.n899 VCC.n654 0.0152714
R50245 VCC.n960 VCC.n959 0.0152714
R50246 VCC.n1037 VCC.n1033 0.0152714
R50247 VCC.n1065 VCC.n1064 0.0152714
R50248 VCC.n1352 VCC.n1351 0.0152714
R50249 VCC.n1391 VCC.n1390 0.0152714
R50250 VCC.n1456 VCC.n1211 0.0152714
R50251 VCC.n1517 VCC.n1516 0.0152714
R50252 VCC.n1600 VCC.n1599 0.0152714
R50253 VCC.n1629 VCC.n1628 0.0152714
R50254 VCC.n1903 VCC.n1902 0.0152714
R50255 VCC.n1942 VCC.n1941 0.0152714
R50256 VCC.n2008 VCC.n1763 0.0152714
R50257 VCC.n2069 VCC.n2068 0.0152714
R50258 VCC.n2146 VCC.n2142 0.0152714
R50259 VCC.n2174 VCC.n2173 0.0152714
R50260 VCC.n2461 VCC.n2460 0.0152714
R50261 VCC.n2500 VCC.n2499 0.0152714
R50262 VCC.n2565 VCC.n2320 0.0152714
R50263 VCC.n2626 VCC.n2625 0.0152714
R50264 VCC.n2709 VCC.n2708 0.0152714
R50265 VCC.n2738 VCC.n2737 0.0152714
R50266 VCC.n3012 VCC.n3011 0.0152714
R50267 VCC.n3051 VCC.n3050 0.0152714
R50268 VCC.n3117 VCC.n2872 0.0152714
R50269 VCC.n3178 VCC.n3177 0.0152714
R50270 VCC.n3255 VCC.n3251 0.0152714
R50271 VCC.n3283 VCC.n3282 0.0152714
R50272 VCC.n3570 VCC.n3569 0.0152714
R50273 VCC.n3609 VCC.n3608 0.0152714
R50274 VCC.n3674 VCC.n3429 0.0152714
R50275 VCC.n3735 VCC.n3734 0.0152714
R50276 VCC.n3818 VCC.n3817 0.0152714
R50277 VCC.n3847 VCC.n3846 0.0152714
R50278 VCC.n4121 VCC.n4120 0.0152714
R50279 VCC.n4160 VCC.n4159 0.0152714
R50280 VCC.n4226 VCC.n3981 0.0152714
R50281 VCC.n4287 VCC.n4286 0.0152714
R50282 VCC.n4364 VCC.n4360 0.0152714
R50283 VCC.n4392 VCC.n4391 0.0152714
R50284 VCC.n4679 VCC.n4678 0.0152714
R50285 VCC.n4718 VCC.n4717 0.0152714
R50286 VCC.n4783 VCC.n4538 0.0152714
R50287 VCC.n4844 VCC.n4843 0.0152714
R50288 VCC.n4927 VCC.n4926 0.0152714
R50289 VCC.n4956 VCC.n4955 0.0152714
R50290 VCC.n5230 VCC.n5229 0.0152714
R50291 VCC.n5269 VCC.n5268 0.0152714
R50292 VCC.n5335 VCC.n5090 0.0152714
R50293 VCC.n5396 VCC.n5395 0.0152714
R50294 VCC.n5473 VCC.n5469 0.0152714
R50295 VCC.n5501 VCC.n5500 0.0152714
R50296 VCC.n5788 VCC.n5787 0.0152714
R50297 VCC.n5827 VCC.n5826 0.0152714
R50298 VCC.n5892 VCC.n5647 0.0152714
R50299 VCC.n5953 VCC.n5952 0.0152714
R50300 VCC.n6036 VCC.n6035 0.0152714
R50301 VCC.n6065 VCC.n6064 0.0152714
R50302 VCC.n6339 VCC.n6338 0.0152714
R50303 VCC.n6378 VCC.n6377 0.0152714
R50304 VCC.n6444 VCC.n6199 0.0152714
R50305 VCC.n6505 VCC.n6504 0.0152714
R50306 VCC.n6582 VCC.n6578 0.0152714
R50307 VCC.n6610 VCC.n6609 0.0152714
R50308 VCC.n6897 VCC.n6896 0.0152714
R50309 VCC.n6936 VCC.n6935 0.0152714
R50310 VCC.n7001 VCC.n6756 0.0152714
R50311 VCC.n7062 VCC.n7061 0.0152714
R50312 VCC.n7145 VCC.n7144 0.0152714
R50313 VCC.n7174 VCC.n7173 0.0152714
R50314 VCC.n7448 VCC.n7447 0.0152714
R50315 VCC.n7487 VCC.n7486 0.0152714
R50316 VCC.n7553 VCC.n7308 0.0152714
R50317 VCC.n7614 VCC.n7613 0.0152714
R50318 VCC.n7691 VCC.n7687 0.0152714
R50319 VCC.n7719 VCC.n7718 0.0152714
R50320 VCC.n8006 VCC.n8005 0.0152714
R50321 VCC.n8045 VCC.n8044 0.0152714
R50322 VCC.n8110 VCC.n7865 0.0152714
R50323 VCC.n8171 VCC.n8170 0.0152714
R50324 VCC.n8254 VCC.n8253 0.0152714
R50325 VCC.n8283 VCC.n8282 0.0152714
R50326 VCC.n8662 VCC.n8417 0.0152714
R50327 VCC.n8723 VCC.n8722 0.0152714
R50328 VCC.n8800 VCC.n8796 0.0152714
R50329 VCC.n8828 VCC.n8827 0.0152714
R50330 VCC.n9115 VCC.n9114 0.0152714
R50331 VCC.n9154 VCC.n9153 0.0152714
R50332 VCC.n9219 VCC.n8974 0.0152714
R50333 VCC.n9280 VCC.n9279 0.0152714
R50334 VCC.n9363 VCC.n9362 0.0152714
R50335 VCC.n9392 VCC.n9391 0.0152714
R50336 VCC.n9666 VCC.n9665 0.0152714
R50337 VCC.n9705 VCC.n9704 0.0152714
R50338 VCC.n9771 VCC.n9526 0.0152714
R50339 VCC.n9832 VCC.n9831 0.0152714
R50340 VCC.n9909 VCC.n9905 0.0152714
R50341 VCC.n9937 VCC.n9936 0.0152714
R50342 VCC.n10223 VCC.n10222 0.0152714
R50343 VCC.n10262 VCC.n10261 0.0152714
R50344 VCC.n10327 VCC.n10082 0.0152714
R50345 VCC.n10388 VCC.n10387 0.0152714
R50346 VCC.n10471 VCC.n10470 0.0152714
R50347 VCC.n10500 VCC.n10499 0.0152714
R50348 VCC.n10773 VCC.n10772 0.0152714
R50349 VCC.n10812 VCC.n10811 0.0152714
R50350 VCC.n10878 VCC.n10633 0.0152714
R50351 VCC.n10939 VCC.n10938 0.0152714
R50352 VCC.n11016 VCC.n11012 0.0152714
R50353 VCC.n11044 VCC.n11043 0.0152714
R50354 VCC.n11330 VCC.n11329 0.0152714
R50355 VCC.n11369 VCC.n11368 0.0152714
R50356 VCC.n11434 VCC.n11189 0.0152714
R50357 VCC.n11495 VCC.n11494 0.0152714
R50358 VCC.n11578 VCC.n11577 0.0152714
R50359 VCC.n11607 VCC.n11606 0.0152714
R50360 VCC.n11880 VCC.n11879 0.0152714
R50361 VCC.n11919 VCC.n11918 0.0152714
R50362 VCC.n11985 VCC.n11740 0.0152714
R50363 VCC.n12046 VCC.n12045 0.0152714
R50364 VCC.n12123 VCC.n12119 0.0152714
R50365 VCC.n12151 VCC.n12150 0.0152714
R50366 VCC.n12437 VCC.n12436 0.0152714
R50367 VCC.n12476 VCC.n12475 0.0152714
R50368 VCC.n12541 VCC.n12296 0.0152714
R50369 VCC.n12602 VCC.n12601 0.0152714
R50370 VCC.n12685 VCC.n12684 0.0152714
R50371 VCC.n12714 VCC.n12713 0.0152714
R50372 VCC.n12987 VCC.n12986 0.0152714
R50373 VCC.n13026 VCC.n13025 0.0152714
R50374 VCC.n13092 VCC.n12847 0.0152714
R50375 VCC.n13153 VCC.n13152 0.0152714
R50376 VCC.n13230 VCC.n13226 0.0152714
R50377 VCC.n13258 VCC.n13257 0.0152714
R50378 VCC.n13544 VCC.n13543 0.0152714
R50379 VCC.n13583 VCC.n13582 0.0152714
R50380 VCC.n13648 VCC.n13403 0.0152714
R50381 VCC.n13709 VCC.n13708 0.0152714
R50382 VCC.n13792 VCC.n13791 0.0152714
R50383 VCC.n13821 VCC.n13820 0.0152714
R50384 VCC.n14094 VCC.n14093 0.0152714
R50385 VCC.n14133 VCC.n14132 0.0152714
R50386 VCC.n14199 VCC.n13954 0.0152714
R50387 VCC.n14260 VCC.n14259 0.0152714
R50388 VCC.n14337 VCC.n14333 0.0152714
R50389 VCC.n14365 VCC.n14364 0.0152714
R50390 VCC.n14651 VCC.n14650 0.0152714
R50391 VCC.n14690 VCC.n14689 0.0152714
R50392 VCC.n14755 VCC.n14510 0.0152714
R50393 VCC.n14816 VCC.n14815 0.0152714
R50394 VCC.n14899 VCC.n14898 0.0152714
R50395 VCC.n14928 VCC.n14927 0.0152714
R50396 VCC.n15201 VCC.n15200 0.0152714
R50397 VCC.n15240 VCC.n15239 0.0152714
R50398 VCC.n15306 VCC.n15061 0.0152714
R50399 VCC.n15367 VCC.n15366 0.0152714
R50400 VCC.n15444 VCC.n15440 0.0152714
R50401 VCC.n15472 VCC.n15471 0.0152714
R50402 VCC.n15758 VCC.n15757 0.0152714
R50403 VCC.n15797 VCC.n15796 0.0152714
R50404 VCC.n15862 VCC.n15617 0.0152714
R50405 VCC.n15923 VCC.n15922 0.0152714
R50406 VCC.n16006 VCC.n16005 0.0152714
R50407 VCC.n16035 VCC.n16034 0.0152714
R50408 VCC.n16308 VCC.n16307 0.0152714
R50409 VCC.n16347 VCC.n16346 0.0152714
R50410 VCC.n16413 VCC.n16168 0.0152714
R50411 VCC.n16474 VCC.n16473 0.0152714
R50412 VCC.n16551 VCC.n16547 0.0152714
R50413 VCC.n16579 VCC.n16578 0.0152714
R50414 VCC.n16865 VCC.n16864 0.0152714
R50415 VCC.n16904 VCC.n16903 0.0152714
R50416 VCC.n16969 VCC.n16724 0.0152714
R50417 VCC.n17030 VCC.n17029 0.0152714
R50418 VCC.n17113 VCC.n17112 0.0152714
R50419 VCC.n17142 VCC.n17141 0.0152714
R50420 VCC.n17333 VCC.n17275 0.0152714
R50421 VCC.n17394 VCC.n17393 0.0152714
R50422 VCC.n17471 VCC.n17467 0.0152714
R50423 VCC.n17499 VCC.n17498 0.0152714
R50424 VCC.n8557 VCC.n8556 0.0151667
R50425 VCC.n8596 VCC.n8595 0.0151667
R50426 VCC.n283 VCC.n282 0.0147857
R50427 VCC.n348 VCC.n113 0.0147857
R50428 VCC.n462 VCC.n52 0.0147857
R50429 VCC.n835 VCC.n834 0.0147857
R50430 VCC.n900 VCC.n665 0.0147857
R50431 VCC.n1014 VCC.n604 0.0147857
R50432 VCC.n1168 VCC.n1157 0.0147857
R50433 VCC.n1457 VCC.n1222 0.0147857
R50434 VCC.n1393 VCC.n1392 0.0147857
R50435 VCC.n1944 VCC.n1943 0.0147857
R50436 VCC.n2009 VCC.n1774 0.0147857
R50437 VCC.n2123 VCC.n1713 0.0147857
R50438 VCC.n2277 VCC.n2266 0.0147857
R50439 VCC.n2566 VCC.n2331 0.0147857
R50440 VCC.n2502 VCC.n2501 0.0147857
R50441 VCC.n3053 VCC.n3052 0.0147857
R50442 VCC.n3118 VCC.n2883 0.0147857
R50443 VCC.n3232 VCC.n2822 0.0147857
R50444 VCC.n3386 VCC.n3375 0.0147857
R50445 VCC.n3675 VCC.n3440 0.0147857
R50446 VCC.n3611 VCC.n3610 0.0147857
R50447 VCC.n4162 VCC.n4161 0.0147857
R50448 VCC.n4227 VCC.n3992 0.0147857
R50449 VCC.n4341 VCC.n3931 0.0147857
R50450 VCC.n4495 VCC.n4484 0.0147857
R50451 VCC.n4784 VCC.n4549 0.0147857
R50452 VCC.n4720 VCC.n4719 0.0147857
R50453 VCC.n5271 VCC.n5270 0.0147857
R50454 VCC.n5336 VCC.n5101 0.0147857
R50455 VCC.n5450 VCC.n5040 0.0147857
R50456 VCC.n5604 VCC.n5593 0.0147857
R50457 VCC.n5893 VCC.n5658 0.0147857
R50458 VCC.n5829 VCC.n5828 0.0147857
R50459 VCC.n6380 VCC.n6379 0.0147857
R50460 VCC.n6445 VCC.n6210 0.0147857
R50461 VCC.n6559 VCC.n6149 0.0147857
R50462 VCC.n6713 VCC.n6702 0.0147857
R50463 VCC.n7002 VCC.n6767 0.0147857
R50464 VCC.n6938 VCC.n6937 0.0147857
R50465 VCC.n7489 VCC.n7488 0.0147857
R50466 VCC.n7554 VCC.n7319 0.0147857
R50467 VCC.n7668 VCC.n7258 0.0147857
R50468 VCC.n7822 VCC.n7811 0.0147857
R50469 VCC.n8111 VCC.n7876 0.0147857
R50470 VCC.n8047 VCC.n8046 0.0147857
R50471 VCC.n8663 VCC.n8428 0.0147857
R50472 VCC.n8777 VCC.n8367 0.0147857
R50473 VCC.n8598 VCC.n8597 0.0147857
R50474 VCC.n8931 VCC.n8920 0.0147857
R50475 VCC.n9220 VCC.n8985 0.0147857
R50476 VCC.n9156 VCC.n9155 0.0147857
R50477 VCC.n9707 VCC.n9706 0.0147857
R50478 VCC.n9772 VCC.n9537 0.0147857
R50479 VCC.n9886 VCC.n9476 0.0147857
R50480 VCC.n10039 VCC.n10028 0.0147857
R50481 VCC.n10328 VCC.n10093 0.0147857
R50482 VCC.n10264 VCC.n10263 0.0147857
R50483 VCC.n10814 VCC.n10813 0.0147857
R50484 VCC.n10879 VCC.n10644 0.0147857
R50485 VCC.n10993 VCC.n10583 0.0147857
R50486 VCC.n11146 VCC.n11135 0.0147857
R50487 VCC.n11435 VCC.n11200 0.0147857
R50488 VCC.n11371 VCC.n11370 0.0147857
R50489 VCC.n11921 VCC.n11920 0.0147857
R50490 VCC.n11986 VCC.n11751 0.0147857
R50491 VCC.n12100 VCC.n11690 0.0147857
R50492 VCC.n12253 VCC.n12242 0.0147857
R50493 VCC.n12542 VCC.n12307 0.0147857
R50494 VCC.n12478 VCC.n12477 0.0147857
R50495 VCC.n13028 VCC.n13027 0.0147857
R50496 VCC.n13093 VCC.n12858 0.0147857
R50497 VCC.n13207 VCC.n12797 0.0147857
R50498 VCC.n13360 VCC.n13349 0.0147857
R50499 VCC.n13649 VCC.n13414 0.0147857
R50500 VCC.n13585 VCC.n13584 0.0147857
R50501 VCC.n14135 VCC.n14134 0.0147857
R50502 VCC.n14200 VCC.n13965 0.0147857
R50503 VCC.n14314 VCC.n13904 0.0147857
R50504 VCC.n14467 VCC.n14456 0.0147857
R50505 VCC.n14756 VCC.n14521 0.0147857
R50506 VCC.n14692 VCC.n14691 0.0147857
R50507 VCC.n15242 VCC.n15241 0.0147857
R50508 VCC.n15307 VCC.n15072 0.0147857
R50509 VCC.n15421 VCC.n15011 0.0147857
R50510 VCC.n15574 VCC.n15563 0.0147857
R50511 VCC.n15863 VCC.n15628 0.0147857
R50512 VCC.n15799 VCC.n15798 0.0147857
R50513 VCC.n16349 VCC.n16348 0.0147857
R50514 VCC.n16414 VCC.n16179 0.0147857
R50515 VCC.n16528 VCC.n16118 0.0147857
R50516 VCC.n16681 VCC.n16670 0.0147857
R50517 VCC.n16970 VCC.n16735 0.0147857
R50518 VCC.n16906 VCC.n16905 0.0147857
R50519 VCC.n17334 VCC.n17286 0.0147857
R50520 VCC.n17448 VCC.n17225 0.0147857
R50521 VCC.n258 VCC.n257 0.0132571
R50522 VCC.n380 VCC.n379 0.0132571
R50523 VCC.n504 VCC.n503 0.0132571
R50524 VCC.n810 VCC.n809 0.0132571
R50525 VCC.n932 VCC.n931 0.0132571
R50526 VCC.n1056 VCC.n1055 0.0132571
R50527 VCC.n1368 VCC.n1367 0.0132571
R50528 VCC.n1489 VCC.n1488 0.0132571
R50529 VCC.n1612 VCC.n1608 0.0132571
R50530 VCC.n1919 VCC.n1918 0.0132571
R50531 VCC.n2041 VCC.n2040 0.0132571
R50532 VCC.n2165 VCC.n2164 0.0132571
R50533 VCC.n2477 VCC.n2476 0.0132571
R50534 VCC.n2598 VCC.n2597 0.0132571
R50535 VCC.n2721 VCC.n2717 0.0132571
R50536 VCC.n3028 VCC.n3027 0.0132571
R50537 VCC.n3150 VCC.n3149 0.0132571
R50538 VCC.n3274 VCC.n3273 0.0132571
R50539 VCC.n3586 VCC.n3585 0.0132571
R50540 VCC.n3707 VCC.n3706 0.0132571
R50541 VCC.n3830 VCC.n3826 0.0132571
R50542 VCC.n4137 VCC.n4136 0.0132571
R50543 VCC.n4259 VCC.n4258 0.0132571
R50544 VCC.n4383 VCC.n4382 0.0132571
R50545 VCC.n4695 VCC.n4694 0.0132571
R50546 VCC.n4816 VCC.n4815 0.0132571
R50547 VCC.n4939 VCC.n4935 0.0132571
R50548 VCC.n5246 VCC.n5245 0.0132571
R50549 VCC.n5368 VCC.n5367 0.0132571
R50550 VCC.n5492 VCC.n5491 0.0132571
R50551 VCC.n5804 VCC.n5803 0.0132571
R50552 VCC.n5925 VCC.n5924 0.0132571
R50553 VCC.n6048 VCC.n6044 0.0132571
R50554 VCC.n6355 VCC.n6354 0.0132571
R50555 VCC.n6477 VCC.n6476 0.0132571
R50556 VCC.n6601 VCC.n6600 0.0132571
R50557 VCC.n6913 VCC.n6912 0.0132571
R50558 VCC.n7034 VCC.n7033 0.0132571
R50559 VCC.n7157 VCC.n7153 0.0132571
R50560 VCC.n7464 VCC.n7463 0.0132571
R50561 VCC.n7586 VCC.n7585 0.0132571
R50562 VCC.n7710 VCC.n7709 0.0132571
R50563 VCC.n8022 VCC.n8021 0.0132571
R50564 VCC.n8143 VCC.n8142 0.0132571
R50565 VCC.n8266 VCC.n8262 0.0132571
R50566 VCC.n8695 VCC.n8694 0.0132571
R50567 VCC.n8819 VCC.n8818 0.0132571
R50568 VCC.n9131 VCC.n9130 0.0132571
R50569 VCC.n9252 VCC.n9251 0.0132571
R50570 VCC.n9375 VCC.n9371 0.0132571
R50571 VCC.n9682 VCC.n9681 0.0132571
R50572 VCC.n9804 VCC.n9803 0.0132571
R50573 VCC.n9928 VCC.n9927 0.0132571
R50574 VCC.n10239 VCC.n10238 0.0132571
R50575 VCC.n10360 VCC.n10359 0.0132571
R50576 VCC.n10483 VCC.n10479 0.0132571
R50577 VCC.n10789 VCC.n10788 0.0132571
R50578 VCC.n10911 VCC.n10910 0.0132571
R50579 VCC.n11035 VCC.n11034 0.0132571
R50580 VCC.n11346 VCC.n11345 0.0132571
R50581 VCC.n11467 VCC.n11466 0.0132571
R50582 VCC.n11590 VCC.n11586 0.0132571
R50583 VCC.n11896 VCC.n11895 0.0132571
R50584 VCC.n12018 VCC.n12017 0.0132571
R50585 VCC.n12142 VCC.n12141 0.0132571
R50586 VCC.n12453 VCC.n12452 0.0132571
R50587 VCC.n12574 VCC.n12573 0.0132571
R50588 VCC.n12697 VCC.n12693 0.0132571
R50589 VCC.n13003 VCC.n13002 0.0132571
R50590 VCC.n13125 VCC.n13124 0.0132571
R50591 VCC.n13249 VCC.n13248 0.0132571
R50592 VCC.n13560 VCC.n13559 0.0132571
R50593 VCC.n13681 VCC.n13680 0.0132571
R50594 VCC.n13804 VCC.n13800 0.0132571
R50595 VCC.n14110 VCC.n14109 0.0132571
R50596 VCC.n14232 VCC.n14231 0.0132571
R50597 VCC.n14356 VCC.n14355 0.0132571
R50598 VCC.n14667 VCC.n14666 0.0132571
R50599 VCC.n14788 VCC.n14787 0.0132571
R50600 VCC.n14911 VCC.n14907 0.0132571
R50601 VCC.n15217 VCC.n15216 0.0132571
R50602 VCC.n15339 VCC.n15338 0.0132571
R50603 VCC.n15463 VCC.n15462 0.0132571
R50604 VCC.n15774 VCC.n15773 0.0132571
R50605 VCC.n15895 VCC.n15894 0.0132571
R50606 VCC.n16018 VCC.n16014 0.0132571
R50607 VCC.n16324 VCC.n16323 0.0132571
R50608 VCC.n16446 VCC.n16445 0.0132571
R50609 VCC.n16570 VCC.n16569 0.0132571
R50610 VCC.n16881 VCC.n16880 0.0132571
R50611 VCC.n17002 VCC.n17001 0.0132571
R50612 VCC.n17125 VCC.n17121 0.0132571
R50613 VCC.n17366 VCC.n17365 0.0132571
R50614 VCC.n17490 VCC.n17489 0.0132571
R50615 VCC.n8573 VCC.n8572 0.0131667
R50616 VCC.n202 VCC.n200 0.013
R50617 VCC.n76 VCC.n74 0.013
R50618 VCC.n542 VCC.n9 0.013
R50619 VCC.n550 VCC.n2 0.013
R50620 VCC.n541 VCC.n540 0.013
R50621 VCC.n754 VCC.n752 0.013
R50622 VCC.n628 VCC.n626 0.013
R50623 VCC.n1096 VCC.n563 0.013
R50624 VCC.n1104 VCC.n556 0.013
R50625 VCC.n1095 VCC.n1094 0.013
R50626 VCC.n1642 VCC.n1641 0.013
R50627 VCC.n1658 VCC.n1110 0.013
R50628 VCC.n1643 VCC.n1121 0.013
R50629 VCC.n1185 VCC.n1183 0.013
R50630 VCC.n1312 VCC.n1310 0.013
R50631 VCC.n1863 VCC.n1861 0.013
R50632 VCC.n1737 VCC.n1735 0.013
R50633 VCC.n2205 VCC.n1672 0.013
R50634 VCC.n2213 VCC.n1665 0.013
R50635 VCC.n2204 VCC.n2203 0.013
R50636 VCC.n2751 VCC.n2750 0.013
R50637 VCC.n2767 VCC.n2219 0.013
R50638 VCC.n2752 VCC.n2230 0.013
R50639 VCC.n2294 VCC.n2292 0.013
R50640 VCC.n2421 VCC.n2419 0.013
R50641 VCC.n2972 VCC.n2970 0.013
R50642 VCC.n2846 VCC.n2844 0.013
R50643 VCC.n3314 VCC.n2781 0.013
R50644 VCC.n3322 VCC.n2774 0.013
R50645 VCC.n3313 VCC.n3312 0.013
R50646 VCC.n3860 VCC.n3859 0.013
R50647 VCC.n3876 VCC.n3328 0.013
R50648 VCC.n3861 VCC.n3339 0.013
R50649 VCC.n3403 VCC.n3401 0.013
R50650 VCC.n3530 VCC.n3528 0.013
R50651 VCC.n4081 VCC.n4079 0.013
R50652 VCC.n3955 VCC.n3953 0.013
R50653 VCC.n4423 VCC.n3890 0.013
R50654 VCC.n4431 VCC.n3883 0.013
R50655 VCC.n4422 VCC.n4421 0.013
R50656 VCC.n4969 VCC.n4968 0.013
R50657 VCC.n4985 VCC.n4437 0.013
R50658 VCC.n4970 VCC.n4448 0.013
R50659 VCC.n4512 VCC.n4510 0.013
R50660 VCC.n4639 VCC.n4637 0.013
R50661 VCC.n5190 VCC.n5188 0.013
R50662 VCC.n5064 VCC.n5062 0.013
R50663 VCC.n5532 VCC.n4999 0.013
R50664 VCC.n5540 VCC.n4992 0.013
R50665 VCC.n5531 VCC.n5530 0.013
R50666 VCC.n6078 VCC.n6077 0.013
R50667 VCC.n6094 VCC.n5546 0.013
R50668 VCC.n6079 VCC.n5557 0.013
R50669 VCC.n5621 VCC.n5619 0.013
R50670 VCC.n5748 VCC.n5746 0.013
R50671 VCC.n6299 VCC.n6297 0.013
R50672 VCC.n6173 VCC.n6171 0.013
R50673 VCC.n6641 VCC.n6108 0.013
R50674 VCC.n6649 VCC.n6101 0.013
R50675 VCC.n6640 VCC.n6639 0.013
R50676 VCC.n7187 VCC.n7186 0.013
R50677 VCC.n7203 VCC.n6655 0.013
R50678 VCC.n7188 VCC.n6666 0.013
R50679 VCC.n6730 VCC.n6728 0.013
R50680 VCC.n6857 VCC.n6855 0.013
R50681 VCC.n7408 VCC.n7406 0.013
R50682 VCC.n7282 VCC.n7280 0.013
R50683 VCC.n7750 VCC.n7217 0.013
R50684 VCC.n7758 VCC.n7210 0.013
R50685 VCC.n7749 VCC.n7748 0.013
R50686 VCC.n8296 VCC.n8295 0.013
R50687 VCC.n8312 VCC.n7764 0.013
R50688 VCC.n8297 VCC.n7775 0.013
R50689 VCC.n7839 VCC.n7837 0.013
R50690 VCC.n7966 VCC.n7964 0.013
R50691 VCC.n8391 VCC.n8389 0.013
R50692 VCC.n8859 VCC.n8326 0.013
R50693 VCC.n8867 VCC.n8319 0.013
R50694 VCC.n8858 VCC.n8857 0.013
R50695 VCC.n8517 VCC.n8515 0.013
R50696 VCC.n9405 VCC.n9404 0.013
R50697 VCC.n9421 VCC.n8873 0.013
R50698 VCC.n9406 VCC.n8884 0.013
R50699 VCC.n8948 VCC.n8946 0.013
R50700 VCC.n9075 VCC.n9073 0.013
R50701 VCC.n9626 VCC.n9624 0.013
R50702 VCC.n9500 VCC.n9498 0.013
R50703 VCC.n9968 VCC.n9435 0.013
R50704 VCC.n9976 VCC.n9428 0.013
R50705 VCC.n9967 VCC.n9966 0.013
R50706 VCC.n10513 VCC.n10512 0.013
R50707 VCC.n10529 VCC.n9981 0.013
R50708 VCC.n10514 VCC.n9992 0.013
R50709 VCC.n10056 VCC.n10054 0.013
R50710 VCC.n10183 VCC.n10181 0.013
R50711 VCC.n10733 VCC.n10731 0.013
R50712 VCC.n10607 VCC.n10605 0.013
R50713 VCC.n11075 VCC.n10542 0.013
R50714 VCC.n11083 VCC.n10535 0.013
R50715 VCC.n11074 VCC.n11073 0.013
R50716 VCC.n11620 VCC.n11619 0.013
R50717 VCC.n11636 VCC.n11088 0.013
R50718 VCC.n11621 VCC.n11099 0.013
R50719 VCC.n11163 VCC.n11161 0.013
R50720 VCC.n11290 VCC.n11288 0.013
R50721 VCC.n11840 VCC.n11838 0.013
R50722 VCC.n11714 VCC.n11712 0.013
R50723 VCC.n12182 VCC.n11649 0.013
R50724 VCC.n12190 VCC.n11642 0.013
R50725 VCC.n12181 VCC.n12180 0.013
R50726 VCC.n12727 VCC.n12726 0.013
R50727 VCC.n12743 VCC.n12195 0.013
R50728 VCC.n12728 VCC.n12206 0.013
R50729 VCC.n12270 VCC.n12268 0.013
R50730 VCC.n12397 VCC.n12395 0.013
R50731 VCC.n12947 VCC.n12945 0.013
R50732 VCC.n12821 VCC.n12819 0.013
R50733 VCC.n13289 VCC.n12756 0.013
R50734 VCC.n13297 VCC.n12749 0.013
R50735 VCC.n13288 VCC.n13287 0.013
R50736 VCC.n13834 VCC.n13833 0.013
R50737 VCC.n13850 VCC.n13302 0.013
R50738 VCC.n13835 VCC.n13313 0.013
R50739 VCC.n13377 VCC.n13375 0.013
R50740 VCC.n13504 VCC.n13502 0.013
R50741 VCC.n14054 VCC.n14052 0.013
R50742 VCC.n13928 VCC.n13926 0.013
R50743 VCC.n14396 VCC.n13863 0.013
R50744 VCC.n14404 VCC.n13856 0.013
R50745 VCC.n14395 VCC.n14394 0.013
R50746 VCC.n14941 VCC.n14940 0.013
R50747 VCC.n14957 VCC.n14409 0.013
R50748 VCC.n14942 VCC.n14420 0.013
R50749 VCC.n14484 VCC.n14482 0.013
R50750 VCC.n14611 VCC.n14609 0.013
R50751 VCC.n15161 VCC.n15159 0.013
R50752 VCC.n15035 VCC.n15033 0.013
R50753 VCC.n15503 VCC.n14970 0.013
R50754 VCC.n15511 VCC.n14963 0.013
R50755 VCC.n15502 VCC.n15501 0.013
R50756 VCC.n16048 VCC.n16047 0.013
R50757 VCC.n16064 VCC.n15516 0.013
R50758 VCC.n16049 VCC.n15527 0.013
R50759 VCC.n15591 VCC.n15589 0.013
R50760 VCC.n15718 VCC.n15716 0.013
R50761 VCC.n16268 VCC.n16266 0.013
R50762 VCC.n16142 VCC.n16140 0.013
R50763 VCC.n16610 VCC.n16077 0.013
R50764 VCC.n16618 VCC.n16070 0.013
R50765 VCC.n16609 VCC.n16608 0.013
R50766 VCC.n17155 VCC.n17154 0.013
R50767 VCC.n17171 VCC.n16623 0.013
R50768 VCC.n17156 VCC.n16634 0.013
R50769 VCC.n16698 VCC.n16696 0.013
R50770 VCC.n16825 VCC.n16823 0.013
R50771 VCC.n17249 VCC.n17247 0.013
R50772 VCC.n17530 VCC.n17184 0.013
R50773 VCC.n17538 VCC.n17177 0.013
R50774 VCC.n17529 VCC.n17528 0.013
R50775 VCC.n137 VCC.n135 0.0121071
R50776 VCC.n205 VCC.n204 0.0121071
R50777 VCC.n327 VCC.n324 0.0121071
R50778 VCC.n446 VCC.n445 0.0121071
R50779 VCC.n435 VCC.n75 0.0121071
R50780 VCC.n458 VCC.n451 0.0121071
R50781 VCC.n456 VCC.n453 0.0121071
R50782 VCC.n455 VCC.n454 0.0121071
R50783 VCC.n18 VCC.n15 0.0121071
R50784 VCC.n689 VCC.n687 0.0121071
R50785 VCC.n757 VCC.n756 0.0121071
R50786 VCC.n879 VCC.n876 0.0121071
R50787 VCC.n998 VCC.n997 0.0121071
R50788 VCC.n987 VCC.n627 0.0121071
R50789 VCC.n1010 VCC.n1003 0.0121071
R50790 VCC.n1008 VCC.n1005 0.0121071
R50791 VCC.n1007 VCC.n1006 0.0121071
R50792 VCC.n570 VCC.n567 0.0121071
R50793 VCC.n1569 VCC.n1561 0.0121071
R50794 VCC.n1567 VCC.n1563 0.0121071
R50795 VCC.n1566 VCC.n1565 0.0121071
R50796 VCC.n1645 VCC.n1120 0.0121071
R50797 VCC.n1436 VCC.n1433 0.0121071
R50798 VCC.n1556 VCC.n1555 0.0121071
R50799 VCC.n1545 VCC.n1184 0.0121071
R50800 VCC.n1247 VCC.n1245 0.0121071
R50801 VCC.n1315 VCC.n1314 0.0121071
R50802 VCC.n1798 VCC.n1796 0.0121071
R50803 VCC.n1866 VCC.n1865 0.0121071
R50804 VCC.n1988 VCC.n1985 0.0121071
R50805 VCC.n2107 VCC.n2106 0.0121071
R50806 VCC.n2096 VCC.n1736 0.0121071
R50807 VCC.n2119 VCC.n2112 0.0121071
R50808 VCC.n2117 VCC.n2114 0.0121071
R50809 VCC.n2116 VCC.n2115 0.0121071
R50810 VCC.n1679 VCC.n1676 0.0121071
R50811 VCC.n2678 VCC.n2670 0.0121071
R50812 VCC.n2676 VCC.n2672 0.0121071
R50813 VCC.n2675 VCC.n2674 0.0121071
R50814 VCC.n2754 VCC.n2229 0.0121071
R50815 VCC.n2545 VCC.n2542 0.0121071
R50816 VCC.n2665 VCC.n2664 0.0121071
R50817 VCC.n2654 VCC.n2293 0.0121071
R50818 VCC.n2356 VCC.n2354 0.0121071
R50819 VCC.n2424 VCC.n2423 0.0121071
R50820 VCC.n2907 VCC.n2905 0.0121071
R50821 VCC.n2975 VCC.n2974 0.0121071
R50822 VCC.n3097 VCC.n3094 0.0121071
R50823 VCC.n3216 VCC.n3215 0.0121071
R50824 VCC.n3205 VCC.n2845 0.0121071
R50825 VCC.n3228 VCC.n3221 0.0121071
R50826 VCC.n3226 VCC.n3223 0.0121071
R50827 VCC.n3225 VCC.n3224 0.0121071
R50828 VCC.n2788 VCC.n2785 0.0121071
R50829 VCC.n3787 VCC.n3779 0.0121071
R50830 VCC.n3785 VCC.n3781 0.0121071
R50831 VCC.n3784 VCC.n3783 0.0121071
R50832 VCC.n3863 VCC.n3338 0.0121071
R50833 VCC.n3654 VCC.n3651 0.0121071
R50834 VCC.n3774 VCC.n3773 0.0121071
R50835 VCC.n3763 VCC.n3402 0.0121071
R50836 VCC.n3465 VCC.n3463 0.0121071
R50837 VCC.n3533 VCC.n3532 0.0121071
R50838 VCC.n4016 VCC.n4014 0.0121071
R50839 VCC.n4084 VCC.n4083 0.0121071
R50840 VCC.n4206 VCC.n4203 0.0121071
R50841 VCC.n4325 VCC.n4324 0.0121071
R50842 VCC.n4314 VCC.n3954 0.0121071
R50843 VCC.n4337 VCC.n4330 0.0121071
R50844 VCC.n4335 VCC.n4332 0.0121071
R50845 VCC.n4334 VCC.n4333 0.0121071
R50846 VCC.n3897 VCC.n3894 0.0121071
R50847 VCC.n4896 VCC.n4888 0.0121071
R50848 VCC.n4894 VCC.n4890 0.0121071
R50849 VCC.n4893 VCC.n4892 0.0121071
R50850 VCC.n4972 VCC.n4447 0.0121071
R50851 VCC.n4763 VCC.n4760 0.0121071
R50852 VCC.n4883 VCC.n4882 0.0121071
R50853 VCC.n4872 VCC.n4511 0.0121071
R50854 VCC.n4574 VCC.n4572 0.0121071
R50855 VCC.n4642 VCC.n4641 0.0121071
R50856 VCC.n5125 VCC.n5123 0.0121071
R50857 VCC.n5193 VCC.n5192 0.0121071
R50858 VCC.n5315 VCC.n5312 0.0121071
R50859 VCC.n5434 VCC.n5433 0.0121071
R50860 VCC.n5423 VCC.n5063 0.0121071
R50861 VCC.n5446 VCC.n5439 0.0121071
R50862 VCC.n5444 VCC.n5441 0.0121071
R50863 VCC.n5443 VCC.n5442 0.0121071
R50864 VCC.n5006 VCC.n5003 0.0121071
R50865 VCC.n6005 VCC.n5997 0.0121071
R50866 VCC.n6003 VCC.n5999 0.0121071
R50867 VCC.n6002 VCC.n6001 0.0121071
R50868 VCC.n6081 VCC.n5556 0.0121071
R50869 VCC.n5872 VCC.n5869 0.0121071
R50870 VCC.n5992 VCC.n5991 0.0121071
R50871 VCC.n5981 VCC.n5620 0.0121071
R50872 VCC.n5683 VCC.n5681 0.0121071
R50873 VCC.n5751 VCC.n5750 0.0121071
R50874 VCC.n6234 VCC.n6232 0.0121071
R50875 VCC.n6302 VCC.n6301 0.0121071
R50876 VCC.n6424 VCC.n6421 0.0121071
R50877 VCC.n6543 VCC.n6542 0.0121071
R50878 VCC.n6532 VCC.n6172 0.0121071
R50879 VCC.n6555 VCC.n6548 0.0121071
R50880 VCC.n6553 VCC.n6550 0.0121071
R50881 VCC.n6552 VCC.n6551 0.0121071
R50882 VCC.n6115 VCC.n6112 0.0121071
R50883 VCC.n7114 VCC.n7106 0.0121071
R50884 VCC.n7112 VCC.n7108 0.0121071
R50885 VCC.n7111 VCC.n7110 0.0121071
R50886 VCC.n7190 VCC.n6665 0.0121071
R50887 VCC.n6981 VCC.n6978 0.0121071
R50888 VCC.n7101 VCC.n7100 0.0121071
R50889 VCC.n7090 VCC.n6729 0.0121071
R50890 VCC.n6792 VCC.n6790 0.0121071
R50891 VCC.n6860 VCC.n6859 0.0121071
R50892 VCC.n7343 VCC.n7341 0.0121071
R50893 VCC.n7411 VCC.n7410 0.0121071
R50894 VCC.n7533 VCC.n7530 0.0121071
R50895 VCC.n7652 VCC.n7651 0.0121071
R50896 VCC.n7641 VCC.n7281 0.0121071
R50897 VCC.n7664 VCC.n7657 0.0121071
R50898 VCC.n7662 VCC.n7659 0.0121071
R50899 VCC.n7661 VCC.n7660 0.0121071
R50900 VCC.n7224 VCC.n7221 0.0121071
R50901 VCC.n8223 VCC.n8215 0.0121071
R50902 VCC.n8221 VCC.n8217 0.0121071
R50903 VCC.n8220 VCC.n8219 0.0121071
R50904 VCC.n8299 VCC.n7774 0.0121071
R50905 VCC.n8090 VCC.n8087 0.0121071
R50906 VCC.n8210 VCC.n8209 0.0121071
R50907 VCC.n8199 VCC.n7838 0.0121071
R50908 VCC.n7901 VCC.n7899 0.0121071
R50909 VCC.n7969 VCC.n7968 0.0121071
R50910 VCC.n8642 VCC.n8639 0.0121071
R50911 VCC.n8761 VCC.n8760 0.0121071
R50912 VCC.n8750 VCC.n8390 0.0121071
R50913 VCC.n8773 VCC.n8766 0.0121071
R50914 VCC.n8771 VCC.n8768 0.0121071
R50915 VCC.n8770 VCC.n8769 0.0121071
R50916 VCC.n8333 VCC.n8330 0.0121071
R50917 VCC.n8452 VCC.n8450 0.0121071
R50918 VCC.n8520 VCC.n8519 0.0121071
R50919 VCC.n9332 VCC.n9324 0.0121071
R50920 VCC.n9330 VCC.n9326 0.0121071
R50921 VCC.n9329 VCC.n9328 0.0121071
R50922 VCC.n9408 VCC.n8883 0.0121071
R50923 VCC.n9199 VCC.n9196 0.0121071
R50924 VCC.n9319 VCC.n9318 0.0121071
R50925 VCC.n9308 VCC.n8947 0.0121071
R50926 VCC.n9010 VCC.n9008 0.0121071
R50927 VCC.n9078 VCC.n9077 0.0121071
R50928 VCC.n9561 VCC.n9559 0.0121071
R50929 VCC.n9629 VCC.n9628 0.0121071
R50930 VCC.n9751 VCC.n9748 0.0121071
R50931 VCC.n9870 VCC.n9869 0.0121071
R50932 VCC.n9859 VCC.n9499 0.0121071
R50933 VCC.n9882 VCC.n9875 0.0121071
R50934 VCC.n9880 VCC.n9877 0.0121071
R50935 VCC.n9879 VCC.n9878 0.0121071
R50936 VCC.n9442 VCC.n9439 0.0121071
R50937 VCC.n10440 VCC.n10432 0.0121071
R50938 VCC.n10438 VCC.n10434 0.0121071
R50939 VCC.n10437 VCC.n10436 0.0121071
R50940 VCC.n10516 VCC.n9991 0.0121071
R50941 VCC.n10307 VCC.n10304 0.0121071
R50942 VCC.n10427 VCC.n10426 0.0121071
R50943 VCC.n10416 VCC.n10055 0.0121071
R50944 VCC.n10118 VCC.n10116 0.0121071
R50945 VCC.n10186 VCC.n10185 0.0121071
R50946 VCC.n10668 VCC.n10666 0.0121071
R50947 VCC.n10736 VCC.n10735 0.0121071
R50948 VCC.n10858 VCC.n10855 0.0121071
R50949 VCC.n10977 VCC.n10976 0.0121071
R50950 VCC.n10966 VCC.n10606 0.0121071
R50951 VCC.n10989 VCC.n10982 0.0121071
R50952 VCC.n10987 VCC.n10984 0.0121071
R50953 VCC.n10986 VCC.n10985 0.0121071
R50954 VCC.n10549 VCC.n10546 0.0121071
R50955 VCC.n11547 VCC.n11539 0.0121071
R50956 VCC.n11545 VCC.n11541 0.0121071
R50957 VCC.n11544 VCC.n11543 0.0121071
R50958 VCC.n11623 VCC.n11098 0.0121071
R50959 VCC.n11414 VCC.n11411 0.0121071
R50960 VCC.n11534 VCC.n11533 0.0121071
R50961 VCC.n11523 VCC.n11162 0.0121071
R50962 VCC.n11225 VCC.n11223 0.0121071
R50963 VCC.n11293 VCC.n11292 0.0121071
R50964 VCC.n11775 VCC.n11773 0.0121071
R50965 VCC.n11843 VCC.n11842 0.0121071
R50966 VCC.n11965 VCC.n11962 0.0121071
R50967 VCC.n12084 VCC.n12083 0.0121071
R50968 VCC.n12073 VCC.n11713 0.0121071
R50969 VCC.n12096 VCC.n12089 0.0121071
R50970 VCC.n12094 VCC.n12091 0.0121071
R50971 VCC.n12093 VCC.n12092 0.0121071
R50972 VCC.n11656 VCC.n11653 0.0121071
R50973 VCC.n12654 VCC.n12646 0.0121071
R50974 VCC.n12652 VCC.n12648 0.0121071
R50975 VCC.n12651 VCC.n12650 0.0121071
R50976 VCC.n12730 VCC.n12205 0.0121071
R50977 VCC.n12521 VCC.n12518 0.0121071
R50978 VCC.n12641 VCC.n12640 0.0121071
R50979 VCC.n12630 VCC.n12269 0.0121071
R50980 VCC.n12332 VCC.n12330 0.0121071
R50981 VCC.n12400 VCC.n12399 0.0121071
R50982 VCC.n12882 VCC.n12880 0.0121071
R50983 VCC.n12950 VCC.n12949 0.0121071
R50984 VCC.n13072 VCC.n13069 0.0121071
R50985 VCC.n13191 VCC.n13190 0.0121071
R50986 VCC.n13180 VCC.n12820 0.0121071
R50987 VCC.n13203 VCC.n13196 0.0121071
R50988 VCC.n13201 VCC.n13198 0.0121071
R50989 VCC.n13200 VCC.n13199 0.0121071
R50990 VCC.n12763 VCC.n12760 0.0121071
R50991 VCC.n13761 VCC.n13753 0.0121071
R50992 VCC.n13759 VCC.n13755 0.0121071
R50993 VCC.n13758 VCC.n13757 0.0121071
R50994 VCC.n13837 VCC.n13312 0.0121071
R50995 VCC.n13628 VCC.n13625 0.0121071
R50996 VCC.n13748 VCC.n13747 0.0121071
R50997 VCC.n13737 VCC.n13376 0.0121071
R50998 VCC.n13439 VCC.n13437 0.0121071
R50999 VCC.n13507 VCC.n13506 0.0121071
R51000 VCC.n13989 VCC.n13987 0.0121071
R51001 VCC.n14057 VCC.n14056 0.0121071
R51002 VCC.n14179 VCC.n14176 0.0121071
R51003 VCC.n14298 VCC.n14297 0.0121071
R51004 VCC.n14287 VCC.n13927 0.0121071
R51005 VCC.n14310 VCC.n14303 0.0121071
R51006 VCC.n14308 VCC.n14305 0.0121071
R51007 VCC.n14307 VCC.n14306 0.0121071
R51008 VCC.n13870 VCC.n13867 0.0121071
R51009 VCC.n14868 VCC.n14860 0.0121071
R51010 VCC.n14866 VCC.n14862 0.0121071
R51011 VCC.n14865 VCC.n14864 0.0121071
R51012 VCC.n14944 VCC.n14419 0.0121071
R51013 VCC.n14735 VCC.n14732 0.0121071
R51014 VCC.n14855 VCC.n14854 0.0121071
R51015 VCC.n14844 VCC.n14483 0.0121071
R51016 VCC.n14546 VCC.n14544 0.0121071
R51017 VCC.n14614 VCC.n14613 0.0121071
R51018 VCC.n15096 VCC.n15094 0.0121071
R51019 VCC.n15164 VCC.n15163 0.0121071
R51020 VCC.n15286 VCC.n15283 0.0121071
R51021 VCC.n15405 VCC.n15404 0.0121071
R51022 VCC.n15394 VCC.n15034 0.0121071
R51023 VCC.n15417 VCC.n15410 0.0121071
R51024 VCC.n15415 VCC.n15412 0.0121071
R51025 VCC.n15414 VCC.n15413 0.0121071
R51026 VCC.n14977 VCC.n14974 0.0121071
R51027 VCC.n15975 VCC.n15967 0.0121071
R51028 VCC.n15973 VCC.n15969 0.0121071
R51029 VCC.n15972 VCC.n15971 0.0121071
R51030 VCC.n16051 VCC.n15526 0.0121071
R51031 VCC.n15842 VCC.n15839 0.0121071
R51032 VCC.n15962 VCC.n15961 0.0121071
R51033 VCC.n15951 VCC.n15590 0.0121071
R51034 VCC.n15653 VCC.n15651 0.0121071
R51035 VCC.n15721 VCC.n15720 0.0121071
R51036 VCC.n16203 VCC.n16201 0.0121071
R51037 VCC.n16271 VCC.n16270 0.0121071
R51038 VCC.n16393 VCC.n16390 0.0121071
R51039 VCC.n16512 VCC.n16511 0.0121071
R51040 VCC.n16501 VCC.n16141 0.0121071
R51041 VCC.n16524 VCC.n16517 0.0121071
R51042 VCC.n16522 VCC.n16519 0.0121071
R51043 VCC.n16521 VCC.n16520 0.0121071
R51044 VCC.n16084 VCC.n16081 0.0121071
R51045 VCC.n17082 VCC.n17074 0.0121071
R51046 VCC.n17080 VCC.n17076 0.0121071
R51047 VCC.n17079 VCC.n17078 0.0121071
R51048 VCC.n17158 VCC.n16633 0.0121071
R51049 VCC.n16949 VCC.n16946 0.0121071
R51050 VCC.n17069 VCC.n17068 0.0121071
R51051 VCC.n17058 VCC.n16697 0.0121071
R51052 VCC.n16760 VCC.n16758 0.0121071
R51053 VCC.n16828 VCC.n16827 0.0121071
R51054 VCC.n17313 VCC.n17310 0.0121071
R51055 VCC.n17432 VCC.n17431 0.0121071
R51056 VCC.n17421 VCC.n17248 0.0121071
R51057 VCC.n17444 VCC.n17437 0.0121071
R51058 VCC.n17442 VCC.n17439 0.0121071
R51059 VCC.n17441 VCC.n17440 0.0121071
R51060 VCC.n17191 VCC.n17188 0.0121071
R51061 VCC.n199 VCC.n185 0.0112143
R51062 VCC.n303 VCC.n135 0.0112143
R51063 VCC.n311 VCC.n310 0.0112143
R51064 VCC.n198 VCC.n186 0.0112143
R51065 VCC.n302 VCC.n301 0.0112143
R51066 VCC.n300 VCC.n136 0.0112143
R51067 VCC.n324 VCC.n323 0.0112143
R51068 VCC.n439 VCC.n438 0.0112143
R51069 VCC.n330 VCC.n329 0.0112143
R51070 VCC.n322 VCC.n321 0.0112143
R51071 VCC.n437 VCC.n72 0.0112143
R51072 VCC.n453 VCC.n452 0.0112143
R51073 VCC.n467 VCC.n59 0.0112143
R51074 VCC.n533 VCC.n532 0.0112143
R51075 VCC.n466 VCC.n465 0.0112143
R51076 VCC.n751 VCC.n737 0.0112143
R51077 VCC.n855 VCC.n687 0.0112143
R51078 VCC.n863 VCC.n862 0.0112143
R51079 VCC.n750 VCC.n738 0.0112143
R51080 VCC.n854 VCC.n853 0.0112143
R51081 VCC.n852 VCC.n688 0.0112143
R51082 VCC.n876 VCC.n875 0.0112143
R51083 VCC.n991 VCC.n990 0.0112143
R51084 VCC.n882 VCC.n881 0.0112143
R51085 VCC.n874 VCC.n873 0.0112143
R51086 VCC.n989 VCC.n624 0.0112143
R51087 VCC.n1005 VCC.n1004 0.0112143
R51088 VCC.n1019 VCC.n611 0.0112143
R51089 VCC.n1085 VCC.n1084 0.0112143
R51090 VCC.n1018 VCC.n1017 0.0112143
R51091 VCC.n1563 VCC.n1562 0.0112143
R51092 VCC.n1576 VCC.n1575 0.0112143
R51093 VCC.n1647 VCC.n1118 0.0112143
R51094 VCC.n1574 VCC.n1167 0.0112143
R51095 VCC.n1433 VCC.n1432 0.0112143
R51096 VCC.n1549 VCC.n1548 0.0112143
R51097 VCC.n1439 VCC.n1438 0.0112143
R51098 VCC.n1431 VCC.n1429 0.0112143
R51099 VCC.n1547 VCC.n1181 0.0112143
R51100 VCC.n1309 VCC.n1295 0.0112143
R51101 VCC.n1413 VCC.n1245 0.0112143
R51102 VCC.n1421 VCC.n1420 0.0112143
R51103 VCC.n1308 VCC.n1296 0.0112143
R51104 VCC.n1412 VCC.n1411 0.0112143
R51105 VCC.n1410 VCC.n1246 0.0112143
R51106 VCC.n1860 VCC.n1846 0.0112143
R51107 VCC.n1964 VCC.n1796 0.0112143
R51108 VCC.n1972 VCC.n1971 0.0112143
R51109 VCC.n1859 VCC.n1847 0.0112143
R51110 VCC.n1963 VCC.n1962 0.0112143
R51111 VCC.n1961 VCC.n1797 0.0112143
R51112 VCC.n1985 VCC.n1984 0.0112143
R51113 VCC.n2100 VCC.n2099 0.0112143
R51114 VCC.n1991 VCC.n1990 0.0112143
R51115 VCC.n1983 VCC.n1982 0.0112143
R51116 VCC.n2098 VCC.n1733 0.0112143
R51117 VCC.n2114 VCC.n2113 0.0112143
R51118 VCC.n2128 VCC.n1720 0.0112143
R51119 VCC.n2194 VCC.n2193 0.0112143
R51120 VCC.n2127 VCC.n2126 0.0112143
R51121 VCC.n2672 VCC.n2671 0.0112143
R51122 VCC.n2685 VCC.n2684 0.0112143
R51123 VCC.n2756 VCC.n2227 0.0112143
R51124 VCC.n2683 VCC.n2276 0.0112143
R51125 VCC.n2542 VCC.n2541 0.0112143
R51126 VCC.n2658 VCC.n2657 0.0112143
R51127 VCC.n2548 VCC.n2547 0.0112143
R51128 VCC.n2540 VCC.n2538 0.0112143
R51129 VCC.n2656 VCC.n2290 0.0112143
R51130 VCC.n2418 VCC.n2404 0.0112143
R51131 VCC.n2522 VCC.n2354 0.0112143
R51132 VCC.n2530 VCC.n2529 0.0112143
R51133 VCC.n2417 VCC.n2405 0.0112143
R51134 VCC.n2521 VCC.n2520 0.0112143
R51135 VCC.n2519 VCC.n2355 0.0112143
R51136 VCC.n2969 VCC.n2955 0.0112143
R51137 VCC.n3073 VCC.n2905 0.0112143
R51138 VCC.n3081 VCC.n3080 0.0112143
R51139 VCC.n2968 VCC.n2956 0.0112143
R51140 VCC.n3072 VCC.n3071 0.0112143
R51141 VCC.n3070 VCC.n2906 0.0112143
R51142 VCC.n3094 VCC.n3093 0.0112143
R51143 VCC.n3209 VCC.n3208 0.0112143
R51144 VCC.n3100 VCC.n3099 0.0112143
R51145 VCC.n3092 VCC.n3091 0.0112143
R51146 VCC.n3207 VCC.n2842 0.0112143
R51147 VCC.n3223 VCC.n3222 0.0112143
R51148 VCC.n3237 VCC.n2829 0.0112143
R51149 VCC.n3303 VCC.n3302 0.0112143
R51150 VCC.n3236 VCC.n3235 0.0112143
R51151 VCC.n3781 VCC.n3780 0.0112143
R51152 VCC.n3794 VCC.n3793 0.0112143
R51153 VCC.n3865 VCC.n3336 0.0112143
R51154 VCC.n3792 VCC.n3385 0.0112143
R51155 VCC.n3651 VCC.n3650 0.0112143
R51156 VCC.n3767 VCC.n3766 0.0112143
R51157 VCC.n3657 VCC.n3656 0.0112143
R51158 VCC.n3649 VCC.n3647 0.0112143
R51159 VCC.n3765 VCC.n3399 0.0112143
R51160 VCC.n3527 VCC.n3513 0.0112143
R51161 VCC.n3631 VCC.n3463 0.0112143
R51162 VCC.n3639 VCC.n3638 0.0112143
R51163 VCC.n3526 VCC.n3514 0.0112143
R51164 VCC.n3630 VCC.n3629 0.0112143
R51165 VCC.n3628 VCC.n3464 0.0112143
R51166 VCC.n4078 VCC.n4064 0.0112143
R51167 VCC.n4182 VCC.n4014 0.0112143
R51168 VCC.n4190 VCC.n4189 0.0112143
R51169 VCC.n4077 VCC.n4065 0.0112143
R51170 VCC.n4181 VCC.n4180 0.0112143
R51171 VCC.n4179 VCC.n4015 0.0112143
R51172 VCC.n4203 VCC.n4202 0.0112143
R51173 VCC.n4318 VCC.n4317 0.0112143
R51174 VCC.n4209 VCC.n4208 0.0112143
R51175 VCC.n4201 VCC.n4200 0.0112143
R51176 VCC.n4316 VCC.n3951 0.0112143
R51177 VCC.n4332 VCC.n4331 0.0112143
R51178 VCC.n4346 VCC.n3938 0.0112143
R51179 VCC.n4412 VCC.n4411 0.0112143
R51180 VCC.n4345 VCC.n4344 0.0112143
R51181 VCC.n4890 VCC.n4889 0.0112143
R51182 VCC.n4903 VCC.n4902 0.0112143
R51183 VCC.n4974 VCC.n4445 0.0112143
R51184 VCC.n4901 VCC.n4494 0.0112143
R51185 VCC.n4760 VCC.n4759 0.0112143
R51186 VCC.n4876 VCC.n4875 0.0112143
R51187 VCC.n4766 VCC.n4765 0.0112143
R51188 VCC.n4758 VCC.n4756 0.0112143
R51189 VCC.n4874 VCC.n4508 0.0112143
R51190 VCC.n4636 VCC.n4622 0.0112143
R51191 VCC.n4740 VCC.n4572 0.0112143
R51192 VCC.n4748 VCC.n4747 0.0112143
R51193 VCC.n4635 VCC.n4623 0.0112143
R51194 VCC.n4739 VCC.n4738 0.0112143
R51195 VCC.n4737 VCC.n4573 0.0112143
R51196 VCC.n5187 VCC.n5173 0.0112143
R51197 VCC.n5291 VCC.n5123 0.0112143
R51198 VCC.n5299 VCC.n5298 0.0112143
R51199 VCC.n5186 VCC.n5174 0.0112143
R51200 VCC.n5290 VCC.n5289 0.0112143
R51201 VCC.n5288 VCC.n5124 0.0112143
R51202 VCC.n5312 VCC.n5311 0.0112143
R51203 VCC.n5427 VCC.n5426 0.0112143
R51204 VCC.n5318 VCC.n5317 0.0112143
R51205 VCC.n5310 VCC.n5309 0.0112143
R51206 VCC.n5425 VCC.n5060 0.0112143
R51207 VCC.n5441 VCC.n5440 0.0112143
R51208 VCC.n5455 VCC.n5047 0.0112143
R51209 VCC.n5521 VCC.n5520 0.0112143
R51210 VCC.n5454 VCC.n5453 0.0112143
R51211 VCC.n5999 VCC.n5998 0.0112143
R51212 VCC.n6012 VCC.n6011 0.0112143
R51213 VCC.n6083 VCC.n5554 0.0112143
R51214 VCC.n6010 VCC.n5603 0.0112143
R51215 VCC.n5869 VCC.n5868 0.0112143
R51216 VCC.n5985 VCC.n5984 0.0112143
R51217 VCC.n5875 VCC.n5874 0.0112143
R51218 VCC.n5867 VCC.n5865 0.0112143
R51219 VCC.n5983 VCC.n5617 0.0112143
R51220 VCC.n5745 VCC.n5731 0.0112143
R51221 VCC.n5849 VCC.n5681 0.0112143
R51222 VCC.n5857 VCC.n5856 0.0112143
R51223 VCC.n5744 VCC.n5732 0.0112143
R51224 VCC.n5848 VCC.n5847 0.0112143
R51225 VCC.n5846 VCC.n5682 0.0112143
R51226 VCC.n6296 VCC.n6282 0.0112143
R51227 VCC.n6400 VCC.n6232 0.0112143
R51228 VCC.n6408 VCC.n6407 0.0112143
R51229 VCC.n6295 VCC.n6283 0.0112143
R51230 VCC.n6399 VCC.n6398 0.0112143
R51231 VCC.n6397 VCC.n6233 0.0112143
R51232 VCC.n6421 VCC.n6420 0.0112143
R51233 VCC.n6536 VCC.n6535 0.0112143
R51234 VCC.n6427 VCC.n6426 0.0112143
R51235 VCC.n6419 VCC.n6418 0.0112143
R51236 VCC.n6534 VCC.n6169 0.0112143
R51237 VCC.n6550 VCC.n6549 0.0112143
R51238 VCC.n6564 VCC.n6156 0.0112143
R51239 VCC.n6630 VCC.n6629 0.0112143
R51240 VCC.n6563 VCC.n6562 0.0112143
R51241 VCC.n7108 VCC.n7107 0.0112143
R51242 VCC.n7121 VCC.n7120 0.0112143
R51243 VCC.n7192 VCC.n6663 0.0112143
R51244 VCC.n7119 VCC.n6712 0.0112143
R51245 VCC.n6978 VCC.n6977 0.0112143
R51246 VCC.n7094 VCC.n7093 0.0112143
R51247 VCC.n6984 VCC.n6983 0.0112143
R51248 VCC.n6976 VCC.n6974 0.0112143
R51249 VCC.n7092 VCC.n6726 0.0112143
R51250 VCC.n6854 VCC.n6840 0.0112143
R51251 VCC.n6958 VCC.n6790 0.0112143
R51252 VCC.n6966 VCC.n6965 0.0112143
R51253 VCC.n6853 VCC.n6841 0.0112143
R51254 VCC.n6957 VCC.n6956 0.0112143
R51255 VCC.n6955 VCC.n6791 0.0112143
R51256 VCC.n7405 VCC.n7391 0.0112143
R51257 VCC.n7509 VCC.n7341 0.0112143
R51258 VCC.n7517 VCC.n7516 0.0112143
R51259 VCC.n7404 VCC.n7392 0.0112143
R51260 VCC.n7508 VCC.n7507 0.0112143
R51261 VCC.n7506 VCC.n7342 0.0112143
R51262 VCC.n7530 VCC.n7529 0.0112143
R51263 VCC.n7645 VCC.n7644 0.0112143
R51264 VCC.n7536 VCC.n7535 0.0112143
R51265 VCC.n7528 VCC.n7527 0.0112143
R51266 VCC.n7643 VCC.n7278 0.0112143
R51267 VCC.n7659 VCC.n7658 0.0112143
R51268 VCC.n7673 VCC.n7265 0.0112143
R51269 VCC.n7739 VCC.n7738 0.0112143
R51270 VCC.n7672 VCC.n7671 0.0112143
R51271 VCC.n8217 VCC.n8216 0.0112143
R51272 VCC.n8230 VCC.n8229 0.0112143
R51273 VCC.n8301 VCC.n7772 0.0112143
R51274 VCC.n8228 VCC.n7821 0.0112143
R51275 VCC.n8087 VCC.n8086 0.0112143
R51276 VCC.n8203 VCC.n8202 0.0112143
R51277 VCC.n8093 VCC.n8092 0.0112143
R51278 VCC.n8085 VCC.n8083 0.0112143
R51279 VCC.n8201 VCC.n7835 0.0112143
R51280 VCC.n7963 VCC.n7949 0.0112143
R51281 VCC.n8067 VCC.n7899 0.0112143
R51282 VCC.n8075 VCC.n8074 0.0112143
R51283 VCC.n7962 VCC.n7950 0.0112143
R51284 VCC.n8066 VCC.n8065 0.0112143
R51285 VCC.n8064 VCC.n7900 0.0112143
R51286 VCC.n8639 VCC.n8638 0.0112143
R51287 VCC.n8754 VCC.n8753 0.0112143
R51288 VCC.n8645 VCC.n8644 0.0112143
R51289 VCC.n8637 VCC.n8636 0.0112143
R51290 VCC.n8752 VCC.n8387 0.0112143
R51291 VCC.n8768 VCC.n8767 0.0112143
R51292 VCC.n8782 VCC.n8374 0.0112143
R51293 VCC.n8848 VCC.n8847 0.0112143
R51294 VCC.n8781 VCC.n8780 0.0112143
R51295 VCC.n8514 VCC.n8500 0.0112143
R51296 VCC.n8618 VCC.n8450 0.0112143
R51297 VCC.n8626 VCC.n8625 0.0112143
R51298 VCC.n8513 VCC.n8501 0.0112143
R51299 VCC.n8617 VCC.n8616 0.0112143
R51300 VCC.n8615 VCC.n8451 0.0112143
R51301 VCC.n9326 VCC.n9325 0.0112143
R51302 VCC.n9339 VCC.n9338 0.0112143
R51303 VCC.n9410 VCC.n8881 0.0112143
R51304 VCC.n9337 VCC.n8930 0.0112143
R51305 VCC.n9196 VCC.n9195 0.0112143
R51306 VCC.n9312 VCC.n9311 0.0112143
R51307 VCC.n9202 VCC.n9201 0.0112143
R51308 VCC.n9194 VCC.n9192 0.0112143
R51309 VCC.n9310 VCC.n8944 0.0112143
R51310 VCC.n9072 VCC.n9058 0.0112143
R51311 VCC.n9176 VCC.n9008 0.0112143
R51312 VCC.n9184 VCC.n9183 0.0112143
R51313 VCC.n9071 VCC.n9059 0.0112143
R51314 VCC.n9175 VCC.n9174 0.0112143
R51315 VCC.n9173 VCC.n9009 0.0112143
R51316 VCC.n9623 VCC.n9609 0.0112143
R51317 VCC.n9727 VCC.n9559 0.0112143
R51318 VCC.n9735 VCC.n9734 0.0112143
R51319 VCC.n9622 VCC.n9610 0.0112143
R51320 VCC.n9726 VCC.n9725 0.0112143
R51321 VCC.n9724 VCC.n9560 0.0112143
R51322 VCC.n9748 VCC.n9747 0.0112143
R51323 VCC.n9863 VCC.n9862 0.0112143
R51324 VCC.n9754 VCC.n9753 0.0112143
R51325 VCC.n9746 VCC.n9745 0.0112143
R51326 VCC.n9861 VCC.n9496 0.0112143
R51327 VCC.n9877 VCC.n9876 0.0112143
R51328 VCC.n9891 VCC.n9483 0.0112143
R51329 VCC.n9957 VCC.n9956 0.0112143
R51330 VCC.n9890 VCC.n9889 0.0112143
R51331 VCC.n10434 VCC.n10433 0.0112143
R51332 VCC.n10447 VCC.n10446 0.0112143
R51333 VCC.n10518 VCC.n9989 0.0112143
R51334 VCC.n10445 VCC.n10038 0.0112143
R51335 VCC.n10304 VCC.n10303 0.0112143
R51336 VCC.n10420 VCC.n10419 0.0112143
R51337 VCC.n10310 VCC.n10309 0.0112143
R51338 VCC.n10302 VCC.n10300 0.0112143
R51339 VCC.n10418 VCC.n10052 0.0112143
R51340 VCC.n10180 VCC.n10166 0.0112143
R51341 VCC.n10284 VCC.n10116 0.0112143
R51342 VCC.n10292 VCC.n10291 0.0112143
R51343 VCC.n10179 VCC.n10167 0.0112143
R51344 VCC.n10283 VCC.n10282 0.0112143
R51345 VCC.n10281 VCC.n10117 0.0112143
R51346 VCC.n10730 VCC.n10716 0.0112143
R51347 VCC.n10834 VCC.n10666 0.0112143
R51348 VCC.n10842 VCC.n10841 0.0112143
R51349 VCC.n10729 VCC.n10717 0.0112143
R51350 VCC.n10833 VCC.n10832 0.0112143
R51351 VCC.n10831 VCC.n10667 0.0112143
R51352 VCC.n10855 VCC.n10854 0.0112143
R51353 VCC.n10970 VCC.n10969 0.0112143
R51354 VCC.n10861 VCC.n10860 0.0112143
R51355 VCC.n10853 VCC.n10852 0.0112143
R51356 VCC.n10968 VCC.n10603 0.0112143
R51357 VCC.n10984 VCC.n10983 0.0112143
R51358 VCC.n10998 VCC.n10590 0.0112143
R51359 VCC.n11064 VCC.n11063 0.0112143
R51360 VCC.n10997 VCC.n10996 0.0112143
R51361 VCC.n11541 VCC.n11540 0.0112143
R51362 VCC.n11554 VCC.n11553 0.0112143
R51363 VCC.n11625 VCC.n11096 0.0112143
R51364 VCC.n11552 VCC.n11145 0.0112143
R51365 VCC.n11411 VCC.n11410 0.0112143
R51366 VCC.n11527 VCC.n11526 0.0112143
R51367 VCC.n11417 VCC.n11416 0.0112143
R51368 VCC.n11409 VCC.n11407 0.0112143
R51369 VCC.n11525 VCC.n11159 0.0112143
R51370 VCC.n11287 VCC.n11273 0.0112143
R51371 VCC.n11391 VCC.n11223 0.0112143
R51372 VCC.n11399 VCC.n11398 0.0112143
R51373 VCC.n11286 VCC.n11274 0.0112143
R51374 VCC.n11390 VCC.n11389 0.0112143
R51375 VCC.n11388 VCC.n11224 0.0112143
R51376 VCC.n11837 VCC.n11823 0.0112143
R51377 VCC.n11941 VCC.n11773 0.0112143
R51378 VCC.n11949 VCC.n11948 0.0112143
R51379 VCC.n11836 VCC.n11824 0.0112143
R51380 VCC.n11940 VCC.n11939 0.0112143
R51381 VCC.n11938 VCC.n11774 0.0112143
R51382 VCC.n11962 VCC.n11961 0.0112143
R51383 VCC.n12077 VCC.n12076 0.0112143
R51384 VCC.n11968 VCC.n11967 0.0112143
R51385 VCC.n11960 VCC.n11959 0.0112143
R51386 VCC.n12075 VCC.n11710 0.0112143
R51387 VCC.n12091 VCC.n12090 0.0112143
R51388 VCC.n12105 VCC.n11697 0.0112143
R51389 VCC.n12171 VCC.n12170 0.0112143
R51390 VCC.n12104 VCC.n12103 0.0112143
R51391 VCC.n12648 VCC.n12647 0.0112143
R51392 VCC.n12661 VCC.n12660 0.0112143
R51393 VCC.n12732 VCC.n12203 0.0112143
R51394 VCC.n12659 VCC.n12252 0.0112143
R51395 VCC.n12518 VCC.n12517 0.0112143
R51396 VCC.n12634 VCC.n12633 0.0112143
R51397 VCC.n12524 VCC.n12523 0.0112143
R51398 VCC.n12516 VCC.n12514 0.0112143
R51399 VCC.n12632 VCC.n12266 0.0112143
R51400 VCC.n12394 VCC.n12380 0.0112143
R51401 VCC.n12498 VCC.n12330 0.0112143
R51402 VCC.n12506 VCC.n12505 0.0112143
R51403 VCC.n12393 VCC.n12381 0.0112143
R51404 VCC.n12497 VCC.n12496 0.0112143
R51405 VCC.n12495 VCC.n12331 0.0112143
R51406 VCC.n12944 VCC.n12930 0.0112143
R51407 VCC.n13048 VCC.n12880 0.0112143
R51408 VCC.n13056 VCC.n13055 0.0112143
R51409 VCC.n12943 VCC.n12931 0.0112143
R51410 VCC.n13047 VCC.n13046 0.0112143
R51411 VCC.n13045 VCC.n12881 0.0112143
R51412 VCC.n13069 VCC.n13068 0.0112143
R51413 VCC.n13184 VCC.n13183 0.0112143
R51414 VCC.n13075 VCC.n13074 0.0112143
R51415 VCC.n13067 VCC.n13066 0.0112143
R51416 VCC.n13182 VCC.n12817 0.0112143
R51417 VCC.n13198 VCC.n13197 0.0112143
R51418 VCC.n13212 VCC.n12804 0.0112143
R51419 VCC.n13278 VCC.n13277 0.0112143
R51420 VCC.n13211 VCC.n13210 0.0112143
R51421 VCC.n13755 VCC.n13754 0.0112143
R51422 VCC.n13768 VCC.n13767 0.0112143
R51423 VCC.n13839 VCC.n13310 0.0112143
R51424 VCC.n13766 VCC.n13359 0.0112143
R51425 VCC.n13625 VCC.n13624 0.0112143
R51426 VCC.n13741 VCC.n13740 0.0112143
R51427 VCC.n13631 VCC.n13630 0.0112143
R51428 VCC.n13623 VCC.n13621 0.0112143
R51429 VCC.n13739 VCC.n13373 0.0112143
R51430 VCC.n13501 VCC.n13487 0.0112143
R51431 VCC.n13605 VCC.n13437 0.0112143
R51432 VCC.n13613 VCC.n13612 0.0112143
R51433 VCC.n13500 VCC.n13488 0.0112143
R51434 VCC.n13604 VCC.n13603 0.0112143
R51435 VCC.n13602 VCC.n13438 0.0112143
R51436 VCC.n14051 VCC.n14037 0.0112143
R51437 VCC.n14155 VCC.n13987 0.0112143
R51438 VCC.n14163 VCC.n14162 0.0112143
R51439 VCC.n14050 VCC.n14038 0.0112143
R51440 VCC.n14154 VCC.n14153 0.0112143
R51441 VCC.n14152 VCC.n13988 0.0112143
R51442 VCC.n14176 VCC.n14175 0.0112143
R51443 VCC.n14291 VCC.n14290 0.0112143
R51444 VCC.n14182 VCC.n14181 0.0112143
R51445 VCC.n14174 VCC.n14173 0.0112143
R51446 VCC.n14289 VCC.n13924 0.0112143
R51447 VCC.n14305 VCC.n14304 0.0112143
R51448 VCC.n14319 VCC.n13911 0.0112143
R51449 VCC.n14385 VCC.n14384 0.0112143
R51450 VCC.n14318 VCC.n14317 0.0112143
R51451 VCC.n14862 VCC.n14861 0.0112143
R51452 VCC.n14875 VCC.n14874 0.0112143
R51453 VCC.n14946 VCC.n14417 0.0112143
R51454 VCC.n14873 VCC.n14466 0.0112143
R51455 VCC.n14732 VCC.n14731 0.0112143
R51456 VCC.n14848 VCC.n14847 0.0112143
R51457 VCC.n14738 VCC.n14737 0.0112143
R51458 VCC.n14730 VCC.n14728 0.0112143
R51459 VCC.n14846 VCC.n14480 0.0112143
R51460 VCC.n14608 VCC.n14594 0.0112143
R51461 VCC.n14712 VCC.n14544 0.0112143
R51462 VCC.n14720 VCC.n14719 0.0112143
R51463 VCC.n14607 VCC.n14595 0.0112143
R51464 VCC.n14711 VCC.n14710 0.0112143
R51465 VCC.n14709 VCC.n14545 0.0112143
R51466 VCC.n15158 VCC.n15144 0.0112143
R51467 VCC.n15262 VCC.n15094 0.0112143
R51468 VCC.n15270 VCC.n15269 0.0112143
R51469 VCC.n15157 VCC.n15145 0.0112143
R51470 VCC.n15261 VCC.n15260 0.0112143
R51471 VCC.n15259 VCC.n15095 0.0112143
R51472 VCC.n15283 VCC.n15282 0.0112143
R51473 VCC.n15398 VCC.n15397 0.0112143
R51474 VCC.n15289 VCC.n15288 0.0112143
R51475 VCC.n15281 VCC.n15280 0.0112143
R51476 VCC.n15396 VCC.n15031 0.0112143
R51477 VCC.n15412 VCC.n15411 0.0112143
R51478 VCC.n15426 VCC.n15018 0.0112143
R51479 VCC.n15492 VCC.n15491 0.0112143
R51480 VCC.n15425 VCC.n15424 0.0112143
R51481 VCC.n15969 VCC.n15968 0.0112143
R51482 VCC.n15982 VCC.n15981 0.0112143
R51483 VCC.n16053 VCC.n15524 0.0112143
R51484 VCC.n15980 VCC.n15573 0.0112143
R51485 VCC.n15839 VCC.n15838 0.0112143
R51486 VCC.n15955 VCC.n15954 0.0112143
R51487 VCC.n15845 VCC.n15844 0.0112143
R51488 VCC.n15837 VCC.n15835 0.0112143
R51489 VCC.n15953 VCC.n15587 0.0112143
R51490 VCC.n15715 VCC.n15701 0.0112143
R51491 VCC.n15819 VCC.n15651 0.0112143
R51492 VCC.n15827 VCC.n15826 0.0112143
R51493 VCC.n15714 VCC.n15702 0.0112143
R51494 VCC.n15818 VCC.n15817 0.0112143
R51495 VCC.n15816 VCC.n15652 0.0112143
R51496 VCC.n16265 VCC.n16251 0.0112143
R51497 VCC.n16369 VCC.n16201 0.0112143
R51498 VCC.n16377 VCC.n16376 0.0112143
R51499 VCC.n16264 VCC.n16252 0.0112143
R51500 VCC.n16368 VCC.n16367 0.0112143
R51501 VCC.n16366 VCC.n16202 0.0112143
R51502 VCC.n16390 VCC.n16389 0.0112143
R51503 VCC.n16505 VCC.n16504 0.0112143
R51504 VCC.n16396 VCC.n16395 0.0112143
R51505 VCC.n16388 VCC.n16387 0.0112143
R51506 VCC.n16503 VCC.n16138 0.0112143
R51507 VCC.n16519 VCC.n16518 0.0112143
R51508 VCC.n16533 VCC.n16125 0.0112143
R51509 VCC.n16599 VCC.n16598 0.0112143
R51510 VCC.n16532 VCC.n16531 0.0112143
R51511 VCC.n17076 VCC.n17075 0.0112143
R51512 VCC.n17089 VCC.n17088 0.0112143
R51513 VCC.n17160 VCC.n16631 0.0112143
R51514 VCC.n17087 VCC.n16680 0.0112143
R51515 VCC.n16946 VCC.n16945 0.0112143
R51516 VCC.n17062 VCC.n17061 0.0112143
R51517 VCC.n16952 VCC.n16951 0.0112143
R51518 VCC.n16944 VCC.n16942 0.0112143
R51519 VCC.n17060 VCC.n16694 0.0112143
R51520 VCC.n16822 VCC.n16808 0.0112143
R51521 VCC.n16926 VCC.n16758 0.0112143
R51522 VCC.n16934 VCC.n16933 0.0112143
R51523 VCC.n16821 VCC.n16809 0.0112143
R51524 VCC.n16925 VCC.n16924 0.0112143
R51525 VCC.n16923 VCC.n16759 0.0112143
R51526 VCC.n17310 VCC.n17309 0.0112143
R51527 VCC.n17425 VCC.n17424 0.0112143
R51528 VCC.n17316 VCC.n17315 0.0112143
R51529 VCC.n17308 VCC.n17307 0.0112143
R51530 VCC.n17423 VCC.n17245 0.0112143
R51531 VCC.n17439 VCC.n17438 0.0112143
R51532 VCC.n17453 VCC.n17232 0.0112143
R51533 VCC.n17519 VCC.n17518 0.0112143
R51534 VCC.n17452 VCC.n17451 0.0112143
R51535 VCC.n200 VCC.n199 0.0103214
R51536 VCC.n235 VCC.n170 0.0103214
R51537 VCC.n161 VCC.n158 0.0103214
R51538 VCC.n278 VCC.n277 0.0103214
R51539 VCC.n304 VCC.n303 0.0103214
R51540 VCC.n198 VCC.n197 0.0103214
R51541 VCC.n234 VCC.n171 0.0103214
R51542 VCC.n279 VCC.n149 0.0103214
R51543 VCC.n302 VCC.n133 0.0103214
R51544 VCC.n136 VCC.n130 0.0103214
R51545 VCC.n332 VCC.n331 0.0103214
R51546 VCC.n323 VCC.n116 0.0103214
R51547 VCC.n351 VCC.n350 0.0103214
R51548 VCC.n390 VCC.n389 0.0103214
R51549 VCC.n405 VCC.n404 0.0103214
R51550 VCC.n438 VCC.n74 0.0103214
R51551 VCC.n330 VCC.n319 0.0103214
R51552 VCC.n322 VCC.n115 0.0103214
R51553 VCC.n349 VCC.n103 0.0103214
R51554 VCC.n406 VCC.n89 0.0103214
R51555 VCC.n437 VCC.n436 0.0103214
R51556 VCC.n467 VCC.n58 0.0103214
R51557 VCC.n463 VCC.n462 0.0103214
R51558 VCC.n488 VCC.n45 0.0103214
R51559 VCC.n510 VCC.n26 0.0103214
R51560 VCC.n543 VCC.n542 0.0103214
R51561 VCC.n466 VCC.n60 0.0103214
R51562 VCC.n487 VCC.n486 0.0103214
R51563 VCC.n482 VCC.n36 0.0103214
R51564 VCC.n511 VCC.n28 0.0103214
R51565 VCC.n519 VCC.n518 0.0103214
R51566 VCC.n752 VCC.n751 0.0103214
R51567 VCC.n787 VCC.n722 0.0103214
R51568 VCC.n713 VCC.n710 0.0103214
R51569 VCC.n830 VCC.n829 0.0103214
R51570 VCC.n856 VCC.n855 0.0103214
R51571 VCC.n750 VCC.n749 0.0103214
R51572 VCC.n786 VCC.n723 0.0103214
R51573 VCC.n831 VCC.n701 0.0103214
R51574 VCC.n854 VCC.n685 0.0103214
R51575 VCC.n688 VCC.n682 0.0103214
R51576 VCC.n884 VCC.n883 0.0103214
R51577 VCC.n875 VCC.n668 0.0103214
R51578 VCC.n903 VCC.n902 0.0103214
R51579 VCC.n942 VCC.n941 0.0103214
R51580 VCC.n957 VCC.n956 0.0103214
R51581 VCC.n990 VCC.n626 0.0103214
R51582 VCC.n882 VCC.n871 0.0103214
R51583 VCC.n874 VCC.n667 0.0103214
R51584 VCC.n901 VCC.n655 0.0103214
R51585 VCC.n958 VCC.n641 0.0103214
R51586 VCC.n989 VCC.n988 0.0103214
R51587 VCC.n1019 VCC.n610 0.0103214
R51588 VCC.n1015 VCC.n1014 0.0103214
R51589 VCC.n1040 VCC.n597 0.0103214
R51590 VCC.n1062 VCC.n578 0.0103214
R51591 VCC.n1097 VCC.n1096 0.0103214
R51592 VCC.n1018 VCC.n612 0.0103214
R51593 VCC.n1039 VCC.n1038 0.0103214
R51594 VCC.n1034 VCC.n588 0.0103214
R51595 VCC.n1063 VCC.n580 0.0103214
R51596 VCC.n1071 VCC.n1070 0.0103214
R51597 VCC.n1576 VCC.n1166 0.0103214
R51598 VCC.n1169 VCC.n1168 0.0103214
R51599 VCC.n1589 VCC.n1152 0.0103214
R51600 VCC.n1626 VCC.n1625 0.0103214
R51601 VCC.n1642 VCC.n1125 0.0103214
R51602 VCC.n1564 VCC.n1167 0.0103214
R51603 VCC.n1590 VCC.n1153 0.0103214
R51604 VCC.n1606 VCC.n1151 0.0103214
R51605 VCC.n1627 VCC.n1132 0.0103214
R51606 VCC.n1137 VCC.n1129 0.0103214
R51607 VCC.n1441 VCC.n1235 0.0103214
R51608 VCC.n1432 VCC.n1225 0.0103214
R51609 VCC.n1460 VCC.n1459 0.0103214
R51610 VCC.n1499 VCC.n1498 0.0103214
R51611 VCC.n1514 VCC.n1513 0.0103214
R51612 VCC.n1548 VCC.n1183 0.0103214
R51613 VCC.n1440 VCC.n1439 0.0103214
R51614 VCC.n1431 VCC.n1224 0.0103214
R51615 VCC.n1458 VCC.n1212 0.0103214
R51616 VCC.n1515 VCC.n1198 0.0103214
R51617 VCC.n1547 VCC.n1546 0.0103214
R51618 VCC.n1310 VCC.n1309 0.0103214
R51619 VCC.n1345 VCC.n1280 0.0103214
R51620 VCC.n1271 VCC.n1268 0.0103214
R51621 VCC.n1388 VCC.n1387 0.0103214
R51622 VCC.n1414 VCC.n1413 0.0103214
R51623 VCC.n1308 VCC.n1307 0.0103214
R51624 VCC.n1344 VCC.n1281 0.0103214
R51625 VCC.n1389 VCC.n1259 0.0103214
R51626 VCC.n1412 VCC.n1243 0.0103214
R51627 VCC.n1246 VCC.n1240 0.0103214
R51628 VCC.n1861 VCC.n1860 0.0103214
R51629 VCC.n1896 VCC.n1831 0.0103214
R51630 VCC.n1822 VCC.n1819 0.0103214
R51631 VCC.n1939 VCC.n1938 0.0103214
R51632 VCC.n1965 VCC.n1964 0.0103214
R51633 VCC.n1859 VCC.n1858 0.0103214
R51634 VCC.n1895 VCC.n1832 0.0103214
R51635 VCC.n1940 VCC.n1810 0.0103214
R51636 VCC.n1963 VCC.n1794 0.0103214
R51637 VCC.n1797 VCC.n1791 0.0103214
R51638 VCC.n1993 VCC.n1992 0.0103214
R51639 VCC.n1984 VCC.n1777 0.0103214
R51640 VCC.n2012 VCC.n2011 0.0103214
R51641 VCC.n2051 VCC.n2050 0.0103214
R51642 VCC.n2066 VCC.n2065 0.0103214
R51643 VCC.n2099 VCC.n1735 0.0103214
R51644 VCC.n1991 VCC.n1980 0.0103214
R51645 VCC.n1983 VCC.n1776 0.0103214
R51646 VCC.n2010 VCC.n1764 0.0103214
R51647 VCC.n2067 VCC.n1750 0.0103214
R51648 VCC.n2098 VCC.n2097 0.0103214
R51649 VCC.n2128 VCC.n1719 0.0103214
R51650 VCC.n2124 VCC.n2123 0.0103214
R51651 VCC.n2149 VCC.n1706 0.0103214
R51652 VCC.n2171 VCC.n1687 0.0103214
R51653 VCC.n2206 VCC.n2205 0.0103214
R51654 VCC.n2127 VCC.n1721 0.0103214
R51655 VCC.n2148 VCC.n2147 0.0103214
R51656 VCC.n2143 VCC.n1697 0.0103214
R51657 VCC.n2172 VCC.n1689 0.0103214
R51658 VCC.n2180 VCC.n2179 0.0103214
R51659 VCC.n2685 VCC.n2275 0.0103214
R51660 VCC.n2278 VCC.n2277 0.0103214
R51661 VCC.n2698 VCC.n2261 0.0103214
R51662 VCC.n2735 VCC.n2734 0.0103214
R51663 VCC.n2751 VCC.n2234 0.0103214
R51664 VCC.n2673 VCC.n2276 0.0103214
R51665 VCC.n2699 VCC.n2262 0.0103214
R51666 VCC.n2715 VCC.n2260 0.0103214
R51667 VCC.n2736 VCC.n2241 0.0103214
R51668 VCC.n2246 VCC.n2238 0.0103214
R51669 VCC.n2550 VCC.n2344 0.0103214
R51670 VCC.n2541 VCC.n2334 0.0103214
R51671 VCC.n2569 VCC.n2568 0.0103214
R51672 VCC.n2608 VCC.n2607 0.0103214
R51673 VCC.n2623 VCC.n2622 0.0103214
R51674 VCC.n2657 VCC.n2292 0.0103214
R51675 VCC.n2549 VCC.n2548 0.0103214
R51676 VCC.n2540 VCC.n2333 0.0103214
R51677 VCC.n2567 VCC.n2321 0.0103214
R51678 VCC.n2624 VCC.n2307 0.0103214
R51679 VCC.n2656 VCC.n2655 0.0103214
R51680 VCC.n2419 VCC.n2418 0.0103214
R51681 VCC.n2454 VCC.n2389 0.0103214
R51682 VCC.n2380 VCC.n2377 0.0103214
R51683 VCC.n2497 VCC.n2496 0.0103214
R51684 VCC.n2523 VCC.n2522 0.0103214
R51685 VCC.n2417 VCC.n2416 0.0103214
R51686 VCC.n2453 VCC.n2390 0.0103214
R51687 VCC.n2498 VCC.n2368 0.0103214
R51688 VCC.n2521 VCC.n2352 0.0103214
R51689 VCC.n2355 VCC.n2349 0.0103214
R51690 VCC.n2970 VCC.n2969 0.0103214
R51691 VCC.n3005 VCC.n2940 0.0103214
R51692 VCC.n2931 VCC.n2928 0.0103214
R51693 VCC.n3048 VCC.n3047 0.0103214
R51694 VCC.n3074 VCC.n3073 0.0103214
R51695 VCC.n2968 VCC.n2967 0.0103214
R51696 VCC.n3004 VCC.n2941 0.0103214
R51697 VCC.n3049 VCC.n2919 0.0103214
R51698 VCC.n3072 VCC.n2903 0.0103214
R51699 VCC.n2906 VCC.n2900 0.0103214
R51700 VCC.n3102 VCC.n3101 0.0103214
R51701 VCC.n3093 VCC.n2886 0.0103214
R51702 VCC.n3121 VCC.n3120 0.0103214
R51703 VCC.n3160 VCC.n3159 0.0103214
R51704 VCC.n3175 VCC.n3174 0.0103214
R51705 VCC.n3208 VCC.n2844 0.0103214
R51706 VCC.n3100 VCC.n3089 0.0103214
R51707 VCC.n3092 VCC.n2885 0.0103214
R51708 VCC.n3119 VCC.n2873 0.0103214
R51709 VCC.n3176 VCC.n2859 0.0103214
R51710 VCC.n3207 VCC.n3206 0.0103214
R51711 VCC.n3237 VCC.n2828 0.0103214
R51712 VCC.n3233 VCC.n3232 0.0103214
R51713 VCC.n3258 VCC.n2815 0.0103214
R51714 VCC.n3280 VCC.n2796 0.0103214
R51715 VCC.n3315 VCC.n3314 0.0103214
R51716 VCC.n3236 VCC.n2830 0.0103214
R51717 VCC.n3257 VCC.n3256 0.0103214
R51718 VCC.n3252 VCC.n2806 0.0103214
R51719 VCC.n3281 VCC.n2798 0.0103214
R51720 VCC.n3289 VCC.n3288 0.0103214
R51721 VCC.n3794 VCC.n3384 0.0103214
R51722 VCC.n3387 VCC.n3386 0.0103214
R51723 VCC.n3807 VCC.n3370 0.0103214
R51724 VCC.n3844 VCC.n3843 0.0103214
R51725 VCC.n3860 VCC.n3343 0.0103214
R51726 VCC.n3782 VCC.n3385 0.0103214
R51727 VCC.n3808 VCC.n3371 0.0103214
R51728 VCC.n3824 VCC.n3369 0.0103214
R51729 VCC.n3845 VCC.n3350 0.0103214
R51730 VCC.n3355 VCC.n3347 0.0103214
R51731 VCC.n3659 VCC.n3453 0.0103214
R51732 VCC.n3650 VCC.n3443 0.0103214
R51733 VCC.n3678 VCC.n3677 0.0103214
R51734 VCC.n3717 VCC.n3716 0.0103214
R51735 VCC.n3732 VCC.n3731 0.0103214
R51736 VCC.n3766 VCC.n3401 0.0103214
R51737 VCC.n3658 VCC.n3657 0.0103214
R51738 VCC.n3649 VCC.n3442 0.0103214
R51739 VCC.n3676 VCC.n3430 0.0103214
R51740 VCC.n3733 VCC.n3416 0.0103214
R51741 VCC.n3765 VCC.n3764 0.0103214
R51742 VCC.n3528 VCC.n3527 0.0103214
R51743 VCC.n3563 VCC.n3498 0.0103214
R51744 VCC.n3489 VCC.n3486 0.0103214
R51745 VCC.n3606 VCC.n3605 0.0103214
R51746 VCC.n3632 VCC.n3631 0.0103214
R51747 VCC.n3526 VCC.n3525 0.0103214
R51748 VCC.n3562 VCC.n3499 0.0103214
R51749 VCC.n3607 VCC.n3477 0.0103214
R51750 VCC.n3630 VCC.n3461 0.0103214
R51751 VCC.n3464 VCC.n3458 0.0103214
R51752 VCC.n4079 VCC.n4078 0.0103214
R51753 VCC.n4114 VCC.n4049 0.0103214
R51754 VCC.n4040 VCC.n4037 0.0103214
R51755 VCC.n4157 VCC.n4156 0.0103214
R51756 VCC.n4183 VCC.n4182 0.0103214
R51757 VCC.n4077 VCC.n4076 0.0103214
R51758 VCC.n4113 VCC.n4050 0.0103214
R51759 VCC.n4158 VCC.n4028 0.0103214
R51760 VCC.n4181 VCC.n4012 0.0103214
R51761 VCC.n4015 VCC.n4009 0.0103214
R51762 VCC.n4211 VCC.n4210 0.0103214
R51763 VCC.n4202 VCC.n3995 0.0103214
R51764 VCC.n4230 VCC.n4229 0.0103214
R51765 VCC.n4269 VCC.n4268 0.0103214
R51766 VCC.n4284 VCC.n4283 0.0103214
R51767 VCC.n4317 VCC.n3953 0.0103214
R51768 VCC.n4209 VCC.n4198 0.0103214
R51769 VCC.n4201 VCC.n3994 0.0103214
R51770 VCC.n4228 VCC.n3982 0.0103214
R51771 VCC.n4285 VCC.n3968 0.0103214
R51772 VCC.n4316 VCC.n4315 0.0103214
R51773 VCC.n4346 VCC.n3937 0.0103214
R51774 VCC.n4342 VCC.n4341 0.0103214
R51775 VCC.n4367 VCC.n3924 0.0103214
R51776 VCC.n4389 VCC.n3905 0.0103214
R51777 VCC.n4424 VCC.n4423 0.0103214
R51778 VCC.n4345 VCC.n3939 0.0103214
R51779 VCC.n4366 VCC.n4365 0.0103214
R51780 VCC.n4361 VCC.n3915 0.0103214
R51781 VCC.n4390 VCC.n3907 0.0103214
R51782 VCC.n4398 VCC.n4397 0.0103214
R51783 VCC.n4903 VCC.n4493 0.0103214
R51784 VCC.n4496 VCC.n4495 0.0103214
R51785 VCC.n4916 VCC.n4479 0.0103214
R51786 VCC.n4953 VCC.n4952 0.0103214
R51787 VCC.n4969 VCC.n4452 0.0103214
R51788 VCC.n4891 VCC.n4494 0.0103214
R51789 VCC.n4917 VCC.n4480 0.0103214
R51790 VCC.n4933 VCC.n4478 0.0103214
R51791 VCC.n4954 VCC.n4459 0.0103214
R51792 VCC.n4464 VCC.n4456 0.0103214
R51793 VCC.n4768 VCC.n4562 0.0103214
R51794 VCC.n4759 VCC.n4552 0.0103214
R51795 VCC.n4787 VCC.n4786 0.0103214
R51796 VCC.n4826 VCC.n4825 0.0103214
R51797 VCC.n4841 VCC.n4840 0.0103214
R51798 VCC.n4875 VCC.n4510 0.0103214
R51799 VCC.n4767 VCC.n4766 0.0103214
R51800 VCC.n4758 VCC.n4551 0.0103214
R51801 VCC.n4785 VCC.n4539 0.0103214
R51802 VCC.n4842 VCC.n4525 0.0103214
R51803 VCC.n4874 VCC.n4873 0.0103214
R51804 VCC.n4637 VCC.n4636 0.0103214
R51805 VCC.n4672 VCC.n4607 0.0103214
R51806 VCC.n4598 VCC.n4595 0.0103214
R51807 VCC.n4715 VCC.n4714 0.0103214
R51808 VCC.n4741 VCC.n4740 0.0103214
R51809 VCC.n4635 VCC.n4634 0.0103214
R51810 VCC.n4671 VCC.n4608 0.0103214
R51811 VCC.n4716 VCC.n4586 0.0103214
R51812 VCC.n4739 VCC.n4570 0.0103214
R51813 VCC.n4573 VCC.n4567 0.0103214
R51814 VCC.n5188 VCC.n5187 0.0103214
R51815 VCC.n5223 VCC.n5158 0.0103214
R51816 VCC.n5149 VCC.n5146 0.0103214
R51817 VCC.n5266 VCC.n5265 0.0103214
R51818 VCC.n5292 VCC.n5291 0.0103214
R51819 VCC.n5186 VCC.n5185 0.0103214
R51820 VCC.n5222 VCC.n5159 0.0103214
R51821 VCC.n5267 VCC.n5137 0.0103214
R51822 VCC.n5290 VCC.n5121 0.0103214
R51823 VCC.n5124 VCC.n5118 0.0103214
R51824 VCC.n5320 VCC.n5319 0.0103214
R51825 VCC.n5311 VCC.n5104 0.0103214
R51826 VCC.n5339 VCC.n5338 0.0103214
R51827 VCC.n5378 VCC.n5377 0.0103214
R51828 VCC.n5393 VCC.n5392 0.0103214
R51829 VCC.n5426 VCC.n5062 0.0103214
R51830 VCC.n5318 VCC.n5307 0.0103214
R51831 VCC.n5310 VCC.n5103 0.0103214
R51832 VCC.n5337 VCC.n5091 0.0103214
R51833 VCC.n5394 VCC.n5077 0.0103214
R51834 VCC.n5425 VCC.n5424 0.0103214
R51835 VCC.n5455 VCC.n5046 0.0103214
R51836 VCC.n5451 VCC.n5450 0.0103214
R51837 VCC.n5476 VCC.n5033 0.0103214
R51838 VCC.n5498 VCC.n5014 0.0103214
R51839 VCC.n5533 VCC.n5532 0.0103214
R51840 VCC.n5454 VCC.n5048 0.0103214
R51841 VCC.n5475 VCC.n5474 0.0103214
R51842 VCC.n5470 VCC.n5024 0.0103214
R51843 VCC.n5499 VCC.n5016 0.0103214
R51844 VCC.n5507 VCC.n5506 0.0103214
R51845 VCC.n6012 VCC.n5602 0.0103214
R51846 VCC.n5605 VCC.n5604 0.0103214
R51847 VCC.n6025 VCC.n5588 0.0103214
R51848 VCC.n6062 VCC.n6061 0.0103214
R51849 VCC.n6078 VCC.n5561 0.0103214
R51850 VCC.n6000 VCC.n5603 0.0103214
R51851 VCC.n6026 VCC.n5589 0.0103214
R51852 VCC.n6042 VCC.n5587 0.0103214
R51853 VCC.n6063 VCC.n5568 0.0103214
R51854 VCC.n5573 VCC.n5565 0.0103214
R51855 VCC.n5877 VCC.n5671 0.0103214
R51856 VCC.n5868 VCC.n5661 0.0103214
R51857 VCC.n5896 VCC.n5895 0.0103214
R51858 VCC.n5935 VCC.n5934 0.0103214
R51859 VCC.n5950 VCC.n5949 0.0103214
R51860 VCC.n5984 VCC.n5619 0.0103214
R51861 VCC.n5876 VCC.n5875 0.0103214
R51862 VCC.n5867 VCC.n5660 0.0103214
R51863 VCC.n5894 VCC.n5648 0.0103214
R51864 VCC.n5951 VCC.n5634 0.0103214
R51865 VCC.n5983 VCC.n5982 0.0103214
R51866 VCC.n5746 VCC.n5745 0.0103214
R51867 VCC.n5781 VCC.n5716 0.0103214
R51868 VCC.n5707 VCC.n5704 0.0103214
R51869 VCC.n5824 VCC.n5823 0.0103214
R51870 VCC.n5850 VCC.n5849 0.0103214
R51871 VCC.n5744 VCC.n5743 0.0103214
R51872 VCC.n5780 VCC.n5717 0.0103214
R51873 VCC.n5825 VCC.n5695 0.0103214
R51874 VCC.n5848 VCC.n5679 0.0103214
R51875 VCC.n5682 VCC.n5676 0.0103214
R51876 VCC.n6297 VCC.n6296 0.0103214
R51877 VCC.n6332 VCC.n6267 0.0103214
R51878 VCC.n6258 VCC.n6255 0.0103214
R51879 VCC.n6375 VCC.n6374 0.0103214
R51880 VCC.n6401 VCC.n6400 0.0103214
R51881 VCC.n6295 VCC.n6294 0.0103214
R51882 VCC.n6331 VCC.n6268 0.0103214
R51883 VCC.n6376 VCC.n6246 0.0103214
R51884 VCC.n6399 VCC.n6230 0.0103214
R51885 VCC.n6233 VCC.n6227 0.0103214
R51886 VCC.n6429 VCC.n6428 0.0103214
R51887 VCC.n6420 VCC.n6213 0.0103214
R51888 VCC.n6448 VCC.n6447 0.0103214
R51889 VCC.n6487 VCC.n6486 0.0103214
R51890 VCC.n6502 VCC.n6501 0.0103214
R51891 VCC.n6535 VCC.n6171 0.0103214
R51892 VCC.n6427 VCC.n6416 0.0103214
R51893 VCC.n6419 VCC.n6212 0.0103214
R51894 VCC.n6446 VCC.n6200 0.0103214
R51895 VCC.n6503 VCC.n6186 0.0103214
R51896 VCC.n6534 VCC.n6533 0.0103214
R51897 VCC.n6564 VCC.n6155 0.0103214
R51898 VCC.n6560 VCC.n6559 0.0103214
R51899 VCC.n6585 VCC.n6142 0.0103214
R51900 VCC.n6607 VCC.n6123 0.0103214
R51901 VCC.n6642 VCC.n6641 0.0103214
R51902 VCC.n6563 VCC.n6157 0.0103214
R51903 VCC.n6584 VCC.n6583 0.0103214
R51904 VCC.n6579 VCC.n6133 0.0103214
R51905 VCC.n6608 VCC.n6125 0.0103214
R51906 VCC.n6616 VCC.n6615 0.0103214
R51907 VCC.n7121 VCC.n6711 0.0103214
R51908 VCC.n6714 VCC.n6713 0.0103214
R51909 VCC.n7134 VCC.n6697 0.0103214
R51910 VCC.n7171 VCC.n7170 0.0103214
R51911 VCC.n7187 VCC.n6670 0.0103214
R51912 VCC.n7109 VCC.n6712 0.0103214
R51913 VCC.n7135 VCC.n6698 0.0103214
R51914 VCC.n7151 VCC.n6696 0.0103214
R51915 VCC.n7172 VCC.n6677 0.0103214
R51916 VCC.n6682 VCC.n6674 0.0103214
R51917 VCC.n6986 VCC.n6780 0.0103214
R51918 VCC.n6977 VCC.n6770 0.0103214
R51919 VCC.n7005 VCC.n7004 0.0103214
R51920 VCC.n7044 VCC.n7043 0.0103214
R51921 VCC.n7059 VCC.n7058 0.0103214
R51922 VCC.n7093 VCC.n6728 0.0103214
R51923 VCC.n6985 VCC.n6984 0.0103214
R51924 VCC.n6976 VCC.n6769 0.0103214
R51925 VCC.n7003 VCC.n6757 0.0103214
R51926 VCC.n7060 VCC.n6743 0.0103214
R51927 VCC.n7092 VCC.n7091 0.0103214
R51928 VCC.n6855 VCC.n6854 0.0103214
R51929 VCC.n6890 VCC.n6825 0.0103214
R51930 VCC.n6816 VCC.n6813 0.0103214
R51931 VCC.n6933 VCC.n6932 0.0103214
R51932 VCC.n6959 VCC.n6958 0.0103214
R51933 VCC.n6853 VCC.n6852 0.0103214
R51934 VCC.n6889 VCC.n6826 0.0103214
R51935 VCC.n6934 VCC.n6804 0.0103214
R51936 VCC.n6957 VCC.n6788 0.0103214
R51937 VCC.n6791 VCC.n6785 0.0103214
R51938 VCC.n7406 VCC.n7405 0.0103214
R51939 VCC.n7441 VCC.n7376 0.0103214
R51940 VCC.n7367 VCC.n7364 0.0103214
R51941 VCC.n7484 VCC.n7483 0.0103214
R51942 VCC.n7510 VCC.n7509 0.0103214
R51943 VCC.n7404 VCC.n7403 0.0103214
R51944 VCC.n7440 VCC.n7377 0.0103214
R51945 VCC.n7485 VCC.n7355 0.0103214
R51946 VCC.n7508 VCC.n7339 0.0103214
R51947 VCC.n7342 VCC.n7336 0.0103214
R51948 VCC.n7538 VCC.n7537 0.0103214
R51949 VCC.n7529 VCC.n7322 0.0103214
R51950 VCC.n7557 VCC.n7556 0.0103214
R51951 VCC.n7596 VCC.n7595 0.0103214
R51952 VCC.n7611 VCC.n7610 0.0103214
R51953 VCC.n7644 VCC.n7280 0.0103214
R51954 VCC.n7536 VCC.n7525 0.0103214
R51955 VCC.n7528 VCC.n7321 0.0103214
R51956 VCC.n7555 VCC.n7309 0.0103214
R51957 VCC.n7612 VCC.n7295 0.0103214
R51958 VCC.n7643 VCC.n7642 0.0103214
R51959 VCC.n7673 VCC.n7264 0.0103214
R51960 VCC.n7669 VCC.n7668 0.0103214
R51961 VCC.n7694 VCC.n7251 0.0103214
R51962 VCC.n7716 VCC.n7232 0.0103214
R51963 VCC.n7751 VCC.n7750 0.0103214
R51964 VCC.n7672 VCC.n7266 0.0103214
R51965 VCC.n7693 VCC.n7692 0.0103214
R51966 VCC.n7688 VCC.n7242 0.0103214
R51967 VCC.n7717 VCC.n7234 0.0103214
R51968 VCC.n7725 VCC.n7724 0.0103214
R51969 VCC.n8230 VCC.n7820 0.0103214
R51970 VCC.n7823 VCC.n7822 0.0103214
R51971 VCC.n8243 VCC.n7806 0.0103214
R51972 VCC.n8280 VCC.n8279 0.0103214
R51973 VCC.n8296 VCC.n7779 0.0103214
R51974 VCC.n8218 VCC.n7821 0.0103214
R51975 VCC.n8244 VCC.n7807 0.0103214
R51976 VCC.n8260 VCC.n7805 0.0103214
R51977 VCC.n8281 VCC.n7786 0.0103214
R51978 VCC.n7791 VCC.n7783 0.0103214
R51979 VCC.n8095 VCC.n7889 0.0103214
R51980 VCC.n8086 VCC.n7879 0.0103214
R51981 VCC.n8114 VCC.n8113 0.0103214
R51982 VCC.n8153 VCC.n8152 0.0103214
R51983 VCC.n8168 VCC.n8167 0.0103214
R51984 VCC.n8202 VCC.n7837 0.0103214
R51985 VCC.n8094 VCC.n8093 0.0103214
R51986 VCC.n8085 VCC.n7878 0.0103214
R51987 VCC.n8112 VCC.n7866 0.0103214
R51988 VCC.n8169 VCC.n7852 0.0103214
R51989 VCC.n8201 VCC.n8200 0.0103214
R51990 VCC.n7964 VCC.n7963 0.0103214
R51991 VCC.n7999 VCC.n7934 0.0103214
R51992 VCC.n7925 VCC.n7922 0.0103214
R51993 VCC.n8042 VCC.n8041 0.0103214
R51994 VCC.n8068 VCC.n8067 0.0103214
R51995 VCC.n7962 VCC.n7961 0.0103214
R51996 VCC.n7998 VCC.n7935 0.0103214
R51997 VCC.n8043 VCC.n7913 0.0103214
R51998 VCC.n8066 VCC.n7897 0.0103214
R51999 VCC.n7900 VCC.n7894 0.0103214
R52000 VCC.n8647 VCC.n8646 0.0103214
R52001 VCC.n8638 VCC.n8431 0.0103214
R52002 VCC.n8666 VCC.n8665 0.0103214
R52003 VCC.n8705 VCC.n8704 0.0103214
R52004 VCC.n8720 VCC.n8719 0.0103214
R52005 VCC.n8753 VCC.n8389 0.0103214
R52006 VCC.n8645 VCC.n8634 0.0103214
R52007 VCC.n8637 VCC.n8430 0.0103214
R52008 VCC.n8664 VCC.n8418 0.0103214
R52009 VCC.n8721 VCC.n8404 0.0103214
R52010 VCC.n8752 VCC.n8751 0.0103214
R52011 VCC.n8782 VCC.n8373 0.0103214
R52012 VCC.n8778 VCC.n8777 0.0103214
R52013 VCC.n8803 VCC.n8360 0.0103214
R52014 VCC.n8825 VCC.n8341 0.0103214
R52015 VCC.n8860 VCC.n8859 0.0103214
R52016 VCC.n8781 VCC.n8375 0.0103214
R52017 VCC.n8802 VCC.n8801 0.0103214
R52018 VCC.n8797 VCC.n8351 0.0103214
R52019 VCC.n8826 VCC.n8343 0.0103214
R52020 VCC.n8834 VCC.n8833 0.0103214
R52021 VCC.n8515 VCC.n8514 0.0103214
R52022 VCC.n8550 VCC.n8485 0.0103214
R52023 VCC.n8476 VCC.n8473 0.0103214
R52024 VCC.n8593 VCC.n8592 0.0103214
R52025 VCC.n8619 VCC.n8618 0.0103214
R52026 VCC.n8513 VCC.n8512 0.0103214
R52027 VCC.n8549 VCC.n8486 0.0103214
R52028 VCC.n8594 VCC.n8464 0.0103214
R52029 VCC.n8617 VCC.n8448 0.0103214
R52030 VCC.n8451 VCC.n8445 0.0103214
R52031 VCC.n9339 VCC.n8929 0.0103214
R52032 VCC.n8932 VCC.n8931 0.0103214
R52033 VCC.n9352 VCC.n8915 0.0103214
R52034 VCC.n9389 VCC.n9388 0.0103214
R52035 VCC.n9405 VCC.n8888 0.0103214
R52036 VCC.n9327 VCC.n8930 0.0103214
R52037 VCC.n9353 VCC.n8916 0.0103214
R52038 VCC.n9369 VCC.n8914 0.0103214
R52039 VCC.n9390 VCC.n8895 0.0103214
R52040 VCC.n8900 VCC.n8892 0.0103214
R52041 VCC.n9204 VCC.n8998 0.0103214
R52042 VCC.n9195 VCC.n8988 0.0103214
R52043 VCC.n9223 VCC.n9222 0.0103214
R52044 VCC.n9262 VCC.n9261 0.0103214
R52045 VCC.n9277 VCC.n9276 0.0103214
R52046 VCC.n9311 VCC.n8946 0.0103214
R52047 VCC.n9203 VCC.n9202 0.0103214
R52048 VCC.n9194 VCC.n8987 0.0103214
R52049 VCC.n9221 VCC.n8975 0.0103214
R52050 VCC.n9278 VCC.n8961 0.0103214
R52051 VCC.n9310 VCC.n9309 0.0103214
R52052 VCC.n9073 VCC.n9072 0.0103214
R52053 VCC.n9108 VCC.n9043 0.0103214
R52054 VCC.n9034 VCC.n9031 0.0103214
R52055 VCC.n9151 VCC.n9150 0.0103214
R52056 VCC.n9177 VCC.n9176 0.0103214
R52057 VCC.n9071 VCC.n9070 0.0103214
R52058 VCC.n9107 VCC.n9044 0.0103214
R52059 VCC.n9152 VCC.n9022 0.0103214
R52060 VCC.n9175 VCC.n9006 0.0103214
R52061 VCC.n9009 VCC.n9003 0.0103214
R52062 VCC.n9624 VCC.n9623 0.0103214
R52063 VCC.n9659 VCC.n9594 0.0103214
R52064 VCC.n9585 VCC.n9582 0.0103214
R52065 VCC.n9702 VCC.n9701 0.0103214
R52066 VCC.n9728 VCC.n9727 0.0103214
R52067 VCC.n9622 VCC.n9621 0.0103214
R52068 VCC.n9658 VCC.n9595 0.0103214
R52069 VCC.n9703 VCC.n9573 0.0103214
R52070 VCC.n9726 VCC.n9557 0.0103214
R52071 VCC.n9560 VCC.n9554 0.0103214
R52072 VCC.n9756 VCC.n9755 0.0103214
R52073 VCC.n9747 VCC.n9540 0.0103214
R52074 VCC.n9775 VCC.n9774 0.0103214
R52075 VCC.n9814 VCC.n9813 0.0103214
R52076 VCC.n9829 VCC.n9828 0.0103214
R52077 VCC.n9862 VCC.n9498 0.0103214
R52078 VCC.n9754 VCC.n9743 0.0103214
R52079 VCC.n9746 VCC.n9539 0.0103214
R52080 VCC.n9773 VCC.n9527 0.0103214
R52081 VCC.n9830 VCC.n9513 0.0103214
R52082 VCC.n9861 VCC.n9860 0.0103214
R52083 VCC.n9891 VCC.n9482 0.0103214
R52084 VCC.n9887 VCC.n9886 0.0103214
R52085 VCC.n9912 VCC.n9469 0.0103214
R52086 VCC.n9934 VCC.n9450 0.0103214
R52087 VCC.n9969 VCC.n9968 0.0103214
R52088 VCC.n9890 VCC.n9484 0.0103214
R52089 VCC.n9911 VCC.n9910 0.0103214
R52090 VCC.n9906 VCC.n9460 0.0103214
R52091 VCC.n9935 VCC.n9452 0.0103214
R52092 VCC.n9943 VCC.n9942 0.0103214
R52093 VCC.n10447 VCC.n10037 0.0103214
R52094 VCC.n10040 VCC.n10039 0.0103214
R52095 VCC.n10460 VCC.n10023 0.0103214
R52096 VCC.n10497 VCC.n10496 0.0103214
R52097 VCC.n10513 VCC.n9996 0.0103214
R52098 VCC.n10435 VCC.n10038 0.0103214
R52099 VCC.n10461 VCC.n10024 0.0103214
R52100 VCC.n10477 VCC.n10022 0.0103214
R52101 VCC.n10498 VCC.n10003 0.0103214
R52102 VCC.n10008 VCC.n10000 0.0103214
R52103 VCC.n10312 VCC.n10106 0.0103214
R52104 VCC.n10303 VCC.n10096 0.0103214
R52105 VCC.n10331 VCC.n10330 0.0103214
R52106 VCC.n10370 VCC.n10369 0.0103214
R52107 VCC.n10385 VCC.n10384 0.0103214
R52108 VCC.n10419 VCC.n10054 0.0103214
R52109 VCC.n10311 VCC.n10310 0.0103214
R52110 VCC.n10302 VCC.n10095 0.0103214
R52111 VCC.n10329 VCC.n10083 0.0103214
R52112 VCC.n10386 VCC.n10069 0.0103214
R52113 VCC.n10418 VCC.n10417 0.0103214
R52114 VCC.n10181 VCC.n10180 0.0103214
R52115 VCC.n10216 VCC.n10151 0.0103214
R52116 VCC.n10142 VCC.n10139 0.0103214
R52117 VCC.n10259 VCC.n10258 0.0103214
R52118 VCC.n10285 VCC.n10284 0.0103214
R52119 VCC.n10179 VCC.n10178 0.0103214
R52120 VCC.n10215 VCC.n10152 0.0103214
R52121 VCC.n10260 VCC.n10130 0.0103214
R52122 VCC.n10283 VCC.n10114 0.0103214
R52123 VCC.n10117 VCC.n10111 0.0103214
R52124 VCC.n10731 VCC.n10730 0.0103214
R52125 VCC.n10766 VCC.n10701 0.0103214
R52126 VCC.n10692 VCC.n10689 0.0103214
R52127 VCC.n10809 VCC.n10808 0.0103214
R52128 VCC.n10835 VCC.n10834 0.0103214
R52129 VCC.n10729 VCC.n10728 0.0103214
R52130 VCC.n10765 VCC.n10702 0.0103214
R52131 VCC.n10810 VCC.n10680 0.0103214
R52132 VCC.n10833 VCC.n10664 0.0103214
R52133 VCC.n10667 VCC.n10661 0.0103214
R52134 VCC.n10863 VCC.n10862 0.0103214
R52135 VCC.n10854 VCC.n10647 0.0103214
R52136 VCC.n10882 VCC.n10881 0.0103214
R52137 VCC.n10921 VCC.n10920 0.0103214
R52138 VCC.n10936 VCC.n10935 0.0103214
R52139 VCC.n10969 VCC.n10605 0.0103214
R52140 VCC.n10861 VCC.n10850 0.0103214
R52141 VCC.n10853 VCC.n10646 0.0103214
R52142 VCC.n10880 VCC.n10634 0.0103214
R52143 VCC.n10937 VCC.n10620 0.0103214
R52144 VCC.n10968 VCC.n10967 0.0103214
R52145 VCC.n10998 VCC.n10589 0.0103214
R52146 VCC.n10994 VCC.n10993 0.0103214
R52147 VCC.n11019 VCC.n10576 0.0103214
R52148 VCC.n11041 VCC.n10557 0.0103214
R52149 VCC.n11076 VCC.n11075 0.0103214
R52150 VCC.n10997 VCC.n10591 0.0103214
R52151 VCC.n11018 VCC.n11017 0.0103214
R52152 VCC.n11013 VCC.n10567 0.0103214
R52153 VCC.n11042 VCC.n10559 0.0103214
R52154 VCC.n11050 VCC.n11049 0.0103214
R52155 VCC.n11554 VCC.n11144 0.0103214
R52156 VCC.n11147 VCC.n11146 0.0103214
R52157 VCC.n11567 VCC.n11130 0.0103214
R52158 VCC.n11604 VCC.n11603 0.0103214
R52159 VCC.n11620 VCC.n11103 0.0103214
R52160 VCC.n11542 VCC.n11145 0.0103214
R52161 VCC.n11568 VCC.n11131 0.0103214
R52162 VCC.n11584 VCC.n11129 0.0103214
R52163 VCC.n11605 VCC.n11110 0.0103214
R52164 VCC.n11115 VCC.n11107 0.0103214
R52165 VCC.n11419 VCC.n11213 0.0103214
R52166 VCC.n11410 VCC.n11203 0.0103214
R52167 VCC.n11438 VCC.n11437 0.0103214
R52168 VCC.n11477 VCC.n11476 0.0103214
R52169 VCC.n11492 VCC.n11491 0.0103214
R52170 VCC.n11526 VCC.n11161 0.0103214
R52171 VCC.n11418 VCC.n11417 0.0103214
R52172 VCC.n11409 VCC.n11202 0.0103214
R52173 VCC.n11436 VCC.n11190 0.0103214
R52174 VCC.n11493 VCC.n11176 0.0103214
R52175 VCC.n11525 VCC.n11524 0.0103214
R52176 VCC.n11288 VCC.n11287 0.0103214
R52177 VCC.n11323 VCC.n11258 0.0103214
R52178 VCC.n11249 VCC.n11246 0.0103214
R52179 VCC.n11366 VCC.n11365 0.0103214
R52180 VCC.n11392 VCC.n11391 0.0103214
R52181 VCC.n11286 VCC.n11285 0.0103214
R52182 VCC.n11322 VCC.n11259 0.0103214
R52183 VCC.n11367 VCC.n11237 0.0103214
R52184 VCC.n11390 VCC.n11221 0.0103214
R52185 VCC.n11224 VCC.n11218 0.0103214
R52186 VCC.n11838 VCC.n11837 0.0103214
R52187 VCC.n11873 VCC.n11808 0.0103214
R52188 VCC.n11799 VCC.n11796 0.0103214
R52189 VCC.n11916 VCC.n11915 0.0103214
R52190 VCC.n11942 VCC.n11941 0.0103214
R52191 VCC.n11836 VCC.n11835 0.0103214
R52192 VCC.n11872 VCC.n11809 0.0103214
R52193 VCC.n11917 VCC.n11787 0.0103214
R52194 VCC.n11940 VCC.n11771 0.0103214
R52195 VCC.n11774 VCC.n11768 0.0103214
R52196 VCC.n11970 VCC.n11969 0.0103214
R52197 VCC.n11961 VCC.n11754 0.0103214
R52198 VCC.n11989 VCC.n11988 0.0103214
R52199 VCC.n12028 VCC.n12027 0.0103214
R52200 VCC.n12043 VCC.n12042 0.0103214
R52201 VCC.n12076 VCC.n11712 0.0103214
R52202 VCC.n11968 VCC.n11957 0.0103214
R52203 VCC.n11960 VCC.n11753 0.0103214
R52204 VCC.n11987 VCC.n11741 0.0103214
R52205 VCC.n12044 VCC.n11727 0.0103214
R52206 VCC.n12075 VCC.n12074 0.0103214
R52207 VCC.n12105 VCC.n11696 0.0103214
R52208 VCC.n12101 VCC.n12100 0.0103214
R52209 VCC.n12126 VCC.n11683 0.0103214
R52210 VCC.n12148 VCC.n11664 0.0103214
R52211 VCC.n12183 VCC.n12182 0.0103214
R52212 VCC.n12104 VCC.n11698 0.0103214
R52213 VCC.n12125 VCC.n12124 0.0103214
R52214 VCC.n12120 VCC.n11674 0.0103214
R52215 VCC.n12149 VCC.n11666 0.0103214
R52216 VCC.n12157 VCC.n12156 0.0103214
R52217 VCC.n12661 VCC.n12251 0.0103214
R52218 VCC.n12254 VCC.n12253 0.0103214
R52219 VCC.n12674 VCC.n12237 0.0103214
R52220 VCC.n12711 VCC.n12710 0.0103214
R52221 VCC.n12727 VCC.n12210 0.0103214
R52222 VCC.n12649 VCC.n12252 0.0103214
R52223 VCC.n12675 VCC.n12238 0.0103214
R52224 VCC.n12691 VCC.n12236 0.0103214
R52225 VCC.n12712 VCC.n12217 0.0103214
R52226 VCC.n12222 VCC.n12214 0.0103214
R52227 VCC.n12526 VCC.n12320 0.0103214
R52228 VCC.n12517 VCC.n12310 0.0103214
R52229 VCC.n12545 VCC.n12544 0.0103214
R52230 VCC.n12584 VCC.n12583 0.0103214
R52231 VCC.n12599 VCC.n12598 0.0103214
R52232 VCC.n12633 VCC.n12268 0.0103214
R52233 VCC.n12525 VCC.n12524 0.0103214
R52234 VCC.n12516 VCC.n12309 0.0103214
R52235 VCC.n12543 VCC.n12297 0.0103214
R52236 VCC.n12600 VCC.n12283 0.0103214
R52237 VCC.n12632 VCC.n12631 0.0103214
R52238 VCC.n12395 VCC.n12394 0.0103214
R52239 VCC.n12430 VCC.n12365 0.0103214
R52240 VCC.n12356 VCC.n12353 0.0103214
R52241 VCC.n12473 VCC.n12472 0.0103214
R52242 VCC.n12499 VCC.n12498 0.0103214
R52243 VCC.n12393 VCC.n12392 0.0103214
R52244 VCC.n12429 VCC.n12366 0.0103214
R52245 VCC.n12474 VCC.n12344 0.0103214
R52246 VCC.n12497 VCC.n12328 0.0103214
R52247 VCC.n12331 VCC.n12325 0.0103214
R52248 VCC.n12945 VCC.n12944 0.0103214
R52249 VCC.n12980 VCC.n12915 0.0103214
R52250 VCC.n12906 VCC.n12903 0.0103214
R52251 VCC.n13023 VCC.n13022 0.0103214
R52252 VCC.n13049 VCC.n13048 0.0103214
R52253 VCC.n12943 VCC.n12942 0.0103214
R52254 VCC.n12979 VCC.n12916 0.0103214
R52255 VCC.n13024 VCC.n12894 0.0103214
R52256 VCC.n13047 VCC.n12878 0.0103214
R52257 VCC.n12881 VCC.n12875 0.0103214
R52258 VCC.n13077 VCC.n13076 0.0103214
R52259 VCC.n13068 VCC.n12861 0.0103214
R52260 VCC.n13096 VCC.n13095 0.0103214
R52261 VCC.n13135 VCC.n13134 0.0103214
R52262 VCC.n13150 VCC.n13149 0.0103214
R52263 VCC.n13183 VCC.n12819 0.0103214
R52264 VCC.n13075 VCC.n13064 0.0103214
R52265 VCC.n13067 VCC.n12860 0.0103214
R52266 VCC.n13094 VCC.n12848 0.0103214
R52267 VCC.n13151 VCC.n12834 0.0103214
R52268 VCC.n13182 VCC.n13181 0.0103214
R52269 VCC.n13212 VCC.n12803 0.0103214
R52270 VCC.n13208 VCC.n13207 0.0103214
R52271 VCC.n13233 VCC.n12790 0.0103214
R52272 VCC.n13255 VCC.n12771 0.0103214
R52273 VCC.n13290 VCC.n13289 0.0103214
R52274 VCC.n13211 VCC.n12805 0.0103214
R52275 VCC.n13232 VCC.n13231 0.0103214
R52276 VCC.n13227 VCC.n12781 0.0103214
R52277 VCC.n13256 VCC.n12773 0.0103214
R52278 VCC.n13264 VCC.n13263 0.0103214
R52279 VCC.n13768 VCC.n13358 0.0103214
R52280 VCC.n13361 VCC.n13360 0.0103214
R52281 VCC.n13781 VCC.n13344 0.0103214
R52282 VCC.n13818 VCC.n13817 0.0103214
R52283 VCC.n13834 VCC.n13317 0.0103214
R52284 VCC.n13756 VCC.n13359 0.0103214
R52285 VCC.n13782 VCC.n13345 0.0103214
R52286 VCC.n13798 VCC.n13343 0.0103214
R52287 VCC.n13819 VCC.n13324 0.0103214
R52288 VCC.n13329 VCC.n13321 0.0103214
R52289 VCC.n13633 VCC.n13427 0.0103214
R52290 VCC.n13624 VCC.n13417 0.0103214
R52291 VCC.n13652 VCC.n13651 0.0103214
R52292 VCC.n13691 VCC.n13690 0.0103214
R52293 VCC.n13706 VCC.n13705 0.0103214
R52294 VCC.n13740 VCC.n13375 0.0103214
R52295 VCC.n13632 VCC.n13631 0.0103214
R52296 VCC.n13623 VCC.n13416 0.0103214
R52297 VCC.n13650 VCC.n13404 0.0103214
R52298 VCC.n13707 VCC.n13390 0.0103214
R52299 VCC.n13739 VCC.n13738 0.0103214
R52300 VCC.n13502 VCC.n13501 0.0103214
R52301 VCC.n13537 VCC.n13472 0.0103214
R52302 VCC.n13463 VCC.n13460 0.0103214
R52303 VCC.n13580 VCC.n13579 0.0103214
R52304 VCC.n13606 VCC.n13605 0.0103214
R52305 VCC.n13500 VCC.n13499 0.0103214
R52306 VCC.n13536 VCC.n13473 0.0103214
R52307 VCC.n13581 VCC.n13451 0.0103214
R52308 VCC.n13604 VCC.n13435 0.0103214
R52309 VCC.n13438 VCC.n13432 0.0103214
R52310 VCC.n14052 VCC.n14051 0.0103214
R52311 VCC.n14087 VCC.n14022 0.0103214
R52312 VCC.n14013 VCC.n14010 0.0103214
R52313 VCC.n14130 VCC.n14129 0.0103214
R52314 VCC.n14156 VCC.n14155 0.0103214
R52315 VCC.n14050 VCC.n14049 0.0103214
R52316 VCC.n14086 VCC.n14023 0.0103214
R52317 VCC.n14131 VCC.n14001 0.0103214
R52318 VCC.n14154 VCC.n13985 0.0103214
R52319 VCC.n13988 VCC.n13982 0.0103214
R52320 VCC.n14184 VCC.n14183 0.0103214
R52321 VCC.n14175 VCC.n13968 0.0103214
R52322 VCC.n14203 VCC.n14202 0.0103214
R52323 VCC.n14242 VCC.n14241 0.0103214
R52324 VCC.n14257 VCC.n14256 0.0103214
R52325 VCC.n14290 VCC.n13926 0.0103214
R52326 VCC.n14182 VCC.n14171 0.0103214
R52327 VCC.n14174 VCC.n13967 0.0103214
R52328 VCC.n14201 VCC.n13955 0.0103214
R52329 VCC.n14258 VCC.n13941 0.0103214
R52330 VCC.n14289 VCC.n14288 0.0103214
R52331 VCC.n14319 VCC.n13910 0.0103214
R52332 VCC.n14315 VCC.n14314 0.0103214
R52333 VCC.n14340 VCC.n13897 0.0103214
R52334 VCC.n14362 VCC.n13878 0.0103214
R52335 VCC.n14397 VCC.n14396 0.0103214
R52336 VCC.n14318 VCC.n13912 0.0103214
R52337 VCC.n14339 VCC.n14338 0.0103214
R52338 VCC.n14334 VCC.n13888 0.0103214
R52339 VCC.n14363 VCC.n13880 0.0103214
R52340 VCC.n14371 VCC.n14370 0.0103214
R52341 VCC.n14875 VCC.n14465 0.0103214
R52342 VCC.n14468 VCC.n14467 0.0103214
R52343 VCC.n14888 VCC.n14451 0.0103214
R52344 VCC.n14925 VCC.n14924 0.0103214
R52345 VCC.n14941 VCC.n14424 0.0103214
R52346 VCC.n14863 VCC.n14466 0.0103214
R52347 VCC.n14889 VCC.n14452 0.0103214
R52348 VCC.n14905 VCC.n14450 0.0103214
R52349 VCC.n14926 VCC.n14431 0.0103214
R52350 VCC.n14436 VCC.n14428 0.0103214
R52351 VCC.n14740 VCC.n14534 0.0103214
R52352 VCC.n14731 VCC.n14524 0.0103214
R52353 VCC.n14759 VCC.n14758 0.0103214
R52354 VCC.n14798 VCC.n14797 0.0103214
R52355 VCC.n14813 VCC.n14812 0.0103214
R52356 VCC.n14847 VCC.n14482 0.0103214
R52357 VCC.n14739 VCC.n14738 0.0103214
R52358 VCC.n14730 VCC.n14523 0.0103214
R52359 VCC.n14757 VCC.n14511 0.0103214
R52360 VCC.n14814 VCC.n14497 0.0103214
R52361 VCC.n14846 VCC.n14845 0.0103214
R52362 VCC.n14609 VCC.n14608 0.0103214
R52363 VCC.n14644 VCC.n14579 0.0103214
R52364 VCC.n14570 VCC.n14567 0.0103214
R52365 VCC.n14687 VCC.n14686 0.0103214
R52366 VCC.n14713 VCC.n14712 0.0103214
R52367 VCC.n14607 VCC.n14606 0.0103214
R52368 VCC.n14643 VCC.n14580 0.0103214
R52369 VCC.n14688 VCC.n14558 0.0103214
R52370 VCC.n14711 VCC.n14542 0.0103214
R52371 VCC.n14545 VCC.n14539 0.0103214
R52372 VCC.n15159 VCC.n15158 0.0103214
R52373 VCC.n15194 VCC.n15129 0.0103214
R52374 VCC.n15120 VCC.n15117 0.0103214
R52375 VCC.n15237 VCC.n15236 0.0103214
R52376 VCC.n15263 VCC.n15262 0.0103214
R52377 VCC.n15157 VCC.n15156 0.0103214
R52378 VCC.n15193 VCC.n15130 0.0103214
R52379 VCC.n15238 VCC.n15108 0.0103214
R52380 VCC.n15261 VCC.n15092 0.0103214
R52381 VCC.n15095 VCC.n15089 0.0103214
R52382 VCC.n15291 VCC.n15290 0.0103214
R52383 VCC.n15282 VCC.n15075 0.0103214
R52384 VCC.n15310 VCC.n15309 0.0103214
R52385 VCC.n15349 VCC.n15348 0.0103214
R52386 VCC.n15364 VCC.n15363 0.0103214
R52387 VCC.n15397 VCC.n15033 0.0103214
R52388 VCC.n15289 VCC.n15278 0.0103214
R52389 VCC.n15281 VCC.n15074 0.0103214
R52390 VCC.n15308 VCC.n15062 0.0103214
R52391 VCC.n15365 VCC.n15048 0.0103214
R52392 VCC.n15396 VCC.n15395 0.0103214
R52393 VCC.n15426 VCC.n15017 0.0103214
R52394 VCC.n15422 VCC.n15421 0.0103214
R52395 VCC.n15447 VCC.n15004 0.0103214
R52396 VCC.n15469 VCC.n14985 0.0103214
R52397 VCC.n15504 VCC.n15503 0.0103214
R52398 VCC.n15425 VCC.n15019 0.0103214
R52399 VCC.n15446 VCC.n15445 0.0103214
R52400 VCC.n15441 VCC.n14995 0.0103214
R52401 VCC.n15470 VCC.n14987 0.0103214
R52402 VCC.n15478 VCC.n15477 0.0103214
R52403 VCC.n15982 VCC.n15572 0.0103214
R52404 VCC.n15575 VCC.n15574 0.0103214
R52405 VCC.n15995 VCC.n15558 0.0103214
R52406 VCC.n16032 VCC.n16031 0.0103214
R52407 VCC.n16048 VCC.n15531 0.0103214
R52408 VCC.n15970 VCC.n15573 0.0103214
R52409 VCC.n15996 VCC.n15559 0.0103214
R52410 VCC.n16012 VCC.n15557 0.0103214
R52411 VCC.n16033 VCC.n15538 0.0103214
R52412 VCC.n15543 VCC.n15535 0.0103214
R52413 VCC.n15847 VCC.n15641 0.0103214
R52414 VCC.n15838 VCC.n15631 0.0103214
R52415 VCC.n15866 VCC.n15865 0.0103214
R52416 VCC.n15905 VCC.n15904 0.0103214
R52417 VCC.n15920 VCC.n15919 0.0103214
R52418 VCC.n15954 VCC.n15589 0.0103214
R52419 VCC.n15846 VCC.n15845 0.0103214
R52420 VCC.n15837 VCC.n15630 0.0103214
R52421 VCC.n15864 VCC.n15618 0.0103214
R52422 VCC.n15921 VCC.n15604 0.0103214
R52423 VCC.n15953 VCC.n15952 0.0103214
R52424 VCC.n15716 VCC.n15715 0.0103214
R52425 VCC.n15751 VCC.n15686 0.0103214
R52426 VCC.n15677 VCC.n15674 0.0103214
R52427 VCC.n15794 VCC.n15793 0.0103214
R52428 VCC.n15820 VCC.n15819 0.0103214
R52429 VCC.n15714 VCC.n15713 0.0103214
R52430 VCC.n15750 VCC.n15687 0.0103214
R52431 VCC.n15795 VCC.n15665 0.0103214
R52432 VCC.n15818 VCC.n15649 0.0103214
R52433 VCC.n15652 VCC.n15646 0.0103214
R52434 VCC.n16266 VCC.n16265 0.0103214
R52435 VCC.n16301 VCC.n16236 0.0103214
R52436 VCC.n16227 VCC.n16224 0.0103214
R52437 VCC.n16344 VCC.n16343 0.0103214
R52438 VCC.n16370 VCC.n16369 0.0103214
R52439 VCC.n16264 VCC.n16263 0.0103214
R52440 VCC.n16300 VCC.n16237 0.0103214
R52441 VCC.n16345 VCC.n16215 0.0103214
R52442 VCC.n16368 VCC.n16199 0.0103214
R52443 VCC.n16202 VCC.n16196 0.0103214
R52444 VCC.n16398 VCC.n16397 0.0103214
R52445 VCC.n16389 VCC.n16182 0.0103214
R52446 VCC.n16417 VCC.n16416 0.0103214
R52447 VCC.n16456 VCC.n16455 0.0103214
R52448 VCC.n16471 VCC.n16470 0.0103214
R52449 VCC.n16504 VCC.n16140 0.0103214
R52450 VCC.n16396 VCC.n16385 0.0103214
R52451 VCC.n16388 VCC.n16181 0.0103214
R52452 VCC.n16415 VCC.n16169 0.0103214
R52453 VCC.n16472 VCC.n16155 0.0103214
R52454 VCC.n16503 VCC.n16502 0.0103214
R52455 VCC.n16533 VCC.n16124 0.0103214
R52456 VCC.n16529 VCC.n16528 0.0103214
R52457 VCC.n16554 VCC.n16111 0.0103214
R52458 VCC.n16576 VCC.n16092 0.0103214
R52459 VCC.n16611 VCC.n16610 0.0103214
R52460 VCC.n16532 VCC.n16126 0.0103214
R52461 VCC.n16553 VCC.n16552 0.0103214
R52462 VCC.n16548 VCC.n16102 0.0103214
R52463 VCC.n16577 VCC.n16094 0.0103214
R52464 VCC.n16585 VCC.n16584 0.0103214
R52465 VCC.n17089 VCC.n16679 0.0103214
R52466 VCC.n16682 VCC.n16681 0.0103214
R52467 VCC.n17102 VCC.n16665 0.0103214
R52468 VCC.n17139 VCC.n17138 0.0103214
R52469 VCC.n17155 VCC.n16638 0.0103214
R52470 VCC.n17077 VCC.n16680 0.0103214
R52471 VCC.n17103 VCC.n16666 0.0103214
R52472 VCC.n17119 VCC.n16664 0.0103214
R52473 VCC.n17140 VCC.n16645 0.0103214
R52474 VCC.n16650 VCC.n16642 0.0103214
R52475 VCC.n16954 VCC.n16748 0.0103214
R52476 VCC.n16945 VCC.n16738 0.0103214
R52477 VCC.n16973 VCC.n16972 0.0103214
R52478 VCC.n17012 VCC.n17011 0.0103214
R52479 VCC.n17027 VCC.n17026 0.0103214
R52480 VCC.n17061 VCC.n16696 0.0103214
R52481 VCC.n16953 VCC.n16952 0.0103214
R52482 VCC.n16944 VCC.n16737 0.0103214
R52483 VCC.n16971 VCC.n16725 0.0103214
R52484 VCC.n17028 VCC.n16711 0.0103214
R52485 VCC.n17060 VCC.n17059 0.0103214
R52486 VCC.n16823 VCC.n16822 0.0103214
R52487 VCC.n16858 VCC.n16793 0.0103214
R52488 VCC.n16784 VCC.n16781 0.0103214
R52489 VCC.n16901 VCC.n16900 0.0103214
R52490 VCC.n16927 VCC.n16926 0.0103214
R52491 VCC.n16821 VCC.n16820 0.0103214
R52492 VCC.n16857 VCC.n16794 0.0103214
R52493 VCC.n16902 VCC.n16772 0.0103214
R52494 VCC.n16925 VCC.n16756 0.0103214
R52495 VCC.n16759 VCC.n16753 0.0103214
R52496 VCC.n17318 VCC.n17317 0.0103214
R52497 VCC.n17309 VCC.n17289 0.0103214
R52498 VCC.n17337 VCC.n17336 0.0103214
R52499 VCC.n17376 VCC.n17375 0.0103214
R52500 VCC.n17391 VCC.n17390 0.0103214
R52501 VCC.n17424 VCC.n17247 0.0103214
R52502 VCC.n17316 VCC.n17305 0.0103214
R52503 VCC.n17308 VCC.n17288 0.0103214
R52504 VCC.n17335 VCC.n17276 0.0103214
R52505 VCC.n17392 VCC.n17262 0.0103214
R52506 VCC.n17423 VCC.n17422 0.0103214
R52507 VCC.n17453 VCC.n17231 0.0103214
R52508 VCC.n17449 VCC.n17448 0.0103214
R52509 VCC.n17474 VCC.n17218 0.0103214
R52510 VCC.n17496 VCC.n17199 0.0103214
R52511 VCC.n17531 VCC.n17530 0.0103214
R52512 VCC.n17452 VCC.n17233 0.0103214
R52513 VCC.n17473 VCC.n17472 0.0103214
R52514 VCC.n17468 VCC.n17209 0.0103214
R52515 VCC.n17497 VCC.n17201 0.0103214
R52516 VCC.n17505 VCC.n17504 0.0103214
R52517 VCC.n206 VCC.n193 0.00942857
R52518 VCC.n246 VCC.n168 0.00942857
R52519 VCC.n262 VCC.n162 0.00942857
R52520 VCC.n294 VCC.n138 0.00942857
R52521 VCC.n205 VCC.n190 0.00942857
R52522 VCC.n261 VCC.n260 0.00942857
R52523 VCC.n367 VCC.n105 0.00942857
R52524 VCC.n383 VCC.n98 0.00942857
R52525 VCC.n77 VCC.n68 0.00942857
R52526 VCC.n382 VCC.n100 0.00942857
R52527 VCC.n75 VCC.n69 0.00942857
R52528 VCC.n457 VCC.n456 0.00942857
R52529 VCC.n534 VCC.n16 0.00942857
R52530 VCC.n19 VCC.n17 0.00942857
R52531 VCC.n455 VCC.n64 0.00942857
R52532 VCC.n479 VCC.n51 0.00942857
R52533 VCC.n507 VCC.n506 0.00942857
R52534 VCC.n18 VCC.n10 0.00942857
R52535 VCC.n758 VCC.n745 0.00942857
R52536 VCC.n798 VCC.n720 0.00942857
R52537 VCC.n814 VCC.n714 0.00942857
R52538 VCC.n846 VCC.n690 0.00942857
R52539 VCC.n757 VCC.n742 0.00942857
R52540 VCC.n813 VCC.n812 0.00942857
R52541 VCC.n919 VCC.n657 0.00942857
R52542 VCC.n935 VCC.n650 0.00942857
R52543 VCC.n629 VCC.n620 0.00942857
R52544 VCC.n934 VCC.n652 0.00942857
R52545 VCC.n627 VCC.n621 0.00942857
R52546 VCC.n1009 VCC.n1008 0.00942857
R52547 VCC.n1086 VCC.n568 0.00942857
R52548 VCC.n571 VCC.n569 0.00942857
R52549 VCC.n1007 VCC.n616 0.00942857
R52550 VCC.n1031 VCC.n603 0.00942857
R52551 VCC.n1059 VCC.n1058 0.00942857
R52552 VCC.n570 VCC.n564 0.00942857
R52553 VCC.n1568 VCC.n1567 0.00942857
R52554 VCC.n1633 VCC.n1632 0.00942857
R52555 VCC.n1646 VCC.n1119 0.00942857
R52556 VCC.n1566 VCC.n1173 0.00942857
R52557 VCC.n1597 VCC.n1156 0.00942857
R52558 VCC.n1610 VCC.n1149 0.00942857
R52559 VCC.n1645 VCC.n1644 0.00942857
R52560 VCC.n1476 VCC.n1214 0.00942857
R52561 VCC.n1492 VCC.n1207 0.00942857
R52562 VCC.n1186 VCC.n1177 0.00942857
R52563 VCC.n1491 VCC.n1209 0.00942857
R52564 VCC.n1184 VCC.n1178 0.00942857
R52565 VCC.n1316 VCC.n1303 0.00942857
R52566 VCC.n1356 VCC.n1278 0.00942857
R52567 VCC.n1372 VCC.n1272 0.00942857
R52568 VCC.n1404 VCC.n1248 0.00942857
R52569 VCC.n1315 VCC.n1300 0.00942857
R52570 VCC.n1371 VCC.n1370 0.00942857
R52571 VCC.n1867 VCC.n1854 0.00942857
R52572 VCC.n1907 VCC.n1829 0.00942857
R52573 VCC.n1923 VCC.n1823 0.00942857
R52574 VCC.n1955 VCC.n1799 0.00942857
R52575 VCC.n1866 VCC.n1851 0.00942857
R52576 VCC.n1922 VCC.n1921 0.00942857
R52577 VCC.n2028 VCC.n1766 0.00942857
R52578 VCC.n2044 VCC.n1759 0.00942857
R52579 VCC.n1738 VCC.n1729 0.00942857
R52580 VCC.n2043 VCC.n1761 0.00942857
R52581 VCC.n1736 VCC.n1730 0.00942857
R52582 VCC.n2118 VCC.n2117 0.00942857
R52583 VCC.n2195 VCC.n1677 0.00942857
R52584 VCC.n1680 VCC.n1678 0.00942857
R52585 VCC.n2116 VCC.n1725 0.00942857
R52586 VCC.n2140 VCC.n1712 0.00942857
R52587 VCC.n2168 VCC.n2167 0.00942857
R52588 VCC.n1679 VCC.n1673 0.00942857
R52589 VCC.n2677 VCC.n2676 0.00942857
R52590 VCC.n2742 VCC.n2741 0.00942857
R52591 VCC.n2755 VCC.n2228 0.00942857
R52592 VCC.n2675 VCC.n2282 0.00942857
R52593 VCC.n2706 VCC.n2265 0.00942857
R52594 VCC.n2719 VCC.n2258 0.00942857
R52595 VCC.n2754 VCC.n2753 0.00942857
R52596 VCC.n2585 VCC.n2323 0.00942857
R52597 VCC.n2601 VCC.n2316 0.00942857
R52598 VCC.n2295 VCC.n2286 0.00942857
R52599 VCC.n2600 VCC.n2318 0.00942857
R52600 VCC.n2293 VCC.n2287 0.00942857
R52601 VCC.n2425 VCC.n2412 0.00942857
R52602 VCC.n2465 VCC.n2387 0.00942857
R52603 VCC.n2481 VCC.n2381 0.00942857
R52604 VCC.n2513 VCC.n2357 0.00942857
R52605 VCC.n2424 VCC.n2409 0.00942857
R52606 VCC.n2480 VCC.n2479 0.00942857
R52607 VCC.n2976 VCC.n2963 0.00942857
R52608 VCC.n3016 VCC.n2938 0.00942857
R52609 VCC.n3032 VCC.n2932 0.00942857
R52610 VCC.n3064 VCC.n2908 0.00942857
R52611 VCC.n2975 VCC.n2960 0.00942857
R52612 VCC.n3031 VCC.n3030 0.00942857
R52613 VCC.n3137 VCC.n2875 0.00942857
R52614 VCC.n3153 VCC.n2868 0.00942857
R52615 VCC.n2847 VCC.n2838 0.00942857
R52616 VCC.n3152 VCC.n2870 0.00942857
R52617 VCC.n2845 VCC.n2839 0.00942857
R52618 VCC.n3227 VCC.n3226 0.00942857
R52619 VCC.n3304 VCC.n2786 0.00942857
R52620 VCC.n2789 VCC.n2787 0.00942857
R52621 VCC.n3225 VCC.n2834 0.00942857
R52622 VCC.n3249 VCC.n2821 0.00942857
R52623 VCC.n3277 VCC.n3276 0.00942857
R52624 VCC.n2788 VCC.n2782 0.00942857
R52625 VCC.n3786 VCC.n3785 0.00942857
R52626 VCC.n3851 VCC.n3850 0.00942857
R52627 VCC.n3864 VCC.n3337 0.00942857
R52628 VCC.n3784 VCC.n3391 0.00942857
R52629 VCC.n3815 VCC.n3374 0.00942857
R52630 VCC.n3828 VCC.n3367 0.00942857
R52631 VCC.n3863 VCC.n3862 0.00942857
R52632 VCC.n3694 VCC.n3432 0.00942857
R52633 VCC.n3710 VCC.n3425 0.00942857
R52634 VCC.n3404 VCC.n3395 0.00942857
R52635 VCC.n3709 VCC.n3427 0.00942857
R52636 VCC.n3402 VCC.n3396 0.00942857
R52637 VCC.n3534 VCC.n3521 0.00942857
R52638 VCC.n3574 VCC.n3496 0.00942857
R52639 VCC.n3590 VCC.n3490 0.00942857
R52640 VCC.n3622 VCC.n3466 0.00942857
R52641 VCC.n3533 VCC.n3518 0.00942857
R52642 VCC.n3589 VCC.n3588 0.00942857
R52643 VCC.n4085 VCC.n4072 0.00942857
R52644 VCC.n4125 VCC.n4047 0.00942857
R52645 VCC.n4141 VCC.n4041 0.00942857
R52646 VCC.n4173 VCC.n4017 0.00942857
R52647 VCC.n4084 VCC.n4069 0.00942857
R52648 VCC.n4140 VCC.n4139 0.00942857
R52649 VCC.n4246 VCC.n3984 0.00942857
R52650 VCC.n4262 VCC.n3977 0.00942857
R52651 VCC.n3956 VCC.n3947 0.00942857
R52652 VCC.n4261 VCC.n3979 0.00942857
R52653 VCC.n3954 VCC.n3948 0.00942857
R52654 VCC.n4336 VCC.n4335 0.00942857
R52655 VCC.n4413 VCC.n3895 0.00942857
R52656 VCC.n3898 VCC.n3896 0.00942857
R52657 VCC.n4334 VCC.n3943 0.00942857
R52658 VCC.n4358 VCC.n3930 0.00942857
R52659 VCC.n4386 VCC.n4385 0.00942857
R52660 VCC.n3897 VCC.n3891 0.00942857
R52661 VCC.n4895 VCC.n4894 0.00942857
R52662 VCC.n4960 VCC.n4959 0.00942857
R52663 VCC.n4973 VCC.n4446 0.00942857
R52664 VCC.n4893 VCC.n4500 0.00942857
R52665 VCC.n4924 VCC.n4483 0.00942857
R52666 VCC.n4937 VCC.n4476 0.00942857
R52667 VCC.n4972 VCC.n4971 0.00942857
R52668 VCC.n4803 VCC.n4541 0.00942857
R52669 VCC.n4819 VCC.n4534 0.00942857
R52670 VCC.n4513 VCC.n4504 0.00942857
R52671 VCC.n4818 VCC.n4536 0.00942857
R52672 VCC.n4511 VCC.n4505 0.00942857
R52673 VCC.n4643 VCC.n4630 0.00942857
R52674 VCC.n4683 VCC.n4605 0.00942857
R52675 VCC.n4699 VCC.n4599 0.00942857
R52676 VCC.n4731 VCC.n4575 0.00942857
R52677 VCC.n4642 VCC.n4627 0.00942857
R52678 VCC.n4698 VCC.n4697 0.00942857
R52679 VCC.n5194 VCC.n5181 0.00942857
R52680 VCC.n5234 VCC.n5156 0.00942857
R52681 VCC.n5250 VCC.n5150 0.00942857
R52682 VCC.n5282 VCC.n5126 0.00942857
R52683 VCC.n5193 VCC.n5178 0.00942857
R52684 VCC.n5249 VCC.n5248 0.00942857
R52685 VCC.n5355 VCC.n5093 0.00942857
R52686 VCC.n5371 VCC.n5086 0.00942857
R52687 VCC.n5065 VCC.n5056 0.00942857
R52688 VCC.n5370 VCC.n5088 0.00942857
R52689 VCC.n5063 VCC.n5057 0.00942857
R52690 VCC.n5445 VCC.n5444 0.00942857
R52691 VCC.n5522 VCC.n5004 0.00942857
R52692 VCC.n5007 VCC.n5005 0.00942857
R52693 VCC.n5443 VCC.n5052 0.00942857
R52694 VCC.n5467 VCC.n5039 0.00942857
R52695 VCC.n5495 VCC.n5494 0.00942857
R52696 VCC.n5006 VCC.n5000 0.00942857
R52697 VCC.n6004 VCC.n6003 0.00942857
R52698 VCC.n6069 VCC.n6068 0.00942857
R52699 VCC.n6082 VCC.n5555 0.00942857
R52700 VCC.n6002 VCC.n5609 0.00942857
R52701 VCC.n6033 VCC.n5592 0.00942857
R52702 VCC.n6046 VCC.n5585 0.00942857
R52703 VCC.n6081 VCC.n6080 0.00942857
R52704 VCC.n5912 VCC.n5650 0.00942857
R52705 VCC.n5928 VCC.n5643 0.00942857
R52706 VCC.n5622 VCC.n5613 0.00942857
R52707 VCC.n5927 VCC.n5645 0.00942857
R52708 VCC.n5620 VCC.n5614 0.00942857
R52709 VCC.n5752 VCC.n5739 0.00942857
R52710 VCC.n5792 VCC.n5714 0.00942857
R52711 VCC.n5808 VCC.n5708 0.00942857
R52712 VCC.n5840 VCC.n5684 0.00942857
R52713 VCC.n5751 VCC.n5736 0.00942857
R52714 VCC.n5807 VCC.n5806 0.00942857
R52715 VCC.n6303 VCC.n6290 0.00942857
R52716 VCC.n6343 VCC.n6265 0.00942857
R52717 VCC.n6359 VCC.n6259 0.00942857
R52718 VCC.n6391 VCC.n6235 0.00942857
R52719 VCC.n6302 VCC.n6287 0.00942857
R52720 VCC.n6358 VCC.n6357 0.00942857
R52721 VCC.n6464 VCC.n6202 0.00942857
R52722 VCC.n6480 VCC.n6195 0.00942857
R52723 VCC.n6174 VCC.n6165 0.00942857
R52724 VCC.n6479 VCC.n6197 0.00942857
R52725 VCC.n6172 VCC.n6166 0.00942857
R52726 VCC.n6554 VCC.n6553 0.00942857
R52727 VCC.n6631 VCC.n6113 0.00942857
R52728 VCC.n6116 VCC.n6114 0.00942857
R52729 VCC.n6552 VCC.n6161 0.00942857
R52730 VCC.n6576 VCC.n6148 0.00942857
R52731 VCC.n6604 VCC.n6603 0.00942857
R52732 VCC.n6115 VCC.n6109 0.00942857
R52733 VCC.n7113 VCC.n7112 0.00942857
R52734 VCC.n7178 VCC.n7177 0.00942857
R52735 VCC.n7191 VCC.n6664 0.00942857
R52736 VCC.n7111 VCC.n6718 0.00942857
R52737 VCC.n7142 VCC.n6701 0.00942857
R52738 VCC.n7155 VCC.n6694 0.00942857
R52739 VCC.n7190 VCC.n7189 0.00942857
R52740 VCC.n7021 VCC.n6759 0.00942857
R52741 VCC.n7037 VCC.n6752 0.00942857
R52742 VCC.n6731 VCC.n6722 0.00942857
R52743 VCC.n7036 VCC.n6754 0.00942857
R52744 VCC.n6729 VCC.n6723 0.00942857
R52745 VCC.n6861 VCC.n6848 0.00942857
R52746 VCC.n6901 VCC.n6823 0.00942857
R52747 VCC.n6917 VCC.n6817 0.00942857
R52748 VCC.n6949 VCC.n6793 0.00942857
R52749 VCC.n6860 VCC.n6845 0.00942857
R52750 VCC.n6916 VCC.n6915 0.00942857
R52751 VCC.n7412 VCC.n7399 0.00942857
R52752 VCC.n7452 VCC.n7374 0.00942857
R52753 VCC.n7468 VCC.n7368 0.00942857
R52754 VCC.n7500 VCC.n7344 0.00942857
R52755 VCC.n7411 VCC.n7396 0.00942857
R52756 VCC.n7467 VCC.n7466 0.00942857
R52757 VCC.n7573 VCC.n7311 0.00942857
R52758 VCC.n7589 VCC.n7304 0.00942857
R52759 VCC.n7283 VCC.n7274 0.00942857
R52760 VCC.n7588 VCC.n7306 0.00942857
R52761 VCC.n7281 VCC.n7275 0.00942857
R52762 VCC.n7663 VCC.n7662 0.00942857
R52763 VCC.n7740 VCC.n7222 0.00942857
R52764 VCC.n7225 VCC.n7223 0.00942857
R52765 VCC.n7661 VCC.n7270 0.00942857
R52766 VCC.n7685 VCC.n7257 0.00942857
R52767 VCC.n7713 VCC.n7712 0.00942857
R52768 VCC.n7224 VCC.n7218 0.00942857
R52769 VCC.n8222 VCC.n8221 0.00942857
R52770 VCC.n8287 VCC.n8286 0.00942857
R52771 VCC.n8300 VCC.n7773 0.00942857
R52772 VCC.n8220 VCC.n7827 0.00942857
R52773 VCC.n8251 VCC.n7810 0.00942857
R52774 VCC.n8264 VCC.n7803 0.00942857
R52775 VCC.n8299 VCC.n8298 0.00942857
R52776 VCC.n8130 VCC.n7868 0.00942857
R52777 VCC.n8146 VCC.n7861 0.00942857
R52778 VCC.n7840 VCC.n7831 0.00942857
R52779 VCC.n8145 VCC.n7863 0.00942857
R52780 VCC.n7838 VCC.n7832 0.00942857
R52781 VCC.n7970 VCC.n7957 0.00942857
R52782 VCC.n8010 VCC.n7932 0.00942857
R52783 VCC.n8026 VCC.n7926 0.00942857
R52784 VCC.n8058 VCC.n7902 0.00942857
R52785 VCC.n7969 VCC.n7954 0.00942857
R52786 VCC.n8025 VCC.n8024 0.00942857
R52787 VCC.n8682 VCC.n8420 0.00942857
R52788 VCC.n8698 VCC.n8413 0.00942857
R52789 VCC.n8392 VCC.n8383 0.00942857
R52790 VCC.n8697 VCC.n8415 0.00942857
R52791 VCC.n8390 VCC.n8384 0.00942857
R52792 VCC.n8772 VCC.n8771 0.00942857
R52793 VCC.n8849 VCC.n8331 0.00942857
R52794 VCC.n8334 VCC.n8332 0.00942857
R52795 VCC.n8770 VCC.n8379 0.00942857
R52796 VCC.n8794 VCC.n8366 0.00942857
R52797 VCC.n8822 VCC.n8821 0.00942857
R52798 VCC.n8333 VCC.n8327 0.00942857
R52799 VCC.n8521 VCC.n8508 0.00942857
R52800 VCC.n8561 VCC.n8483 0.00942857
R52801 VCC.n8577 VCC.n8477 0.00942857
R52802 VCC.n8609 VCC.n8453 0.00942857
R52803 VCC.n8520 VCC.n8505 0.00942857
R52804 VCC.n8576 VCC.n8575 0.00942857
R52805 VCC.n9331 VCC.n9330 0.00942857
R52806 VCC.n9396 VCC.n9395 0.00942857
R52807 VCC.n9409 VCC.n8882 0.00942857
R52808 VCC.n9329 VCC.n8936 0.00942857
R52809 VCC.n9360 VCC.n8919 0.00942857
R52810 VCC.n9373 VCC.n8912 0.00942857
R52811 VCC.n9408 VCC.n9407 0.00942857
R52812 VCC.n9239 VCC.n8977 0.00942857
R52813 VCC.n9255 VCC.n8970 0.00942857
R52814 VCC.n8949 VCC.n8940 0.00942857
R52815 VCC.n9254 VCC.n8972 0.00942857
R52816 VCC.n8947 VCC.n8941 0.00942857
R52817 VCC.n9079 VCC.n9066 0.00942857
R52818 VCC.n9119 VCC.n9041 0.00942857
R52819 VCC.n9135 VCC.n9035 0.00942857
R52820 VCC.n9167 VCC.n9011 0.00942857
R52821 VCC.n9078 VCC.n9063 0.00942857
R52822 VCC.n9134 VCC.n9133 0.00942857
R52823 VCC.n9630 VCC.n9617 0.00942857
R52824 VCC.n9670 VCC.n9592 0.00942857
R52825 VCC.n9686 VCC.n9586 0.00942857
R52826 VCC.n9718 VCC.n9562 0.00942857
R52827 VCC.n9629 VCC.n9614 0.00942857
R52828 VCC.n9685 VCC.n9684 0.00942857
R52829 VCC.n9791 VCC.n9529 0.00942857
R52830 VCC.n9807 VCC.n9522 0.00942857
R52831 VCC.n9501 VCC.n9492 0.00942857
R52832 VCC.n9806 VCC.n9524 0.00942857
R52833 VCC.n9499 VCC.n9493 0.00942857
R52834 VCC.n9881 VCC.n9880 0.00942857
R52835 VCC.n9958 VCC.n9440 0.00942857
R52836 VCC.n9443 VCC.n9441 0.00942857
R52837 VCC.n9879 VCC.n9488 0.00942857
R52838 VCC.n9903 VCC.n9475 0.00942857
R52839 VCC.n9931 VCC.n9930 0.00942857
R52840 VCC.n9442 VCC.n9436 0.00942857
R52841 VCC.n10439 VCC.n10438 0.00942857
R52842 VCC.n10504 VCC.n10503 0.00942857
R52843 VCC.n10517 VCC.n9990 0.00942857
R52844 VCC.n10437 VCC.n10044 0.00942857
R52845 VCC.n10468 VCC.n10027 0.00942857
R52846 VCC.n10481 VCC.n10020 0.00942857
R52847 VCC.n10516 VCC.n10515 0.00942857
R52848 VCC.n10347 VCC.n10085 0.00942857
R52849 VCC.n10363 VCC.n10078 0.00942857
R52850 VCC.n10057 VCC.n10048 0.00942857
R52851 VCC.n10362 VCC.n10080 0.00942857
R52852 VCC.n10055 VCC.n10049 0.00942857
R52853 VCC.n10187 VCC.n10174 0.00942857
R52854 VCC.n10227 VCC.n10149 0.00942857
R52855 VCC.n10243 VCC.n10143 0.00942857
R52856 VCC.n10275 VCC.n10119 0.00942857
R52857 VCC.n10186 VCC.n10171 0.00942857
R52858 VCC.n10242 VCC.n10241 0.00942857
R52859 VCC.n10737 VCC.n10724 0.00942857
R52860 VCC.n10777 VCC.n10699 0.00942857
R52861 VCC.n10793 VCC.n10693 0.00942857
R52862 VCC.n10825 VCC.n10669 0.00942857
R52863 VCC.n10736 VCC.n10721 0.00942857
R52864 VCC.n10792 VCC.n10791 0.00942857
R52865 VCC.n10898 VCC.n10636 0.00942857
R52866 VCC.n10914 VCC.n10629 0.00942857
R52867 VCC.n10608 VCC.n10599 0.00942857
R52868 VCC.n10913 VCC.n10631 0.00942857
R52869 VCC.n10606 VCC.n10600 0.00942857
R52870 VCC.n10988 VCC.n10987 0.00942857
R52871 VCC.n11065 VCC.n10547 0.00942857
R52872 VCC.n10550 VCC.n10548 0.00942857
R52873 VCC.n10986 VCC.n10595 0.00942857
R52874 VCC.n11010 VCC.n10582 0.00942857
R52875 VCC.n11038 VCC.n11037 0.00942857
R52876 VCC.n10549 VCC.n10543 0.00942857
R52877 VCC.n11546 VCC.n11545 0.00942857
R52878 VCC.n11611 VCC.n11610 0.00942857
R52879 VCC.n11624 VCC.n11097 0.00942857
R52880 VCC.n11544 VCC.n11151 0.00942857
R52881 VCC.n11575 VCC.n11134 0.00942857
R52882 VCC.n11588 VCC.n11127 0.00942857
R52883 VCC.n11623 VCC.n11622 0.00942857
R52884 VCC.n11454 VCC.n11192 0.00942857
R52885 VCC.n11470 VCC.n11185 0.00942857
R52886 VCC.n11164 VCC.n11155 0.00942857
R52887 VCC.n11469 VCC.n11187 0.00942857
R52888 VCC.n11162 VCC.n11156 0.00942857
R52889 VCC.n11294 VCC.n11281 0.00942857
R52890 VCC.n11334 VCC.n11256 0.00942857
R52891 VCC.n11350 VCC.n11250 0.00942857
R52892 VCC.n11382 VCC.n11226 0.00942857
R52893 VCC.n11293 VCC.n11278 0.00942857
R52894 VCC.n11349 VCC.n11348 0.00942857
R52895 VCC.n11844 VCC.n11831 0.00942857
R52896 VCC.n11884 VCC.n11806 0.00942857
R52897 VCC.n11900 VCC.n11800 0.00942857
R52898 VCC.n11932 VCC.n11776 0.00942857
R52899 VCC.n11843 VCC.n11828 0.00942857
R52900 VCC.n11899 VCC.n11898 0.00942857
R52901 VCC.n12005 VCC.n11743 0.00942857
R52902 VCC.n12021 VCC.n11736 0.00942857
R52903 VCC.n11715 VCC.n11706 0.00942857
R52904 VCC.n12020 VCC.n11738 0.00942857
R52905 VCC.n11713 VCC.n11707 0.00942857
R52906 VCC.n12095 VCC.n12094 0.00942857
R52907 VCC.n12172 VCC.n11654 0.00942857
R52908 VCC.n11657 VCC.n11655 0.00942857
R52909 VCC.n12093 VCC.n11702 0.00942857
R52910 VCC.n12117 VCC.n11689 0.00942857
R52911 VCC.n12145 VCC.n12144 0.00942857
R52912 VCC.n11656 VCC.n11650 0.00942857
R52913 VCC.n12653 VCC.n12652 0.00942857
R52914 VCC.n12718 VCC.n12717 0.00942857
R52915 VCC.n12731 VCC.n12204 0.00942857
R52916 VCC.n12651 VCC.n12258 0.00942857
R52917 VCC.n12682 VCC.n12241 0.00942857
R52918 VCC.n12695 VCC.n12234 0.00942857
R52919 VCC.n12730 VCC.n12729 0.00942857
R52920 VCC.n12561 VCC.n12299 0.00942857
R52921 VCC.n12577 VCC.n12292 0.00942857
R52922 VCC.n12271 VCC.n12262 0.00942857
R52923 VCC.n12576 VCC.n12294 0.00942857
R52924 VCC.n12269 VCC.n12263 0.00942857
R52925 VCC.n12401 VCC.n12388 0.00942857
R52926 VCC.n12441 VCC.n12363 0.00942857
R52927 VCC.n12457 VCC.n12357 0.00942857
R52928 VCC.n12489 VCC.n12333 0.00942857
R52929 VCC.n12400 VCC.n12385 0.00942857
R52930 VCC.n12456 VCC.n12455 0.00942857
R52931 VCC.n12951 VCC.n12938 0.00942857
R52932 VCC.n12991 VCC.n12913 0.00942857
R52933 VCC.n13007 VCC.n12907 0.00942857
R52934 VCC.n13039 VCC.n12883 0.00942857
R52935 VCC.n12950 VCC.n12935 0.00942857
R52936 VCC.n13006 VCC.n13005 0.00942857
R52937 VCC.n13112 VCC.n12850 0.00942857
R52938 VCC.n13128 VCC.n12843 0.00942857
R52939 VCC.n12822 VCC.n12813 0.00942857
R52940 VCC.n13127 VCC.n12845 0.00942857
R52941 VCC.n12820 VCC.n12814 0.00942857
R52942 VCC.n13202 VCC.n13201 0.00942857
R52943 VCC.n13279 VCC.n12761 0.00942857
R52944 VCC.n12764 VCC.n12762 0.00942857
R52945 VCC.n13200 VCC.n12809 0.00942857
R52946 VCC.n13224 VCC.n12796 0.00942857
R52947 VCC.n13252 VCC.n13251 0.00942857
R52948 VCC.n12763 VCC.n12757 0.00942857
R52949 VCC.n13760 VCC.n13759 0.00942857
R52950 VCC.n13825 VCC.n13824 0.00942857
R52951 VCC.n13838 VCC.n13311 0.00942857
R52952 VCC.n13758 VCC.n13365 0.00942857
R52953 VCC.n13789 VCC.n13348 0.00942857
R52954 VCC.n13802 VCC.n13341 0.00942857
R52955 VCC.n13837 VCC.n13836 0.00942857
R52956 VCC.n13668 VCC.n13406 0.00942857
R52957 VCC.n13684 VCC.n13399 0.00942857
R52958 VCC.n13378 VCC.n13369 0.00942857
R52959 VCC.n13683 VCC.n13401 0.00942857
R52960 VCC.n13376 VCC.n13370 0.00942857
R52961 VCC.n13508 VCC.n13495 0.00942857
R52962 VCC.n13548 VCC.n13470 0.00942857
R52963 VCC.n13564 VCC.n13464 0.00942857
R52964 VCC.n13596 VCC.n13440 0.00942857
R52965 VCC.n13507 VCC.n13492 0.00942857
R52966 VCC.n13563 VCC.n13562 0.00942857
R52967 VCC.n14058 VCC.n14045 0.00942857
R52968 VCC.n14098 VCC.n14020 0.00942857
R52969 VCC.n14114 VCC.n14014 0.00942857
R52970 VCC.n14146 VCC.n13990 0.00942857
R52971 VCC.n14057 VCC.n14042 0.00942857
R52972 VCC.n14113 VCC.n14112 0.00942857
R52973 VCC.n14219 VCC.n13957 0.00942857
R52974 VCC.n14235 VCC.n13950 0.00942857
R52975 VCC.n13929 VCC.n13920 0.00942857
R52976 VCC.n14234 VCC.n13952 0.00942857
R52977 VCC.n13927 VCC.n13921 0.00942857
R52978 VCC.n14309 VCC.n14308 0.00942857
R52979 VCC.n14386 VCC.n13868 0.00942857
R52980 VCC.n13871 VCC.n13869 0.00942857
R52981 VCC.n14307 VCC.n13916 0.00942857
R52982 VCC.n14331 VCC.n13903 0.00942857
R52983 VCC.n14359 VCC.n14358 0.00942857
R52984 VCC.n13870 VCC.n13864 0.00942857
R52985 VCC.n14867 VCC.n14866 0.00942857
R52986 VCC.n14932 VCC.n14931 0.00942857
R52987 VCC.n14945 VCC.n14418 0.00942857
R52988 VCC.n14865 VCC.n14472 0.00942857
R52989 VCC.n14896 VCC.n14455 0.00942857
R52990 VCC.n14909 VCC.n14448 0.00942857
R52991 VCC.n14944 VCC.n14943 0.00942857
R52992 VCC.n14775 VCC.n14513 0.00942857
R52993 VCC.n14791 VCC.n14506 0.00942857
R52994 VCC.n14485 VCC.n14476 0.00942857
R52995 VCC.n14790 VCC.n14508 0.00942857
R52996 VCC.n14483 VCC.n14477 0.00942857
R52997 VCC.n14615 VCC.n14602 0.00942857
R52998 VCC.n14655 VCC.n14577 0.00942857
R52999 VCC.n14671 VCC.n14571 0.00942857
R53000 VCC.n14703 VCC.n14547 0.00942857
R53001 VCC.n14614 VCC.n14599 0.00942857
R53002 VCC.n14670 VCC.n14669 0.00942857
R53003 VCC.n15165 VCC.n15152 0.00942857
R53004 VCC.n15205 VCC.n15127 0.00942857
R53005 VCC.n15221 VCC.n15121 0.00942857
R53006 VCC.n15253 VCC.n15097 0.00942857
R53007 VCC.n15164 VCC.n15149 0.00942857
R53008 VCC.n15220 VCC.n15219 0.00942857
R53009 VCC.n15326 VCC.n15064 0.00942857
R53010 VCC.n15342 VCC.n15057 0.00942857
R53011 VCC.n15036 VCC.n15027 0.00942857
R53012 VCC.n15341 VCC.n15059 0.00942857
R53013 VCC.n15034 VCC.n15028 0.00942857
R53014 VCC.n15416 VCC.n15415 0.00942857
R53015 VCC.n15493 VCC.n14975 0.00942857
R53016 VCC.n14978 VCC.n14976 0.00942857
R53017 VCC.n15414 VCC.n15023 0.00942857
R53018 VCC.n15438 VCC.n15010 0.00942857
R53019 VCC.n15466 VCC.n15465 0.00942857
R53020 VCC.n14977 VCC.n14971 0.00942857
R53021 VCC.n15974 VCC.n15973 0.00942857
R53022 VCC.n16039 VCC.n16038 0.00942857
R53023 VCC.n16052 VCC.n15525 0.00942857
R53024 VCC.n15972 VCC.n15579 0.00942857
R53025 VCC.n16003 VCC.n15562 0.00942857
R53026 VCC.n16016 VCC.n15555 0.00942857
R53027 VCC.n16051 VCC.n16050 0.00942857
R53028 VCC.n15882 VCC.n15620 0.00942857
R53029 VCC.n15898 VCC.n15613 0.00942857
R53030 VCC.n15592 VCC.n15583 0.00942857
R53031 VCC.n15897 VCC.n15615 0.00942857
R53032 VCC.n15590 VCC.n15584 0.00942857
R53033 VCC.n15722 VCC.n15709 0.00942857
R53034 VCC.n15762 VCC.n15684 0.00942857
R53035 VCC.n15778 VCC.n15678 0.00942857
R53036 VCC.n15810 VCC.n15654 0.00942857
R53037 VCC.n15721 VCC.n15706 0.00942857
R53038 VCC.n15777 VCC.n15776 0.00942857
R53039 VCC.n16272 VCC.n16259 0.00942857
R53040 VCC.n16312 VCC.n16234 0.00942857
R53041 VCC.n16328 VCC.n16228 0.00942857
R53042 VCC.n16360 VCC.n16204 0.00942857
R53043 VCC.n16271 VCC.n16256 0.00942857
R53044 VCC.n16327 VCC.n16326 0.00942857
R53045 VCC.n16433 VCC.n16171 0.00942857
R53046 VCC.n16449 VCC.n16164 0.00942857
R53047 VCC.n16143 VCC.n16134 0.00942857
R53048 VCC.n16448 VCC.n16166 0.00942857
R53049 VCC.n16141 VCC.n16135 0.00942857
R53050 VCC.n16523 VCC.n16522 0.00942857
R53051 VCC.n16600 VCC.n16082 0.00942857
R53052 VCC.n16085 VCC.n16083 0.00942857
R53053 VCC.n16521 VCC.n16130 0.00942857
R53054 VCC.n16545 VCC.n16117 0.00942857
R53055 VCC.n16573 VCC.n16572 0.00942857
R53056 VCC.n16084 VCC.n16078 0.00942857
R53057 VCC.n17081 VCC.n17080 0.00942857
R53058 VCC.n17146 VCC.n17145 0.00942857
R53059 VCC.n17159 VCC.n16632 0.00942857
R53060 VCC.n17079 VCC.n16686 0.00942857
R53061 VCC.n17110 VCC.n16669 0.00942857
R53062 VCC.n17123 VCC.n16662 0.00942857
R53063 VCC.n17158 VCC.n17157 0.00942857
R53064 VCC.n16989 VCC.n16727 0.00942857
R53065 VCC.n17005 VCC.n16720 0.00942857
R53066 VCC.n16699 VCC.n16690 0.00942857
R53067 VCC.n17004 VCC.n16722 0.00942857
R53068 VCC.n16697 VCC.n16691 0.00942857
R53069 VCC.n16829 VCC.n16816 0.00942857
R53070 VCC.n16869 VCC.n16791 0.00942857
R53071 VCC.n16885 VCC.n16785 0.00942857
R53072 VCC.n16917 VCC.n16761 0.00942857
R53073 VCC.n16828 VCC.n16813 0.00942857
R53074 VCC.n16884 VCC.n16883 0.00942857
R53075 VCC.n17353 VCC.n17278 0.00942857
R53076 VCC.n17369 VCC.n17271 0.00942857
R53077 VCC.n17250 VCC.n17241 0.00942857
R53078 VCC.n17368 VCC.n17273 0.00942857
R53079 VCC.n17248 VCC.n17242 0.00942857
R53080 VCC.n17443 VCC.n17442 0.00942857
R53081 VCC.n17520 VCC.n17189 0.00942857
R53082 VCC.n17192 VCC.n17190 0.00942857
R53083 VCC.n17441 VCC.n17237 0.00942857
R53084 VCC.n17465 VCC.n17224 0.00942857
R53085 VCC.n17493 VCC.n17492 0.00942857
R53086 VCC.n17191 VCC.n17185 0.00942857
R53087 VCC.n222 VCC.n221 0.00853571
R53088 VCC.n233 VCC.n176 0.00853571
R53089 VCC.n251 VCC.n250 0.00853571
R53090 VCC.n284 VCC.n145 0.00853571
R53091 VCC.n172 VCC.n166 0.00853571
R53092 VCC.n342 VCC.n117 0.00853571
R53093 VCC.n356 VCC.n111 0.00853571
R53094 VCC.n388 VCC.n96 0.00853571
R53095 VCC.n411 VCC.n85 0.00853571
R53096 VCC.n375 VCC.n374 0.00853571
R53097 VCC.n478 VCC.n52 0.00853571
R53098 VCC.n540 VCC.n539 0.00853571
R53099 VCC.n551 VCC.n1 0.00853571
R53100 VCC.n774 VCC.n773 0.00853571
R53101 VCC.n785 VCC.n728 0.00853571
R53102 VCC.n803 VCC.n802 0.00853571
R53103 VCC.n836 VCC.n697 0.00853571
R53104 VCC.n724 VCC.n718 0.00853571
R53105 VCC.n894 VCC.n669 0.00853571
R53106 VCC.n908 VCC.n663 0.00853571
R53107 VCC.n940 VCC.n648 0.00853571
R53108 VCC.n963 VCC.n637 0.00853571
R53109 VCC.n927 VCC.n926 0.00853571
R53110 VCC.n1030 VCC.n604 0.00853571
R53111 VCC.n1094 VCC.n1093 0.00853571
R53112 VCC.n1105 VCC.n555 0.00853571
R53113 VCC.n1596 VCC.n1157 0.00853571
R53114 VCC.n1638 VCC.n1121 0.00853571
R53115 VCC.n1659 VCC.n1109 0.00853571
R53116 VCC.n1451 VCC.n1226 0.00853571
R53117 VCC.n1465 VCC.n1220 0.00853571
R53118 VCC.n1497 VCC.n1205 0.00853571
R53119 VCC.n1520 VCC.n1194 0.00853571
R53120 VCC.n1484 VCC.n1483 0.00853571
R53121 VCC.n1332 VCC.n1331 0.00853571
R53122 VCC.n1343 VCC.n1286 0.00853571
R53123 VCC.n1361 VCC.n1360 0.00853571
R53124 VCC.n1394 VCC.n1255 0.00853571
R53125 VCC.n1282 VCC.n1276 0.00853571
R53126 VCC.n1883 VCC.n1882 0.00853571
R53127 VCC.n1894 VCC.n1837 0.00853571
R53128 VCC.n1912 VCC.n1911 0.00853571
R53129 VCC.n1945 VCC.n1806 0.00853571
R53130 VCC.n1833 VCC.n1827 0.00853571
R53131 VCC.n2003 VCC.n1778 0.00853571
R53132 VCC.n2017 VCC.n1772 0.00853571
R53133 VCC.n2049 VCC.n1757 0.00853571
R53134 VCC.n2072 VCC.n1746 0.00853571
R53135 VCC.n2036 VCC.n2035 0.00853571
R53136 VCC.n2139 VCC.n1713 0.00853571
R53137 VCC.n2203 VCC.n2202 0.00853571
R53138 VCC.n2214 VCC.n1664 0.00853571
R53139 VCC.n2705 VCC.n2266 0.00853571
R53140 VCC.n2747 VCC.n2230 0.00853571
R53141 VCC.n2768 VCC.n2218 0.00853571
R53142 VCC.n2560 VCC.n2335 0.00853571
R53143 VCC.n2574 VCC.n2329 0.00853571
R53144 VCC.n2606 VCC.n2314 0.00853571
R53145 VCC.n2629 VCC.n2303 0.00853571
R53146 VCC.n2593 VCC.n2592 0.00853571
R53147 VCC.n2441 VCC.n2440 0.00853571
R53148 VCC.n2452 VCC.n2395 0.00853571
R53149 VCC.n2470 VCC.n2469 0.00853571
R53150 VCC.n2503 VCC.n2364 0.00853571
R53151 VCC.n2391 VCC.n2385 0.00853571
R53152 VCC.n2992 VCC.n2991 0.00853571
R53153 VCC.n3003 VCC.n2946 0.00853571
R53154 VCC.n3021 VCC.n3020 0.00853571
R53155 VCC.n3054 VCC.n2915 0.00853571
R53156 VCC.n2942 VCC.n2936 0.00853571
R53157 VCC.n3112 VCC.n2887 0.00853571
R53158 VCC.n3126 VCC.n2881 0.00853571
R53159 VCC.n3158 VCC.n2866 0.00853571
R53160 VCC.n3181 VCC.n2855 0.00853571
R53161 VCC.n3145 VCC.n3144 0.00853571
R53162 VCC.n3248 VCC.n2822 0.00853571
R53163 VCC.n3312 VCC.n3311 0.00853571
R53164 VCC.n3323 VCC.n2773 0.00853571
R53165 VCC.n3814 VCC.n3375 0.00853571
R53166 VCC.n3856 VCC.n3339 0.00853571
R53167 VCC.n3877 VCC.n3327 0.00853571
R53168 VCC.n3669 VCC.n3444 0.00853571
R53169 VCC.n3683 VCC.n3438 0.00853571
R53170 VCC.n3715 VCC.n3423 0.00853571
R53171 VCC.n3738 VCC.n3412 0.00853571
R53172 VCC.n3702 VCC.n3701 0.00853571
R53173 VCC.n3550 VCC.n3549 0.00853571
R53174 VCC.n3561 VCC.n3504 0.00853571
R53175 VCC.n3579 VCC.n3578 0.00853571
R53176 VCC.n3612 VCC.n3473 0.00853571
R53177 VCC.n3500 VCC.n3494 0.00853571
R53178 VCC.n4101 VCC.n4100 0.00853571
R53179 VCC.n4112 VCC.n4055 0.00853571
R53180 VCC.n4130 VCC.n4129 0.00853571
R53181 VCC.n4163 VCC.n4024 0.00853571
R53182 VCC.n4051 VCC.n4045 0.00853571
R53183 VCC.n4221 VCC.n3996 0.00853571
R53184 VCC.n4235 VCC.n3990 0.00853571
R53185 VCC.n4267 VCC.n3975 0.00853571
R53186 VCC.n4290 VCC.n3964 0.00853571
R53187 VCC.n4254 VCC.n4253 0.00853571
R53188 VCC.n4357 VCC.n3931 0.00853571
R53189 VCC.n4421 VCC.n4420 0.00853571
R53190 VCC.n4432 VCC.n3882 0.00853571
R53191 VCC.n4923 VCC.n4484 0.00853571
R53192 VCC.n4965 VCC.n4448 0.00853571
R53193 VCC.n4986 VCC.n4436 0.00853571
R53194 VCC.n4778 VCC.n4553 0.00853571
R53195 VCC.n4792 VCC.n4547 0.00853571
R53196 VCC.n4824 VCC.n4532 0.00853571
R53197 VCC.n4847 VCC.n4521 0.00853571
R53198 VCC.n4811 VCC.n4810 0.00853571
R53199 VCC.n4659 VCC.n4658 0.00853571
R53200 VCC.n4670 VCC.n4613 0.00853571
R53201 VCC.n4688 VCC.n4687 0.00853571
R53202 VCC.n4721 VCC.n4582 0.00853571
R53203 VCC.n4609 VCC.n4603 0.00853571
R53204 VCC.n5210 VCC.n5209 0.00853571
R53205 VCC.n5221 VCC.n5164 0.00853571
R53206 VCC.n5239 VCC.n5238 0.00853571
R53207 VCC.n5272 VCC.n5133 0.00853571
R53208 VCC.n5160 VCC.n5154 0.00853571
R53209 VCC.n5330 VCC.n5105 0.00853571
R53210 VCC.n5344 VCC.n5099 0.00853571
R53211 VCC.n5376 VCC.n5084 0.00853571
R53212 VCC.n5399 VCC.n5073 0.00853571
R53213 VCC.n5363 VCC.n5362 0.00853571
R53214 VCC.n5466 VCC.n5040 0.00853571
R53215 VCC.n5530 VCC.n5529 0.00853571
R53216 VCC.n5541 VCC.n4991 0.00853571
R53217 VCC.n6032 VCC.n5593 0.00853571
R53218 VCC.n6074 VCC.n5557 0.00853571
R53219 VCC.n6095 VCC.n5545 0.00853571
R53220 VCC.n5887 VCC.n5662 0.00853571
R53221 VCC.n5901 VCC.n5656 0.00853571
R53222 VCC.n5933 VCC.n5641 0.00853571
R53223 VCC.n5956 VCC.n5630 0.00853571
R53224 VCC.n5920 VCC.n5919 0.00853571
R53225 VCC.n5768 VCC.n5767 0.00853571
R53226 VCC.n5779 VCC.n5722 0.00853571
R53227 VCC.n5797 VCC.n5796 0.00853571
R53228 VCC.n5830 VCC.n5691 0.00853571
R53229 VCC.n5718 VCC.n5712 0.00853571
R53230 VCC.n6319 VCC.n6318 0.00853571
R53231 VCC.n6330 VCC.n6273 0.00853571
R53232 VCC.n6348 VCC.n6347 0.00853571
R53233 VCC.n6381 VCC.n6242 0.00853571
R53234 VCC.n6269 VCC.n6263 0.00853571
R53235 VCC.n6439 VCC.n6214 0.00853571
R53236 VCC.n6453 VCC.n6208 0.00853571
R53237 VCC.n6485 VCC.n6193 0.00853571
R53238 VCC.n6508 VCC.n6182 0.00853571
R53239 VCC.n6472 VCC.n6471 0.00853571
R53240 VCC.n6575 VCC.n6149 0.00853571
R53241 VCC.n6639 VCC.n6638 0.00853571
R53242 VCC.n6650 VCC.n6100 0.00853571
R53243 VCC.n7141 VCC.n6702 0.00853571
R53244 VCC.n7183 VCC.n6666 0.00853571
R53245 VCC.n7204 VCC.n6654 0.00853571
R53246 VCC.n6996 VCC.n6771 0.00853571
R53247 VCC.n7010 VCC.n6765 0.00853571
R53248 VCC.n7042 VCC.n6750 0.00853571
R53249 VCC.n7065 VCC.n6739 0.00853571
R53250 VCC.n7029 VCC.n7028 0.00853571
R53251 VCC.n6877 VCC.n6876 0.00853571
R53252 VCC.n6888 VCC.n6831 0.00853571
R53253 VCC.n6906 VCC.n6905 0.00853571
R53254 VCC.n6939 VCC.n6800 0.00853571
R53255 VCC.n6827 VCC.n6821 0.00853571
R53256 VCC.n7428 VCC.n7427 0.00853571
R53257 VCC.n7439 VCC.n7382 0.00853571
R53258 VCC.n7457 VCC.n7456 0.00853571
R53259 VCC.n7490 VCC.n7351 0.00853571
R53260 VCC.n7378 VCC.n7372 0.00853571
R53261 VCC.n7548 VCC.n7323 0.00853571
R53262 VCC.n7562 VCC.n7317 0.00853571
R53263 VCC.n7594 VCC.n7302 0.00853571
R53264 VCC.n7617 VCC.n7291 0.00853571
R53265 VCC.n7581 VCC.n7580 0.00853571
R53266 VCC.n7684 VCC.n7258 0.00853571
R53267 VCC.n7748 VCC.n7747 0.00853571
R53268 VCC.n7759 VCC.n7209 0.00853571
R53269 VCC.n8250 VCC.n7811 0.00853571
R53270 VCC.n8292 VCC.n7775 0.00853571
R53271 VCC.n8313 VCC.n7763 0.00853571
R53272 VCC.n8105 VCC.n7880 0.00853571
R53273 VCC.n8119 VCC.n7874 0.00853571
R53274 VCC.n8151 VCC.n7859 0.00853571
R53275 VCC.n8174 VCC.n7848 0.00853571
R53276 VCC.n8138 VCC.n8137 0.00853571
R53277 VCC.n7986 VCC.n7985 0.00853571
R53278 VCC.n7997 VCC.n7940 0.00853571
R53279 VCC.n8015 VCC.n8014 0.00853571
R53280 VCC.n8048 VCC.n7909 0.00853571
R53281 VCC.n7936 VCC.n7930 0.00853571
R53282 VCC.n8657 VCC.n8432 0.00853571
R53283 VCC.n8671 VCC.n8426 0.00853571
R53284 VCC.n8703 VCC.n8411 0.00853571
R53285 VCC.n8726 VCC.n8400 0.00853571
R53286 VCC.n8690 VCC.n8689 0.00853571
R53287 VCC.n8793 VCC.n8367 0.00853571
R53288 VCC.n8857 VCC.n8856 0.00853571
R53289 VCC.n8868 VCC.n8318 0.00853571
R53290 VCC.n8537 VCC.n8536 0.00853571
R53291 VCC.n8548 VCC.n8491 0.00853571
R53292 VCC.n8566 VCC.n8565 0.00853571
R53293 VCC.n8599 VCC.n8460 0.00853571
R53294 VCC.n8487 VCC.n8481 0.00853571
R53295 VCC.n9359 VCC.n8920 0.00853571
R53296 VCC.n9401 VCC.n8884 0.00853571
R53297 VCC.n9422 VCC.n8872 0.00853571
R53298 VCC.n9214 VCC.n8989 0.00853571
R53299 VCC.n9228 VCC.n8983 0.00853571
R53300 VCC.n9260 VCC.n8968 0.00853571
R53301 VCC.n9283 VCC.n8957 0.00853571
R53302 VCC.n9247 VCC.n9246 0.00853571
R53303 VCC.n9095 VCC.n9094 0.00853571
R53304 VCC.n9106 VCC.n9049 0.00853571
R53305 VCC.n9124 VCC.n9123 0.00853571
R53306 VCC.n9157 VCC.n9018 0.00853571
R53307 VCC.n9045 VCC.n9039 0.00853571
R53308 VCC.n9646 VCC.n9645 0.00853571
R53309 VCC.n9657 VCC.n9600 0.00853571
R53310 VCC.n9675 VCC.n9674 0.00853571
R53311 VCC.n9708 VCC.n9569 0.00853571
R53312 VCC.n9596 VCC.n9590 0.00853571
R53313 VCC.n9766 VCC.n9541 0.00853571
R53314 VCC.n9780 VCC.n9535 0.00853571
R53315 VCC.n9812 VCC.n9520 0.00853571
R53316 VCC.n9835 VCC.n9509 0.00853571
R53317 VCC.n9799 VCC.n9798 0.00853571
R53318 VCC.n9902 VCC.n9476 0.00853571
R53319 VCC.n9966 VCC.n9965 0.00853571
R53320 VCC.n9977 VCC.n9427 0.00853571
R53321 VCC.n10467 VCC.n10028 0.00853571
R53322 VCC.n10509 VCC.n9992 0.00853571
R53323 VCC.n10530 VCC.n9980 0.00853571
R53324 VCC.n10322 VCC.n10097 0.00853571
R53325 VCC.n10336 VCC.n10091 0.00853571
R53326 VCC.n10368 VCC.n10076 0.00853571
R53327 VCC.n10391 VCC.n10065 0.00853571
R53328 VCC.n10355 VCC.n10354 0.00853571
R53329 VCC.n10203 VCC.n10202 0.00853571
R53330 VCC.n10214 VCC.n10157 0.00853571
R53331 VCC.n10232 VCC.n10231 0.00853571
R53332 VCC.n10265 VCC.n10126 0.00853571
R53333 VCC.n10153 VCC.n10147 0.00853571
R53334 VCC.n10753 VCC.n10752 0.00853571
R53335 VCC.n10764 VCC.n10707 0.00853571
R53336 VCC.n10782 VCC.n10781 0.00853571
R53337 VCC.n10815 VCC.n10676 0.00853571
R53338 VCC.n10703 VCC.n10697 0.00853571
R53339 VCC.n10873 VCC.n10648 0.00853571
R53340 VCC.n10887 VCC.n10642 0.00853571
R53341 VCC.n10919 VCC.n10627 0.00853571
R53342 VCC.n10942 VCC.n10616 0.00853571
R53343 VCC.n10906 VCC.n10905 0.00853571
R53344 VCC.n11009 VCC.n10583 0.00853571
R53345 VCC.n11073 VCC.n11072 0.00853571
R53346 VCC.n11084 VCC.n10534 0.00853571
R53347 VCC.n11574 VCC.n11135 0.00853571
R53348 VCC.n11616 VCC.n11099 0.00853571
R53349 VCC.n11637 VCC.n11087 0.00853571
R53350 VCC.n11429 VCC.n11204 0.00853571
R53351 VCC.n11443 VCC.n11198 0.00853571
R53352 VCC.n11475 VCC.n11183 0.00853571
R53353 VCC.n11498 VCC.n11172 0.00853571
R53354 VCC.n11462 VCC.n11461 0.00853571
R53355 VCC.n11310 VCC.n11309 0.00853571
R53356 VCC.n11321 VCC.n11264 0.00853571
R53357 VCC.n11339 VCC.n11338 0.00853571
R53358 VCC.n11372 VCC.n11233 0.00853571
R53359 VCC.n11260 VCC.n11254 0.00853571
R53360 VCC.n11860 VCC.n11859 0.00853571
R53361 VCC.n11871 VCC.n11814 0.00853571
R53362 VCC.n11889 VCC.n11888 0.00853571
R53363 VCC.n11922 VCC.n11783 0.00853571
R53364 VCC.n11810 VCC.n11804 0.00853571
R53365 VCC.n11980 VCC.n11755 0.00853571
R53366 VCC.n11994 VCC.n11749 0.00853571
R53367 VCC.n12026 VCC.n11734 0.00853571
R53368 VCC.n12049 VCC.n11723 0.00853571
R53369 VCC.n12013 VCC.n12012 0.00853571
R53370 VCC.n12116 VCC.n11690 0.00853571
R53371 VCC.n12180 VCC.n12179 0.00853571
R53372 VCC.n12191 VCC.n11641 0.00853571
R53373 VCC.n12681 VCC.n12242 0.00853571
R53374 VCC.n12723 VCC.n12206 0.00853571
R53375 VCC.n12744 VCC.n12194 0.00853571
R53376 VCC.n12536 VCC.n12311 0.00853571
R53377 VCC.n12550 VCC.n12305 0.00853571
R53378 VCC.n12582 VCC.n12290 0.00853571
R53379 VCC.n12605 VCC.n12279 0.00853571
R53380 VCC.n12569 VCC.n12568 0.00853571
R53381 VCC.n12417 VCC.n12416 0.00853571
R53382 VCC.n12428 VCC.n12371 0.00853571
R53383 VCC.n12446 VCC.n12445 0.00853571
R53384 VCC.n12479 VCC.n12340 0.00853571
R53385 VCC.n12367 VCC.n12361 0.00853571
R53386 VCC.n12967 VCC.n12966 0.00853571
R53387 VCC.n12978 VCC.n12921 0.00853571
R53388 VCC.n12996 VCC.n12995 0.00853571
R53389 VCC.n13029 VCC.n12890 0.00853571
R53390 VCC.n12917 VCC.n12911 0.00853571
R53391 VCC.n13087 VCC.n12862 0.00853571
R53392 VCC.n13101 VCC.n12856 0.00853571
R53393 VCC.n13133 VCC.n12841 0.00853571
R53394 VCC.n13156 VCC.n12830 0.00853571
R53395 VCC.n13120 VCC.n13119 0.00853571
R53396 VCC.n13223 VCC.n12797 0.00853571
R53397 VCC.n13287 VCC.n13286 0.00853571
R53398 VCC.n13298 VCC.n12748 0.00853571
R53399 VCC.n13788 VCC.n13349 0.00853571
R53400 VCC.n13830 VCC.n13313 0.00853571
R53401 VCC.n13851 VCC.n13301 0.00853571
R53402 VCC.n13643 VCC.n13418 0.00853571
R53403 VCC.n13657 VCC.n13412 0.00853571
R53404 VCC.n13689 VCC.n13397 0.00853571
R53405 VCC.n13712 VCC.n13386 0.00853571
R53406 VCC.n13676 VCC.n13675 0.00853571
R53407 VCC.n13524 VCC.n13523 0.00853571
R53408 VCC.n13535 VCC.n13478 0.00853571
R53409 VCC.n13553 VCC.n13552 0.00853571
R53410 VCC.n13586 VCC.n13447 0.00853571
R53411 VCC.n13474 VCC.n13468 0.00853571
R53412 VCC.n14074 VCC.n14073 0.00853571
R53413 VCC.n14085 VCC.n14028 0.00853571
R53414 VCC.n14103 VCC.n14102 0.00853571
R53415 VCC.n14136 VCC.n13997 0.00853571
R53416 VCC.n14024 VCC.n14018 0.00853571
R53417 VCC.n14194 VCC.n13969 0.00853571
R53418 VCC.n14208 VCC.n13963 0.00853571
R53419 VCC.n14240 VCC.n13948 0.00853571
R53420 VCC.n14263 VCC.n13937 0.00853571
R53421 VCC.n14227 VCC.n14226 0.00853571
R53422 VCC.n14330 VCC.n13904 0.00853571
R53423 VCC.n14394 VCC.n14393 0.00853571
R53424 VCC.n14405 VCC.n13855 0.00853571
R53425 VCC.n14895 VCC.n14456 0.00853571
R53426 VCC.n14937 VCC.n14420 0.00853571
R53427 VCC.n14958 VCC.n14408 0.00853571
R53428 VCC.n14750 VCC.n14525 0.00853571
R53429 VCC.n14764 VCC.n14519 0.00853571
R53430 VCC.n14796 VCC.n14504 0.00853571
R53431 VCC.n14819 VCC.n14493 0.00853571
R53432 VCC.n14783 VCC.n14782 0.00853571
R53433 VCC.n14631 VCC.n14630 0.00853571
R53434 VCC.n14642 VCC.n14585 0.00853571
R53435 VCC.n14660 VCC.n14659 0.00853571
R53436 VCC.n14693 VCC.n14554 0.00853571
R53437 VCC.n14581 VCC.n14575 0.00853571
R53438 VCC.n15181 VCC.n15180 0.00853571
R53439 VCC.n15192 VCC.n15135 0.00853571
R53440 VCC.n15210 VCC.n15209 0.00853571
R53441 VCC.n15243 VCC.n15104 0.00853571
R53442 VCC.n15131 VCC.n15125 0.00853571
R53443 VCC.n15301 VCC.n15076 0.00853571
R53444 VCC.n15315 VCC.n15070 0.00853571
R53445 VCC.n15347 VCC.n15055 0.00853571
R53446 VCC.n15370 VCC.n15044 0.00853571
R53447 VCC.n15334 VCC.n15333 0.00853571
R53448 VCC.n15437 VCC.n15011 0.00853571
R53449 VCC.n15501 VCC.n15500 0.00853571
R53450 VCC.n15512 VCC.n14962 0.00853571
R53451 VCC.n16002 VCC.n15563 0.00853571
R53452 VCC.n16044 VCC.n15527 0.00853571
R53453 VCC.n16065 VCC.n15515 0.00853571
R53454 VCC.n15857 VCC.n15632 0.00853571
R53455 VCC.n15871 VCC.n15626 0.00853571
R53456 VCC.n15903 VCC.n15611 0.00853571
R53457 VCC.n15926 VCC.n15600 0.00853571
R53458 VCC.n15890 VCC.n15889 0.00853571
R53459 VCC.n15738 VCC.n15737 0.00853571
R53460 VCC.n15749 VCC.n15692 0.00853571
R53461 VCC.n15767 VCC.n15766 0.00853571
R53462 VCC.n15800 VCC.n15661 0.00853571
R53463 VCC.n15688 VCC.n15682 0.00853571
R53464 VCC.n16288 VCC.n16287 0.00853571
R53465 VCC.n16299 VCC.n16242 0.00853571
R53466 VCC.n16317 VCC.n16316 0.00853571
R53467 VCC.n16350 VCC.n16211 0.00853571
R53468 VCC.n16238 VCC.n16232 0.00853571
R53469 VCC.n16408 VCC.n16183 0.00853571
R53470 VCC.n16422 VCC.n16177 0.00853571
R53471 VCC.n16454 VCC.n16162 0.00853571
R53472 VCC.n16477 VCC.n16151 0.00853571
R53473 VCC.n16441 VCC.n16440 0.00853571
R53474 VCC.n16544 VCC.n16118 0.00853571
R53475 VCC.n16608 VCC.n16607 0.00853571
R53476 VCC.n16619 VCC.n16069 0.00853571
R53477 VCC.n17109 VCC.n16670 0.00853571
R53478 VCC.n17151 VCC.n16634 0.00853571
R53479 VCC.n17172 VCC.n16622 0.00853571
R53480 VCC.n16964 VCC.n16739 0.00853571
R53481 VCC.n16978 VCC.n16733 0.00853571
R53482 VCC.n17010 VCC.n16718 0.00853571
R53483 VCC.n17033 VCC.n16707 0.00853571
R53484 VCC.n16997 VCC.n16996 0.00853571
R53485 VCC.n16845 VCC.n16844 0.00853571
R53486 VCC.n16856 VCC.n16799 0.00853571
R53487 VCC.n16874 VCC.n16873 0.00853571
R53488 VCC.n16907 VCC.n16768 0.00853571
R53489 VCC.n16795 VCC.n16789 0.00853571
R53490 VCC.n17328 VCC.n17290 0.00853571
R53491 VCC.n17342 VCC.n17284 0.00853571
R53492 VCC.n17374 VCC.n17269 0.00853571
R53493 VCC.n17397 VCC.n17258 0.00853571
R53494 VCC.n17361 VCC.n17360 0.00853571
R53495 VCC.n17464 VCC.n17225 0.00853571
R53496 VCC.n17528 VCC.n17527 0.00853571
R53497 VCC.n17539 VCC.n17176 0.00853571
R53498 VCC.n191 VCC.n188 0.00822143
R53499 VCC.n241 VCC.n173 0.00822143
R53500 VCC.n281 VCC.n131 0.00822143
R53501 VCC.n313 VCC.n127 0.00822143
R53502 VCC.n316 VCC.n315 0.00822143
R53503 VCC.n347 VCC.n346 0.00822143
R53504 VCC.n408 VCC.n70 0.00822143
R53505 VCC.n448 VCC.n66 0.00822143
R53506 VCC.n449 VCC.n62 0.00822143
R53507 VCC.n481 VCC.n49 0.00822143
R53508 VCC.n513 VCC.n13 0.00822143
R53509 VCC.n552 VCC.n0 0.00822143
R53510 VCC.n743 VCC.n740 0.00822143
R53511 VCC.n793 VCC.n725 0.00822143
R53512 VCC.n833 VCC.n683 0.00822143
R53513 VCC.n865 VCC.n679 0.00822143
R53514 VCC.n868 VCC.n867 0.00822143
R53515 VCC.n899 VCC.n898 0.00822143
R53516 VCC.n960 VCC.n622 0.00822143
R53517 VCC.n1000 VCC.n618 0.00822143
R53518 VCC.n1001 VCC.n614 0.00822143
R53519 VCC.n1033 VCC.n601 0.00822143
R53520 VCC.n1065 VCC.n565 0.00822143
R53521 VCC.n1106 VCC.n554 0.00822143
R53522 VCC.n1301 VCC.n1298 0.00822143
R53523 VCC.n1351 VCC.n1283 0.00822143
R53524 VCC.n1391 VCC.n1241 0.00822143
R53525 VCC.n1423 VCC.n1237 0.00822143
R53526 VCC.n1426 VCC.n1425 0.00822143
R53527 VCC.n1456 VCC.n1455 0.00822143
R53528 VCC.n1517 VCC.n1179 0.00822143
R53529 VCC.n1558 VCC.n1175 0.00822143
R53530 VCC.n1559 VCC.n1171 0.00822143
R53531 VCC.n1599 VCC.n1154 0.00822143
R53532 VCC.n1629 VCC.n1126 0.00822143
R53533 VCC.n1660 VCC.n1108 0.00822143
R53534 VCC.n1852 VCC.n1849 0.00822143
R53535 VCC.n1902 VCC.n1834 0.00822143
R53536 VCC.n1942 VCC.n1792 0.00822143
R53537 VCC.n1974 VCC.n1788 0.00822143
R53538 VCC.n1977 VCC.n1976 0.00822143
R53539 VCC.n2008 VCC.n2007 0.00822143
R53540 VCC.n2069 VCC.n1731 0.00822143
R53541 VCC.n2109 VCC.n1727 0.00822143
R53542 VCC.n2110 VCC.n1723 0.00822143
R53543 VCC.n2142 VCC.n1710 0.00822143
R53544 VCC.n2174 VCC.n1674 0.00822143
R53545 VCC.n2215 VCC.n1663 0.00822143
R53546 VCC.n2410 VCC.n2407 0.00822143
R53547 VCC.n2460 VCC.n2392 0.00822143
R53548 VCC.n2500 VCC.n2350 0.00822143
R53549 VCC.n2532 VCC.n2346 0.00822143
R53550 VCC.n2535 VCC.n2534 0.00822143
R53551 VCC.n2565 VCC.n2564 0.00822143
R53552 VCC.n2626 VCC.n2288 0.00822143
R53553 VCC.n2667 VCC.n2284 0.00822143
R53554 VCC.n2668 VCC.n2280 0.00822143
R53555 VCC.n2708 VCC.n2263 0.00822143
R53556 VCC.n2738 VCC.n2235 0.00822143
R53557 VCC.n2769 VCC.n2217 0.00822143
R53558 VCC.n2961 VCC.n2958 0.00822143
R53559 VCC.n3011 VCC.n2943 0.00822143
R53560 VCC.n3051 VCC.n2901 0.00822143
R53561 VCC.n3083 VCC.n2897 0.00822143
R53562 VCC.n3086 VCC.n3085 0.00822143
R53563 VCC.n3117 VCC.n3116 0.00822143
R53564 VCC.n3178 VCC.n2840 0.00822143
R53565 VCC.n3218 VCC.n2836 0.00822143
R53566 VCC.n3219 VCC.n2832 0.00822143
R53567 VCC.n3251 VCC.n2819 0.00822143
R53568 VCC.n3283 VCC.n2783 0.00822143
R53569 VCC.n3324 VCC.n2772 0.00822143
R53570 VCC.n3519 VCC.n3516 0.00822143
R53571 VCC.n3569 VCC.n3501 0.00822143
R53572 VCC.n3609 VCC.n3459 0.00822143
R53573 VCC.n3641 VCC.n3455 0.00822143
R53574 VCC.n3644 VCC.n3643 0.00822143
R53575 VCC.n3674 VCC.n3673 0.00822143
R53576 VCC.n3735 VCC.n3397 0.00822143
R53577 VCC.n3776 VCC.n3393 0.00822143
R53578 VCC.n3777 VCC.n3389 0.00822143
R53579 VCC.n3817 VCC.n3372 0.00822143
R53580 VCC.n3847 VCC.n3344 0.00822143
R53581 VCC.n3878 VCC.n3326 0.00822143
R53582 VCC.n4070 VCC.n4067 0.00822143
R53583 VCC.n4120 VCC.n4052 0.00822143
R53584 VCC.n4160 VCC.n4010 0.00822143
R53585 VCC.n4192 VCC.n4006 0.00822143
R53586 VCC.n4195 VCC.n4194 0.00822143
R53587 VCC.n4226 VCC.n4225 0.00822143
R53588 VCC.n4287 VCC.n3949 0.00822143
R53589 VCC.n4327 VCC.n3945 0.00822143
R53590 VCC.n4328 VCC.n3941 0.00822143
R53591 VCC.n4360 VCC.n3928 0.00822143
R53592 VCC.n4392 VCC.n3892 0.00822143
R53593 VCC.n4433 VCC.n3881 0.00822143
R53594 VCC.n4628 VCC.n4625 0.00822143
R53595 VCC.n4678 VCC.n4610 0.00822143
R53596 VCC.n4718 VCC.n4568 0.00822143
R53597 VCC.n4750 VCC.n4564 0.00822143
R53598 VCC.n4753 VCC.n4752 0.00822143
R53599 VCC.n4783 VCC.n4782 0.00822143
R53600 VCC.n4844 VCC.n4506 0.00822143
R53601 VCC.n4885 VCC.n4502 0.00822143
R53602 VCC.n4886 VCC.n4498 0.00822143
R53603 VCC.n4926 VCC.n4481 0.00822143
R53604 VCC.n4956 VCC.n4453 0.00822143
R53605 VCC.n4987 VCC.n4435 0.00822143
R53606 VCC.n5179 VCC.n5176 0.00822143
R53607 VCC.n5229 VCC.n5161 0.00822143
R53608 VCC.n5269 VCC.n5119 0.00822143
R53609 VCC.n5301 VCC.n5115 0.00822143
R53610 VCC.n5304 VCC.n5303 0.00822143
R53611 VCC.n5335 VCC.n5334 0.00822143
R53612 VCC.n5396 VCC.n5058 0.00822143
R53613 VCC.n5436 VCC.n5054 0.00822143
R53614 VCC.n5437 VCC.n5050 0.00822143
R53615 VCC.n5469 VCC.n5037 0.00822143
R53616 VCC.n5501 VCC.n5001 0.00822143
R53617 VCC.n5542 VCC.n4990 0.00822143
R53618 VCC.n5737 VCC.n5734 0.00822143
R53619 VCC.n5787 VCC.n5719 0.00822143
R53620 VCC.n5827 VCC.n5677 0.00822143
R53621 VCC.n5859 VCC.n5673 0.00822143
R53622 VCC.n5862 VCC.n5861 0.00822143
R53623 VCC.n5892 VCC.n5891 0.00822143
R53624 VCC.n5953 VCC.n5615 0.00822143
R53625 VCC.n5994 VCC.n5611 0.00822143
R53626 VCC.n5995 VCC.n5607 0.00822143
R53627 VCC.n6035 VCC.n5590 0.00822143
R53628 VCC.n6065 VCC.n5562 0.00822143
R53629 VCC.n6096 VCC.n5544 0.00822143
R53630 VCC.n6288 VCC.n6285 0.00822143
R53631 VCC.n6338 VCC.n6270 0.00822143
R53632 VCC.n6378 VCC.n6228 0.00822143
R53633 VCC.n6410 VCC.n6224 0.00822143
R53634 VCC.n6413 VCC.n6412 0.00822143
R53635 VCC.n6444 VCC.n6443 0.00822143
R53636 VCC.n6505 VCC.n6167 0.00822143
R53637 VCC.n6545 VCC.n6163 0.00822143
R53638 VCC.n6546 VCC.n6159 0.00822143
R53639 VCC.n6578 VCC.n6146 0.00822143
R53640 VCC.n6610 VCC.n6110 0.00822143
R53641 VCC.n6651 VCC.n6099 0.00822143
R53642 VCC.n6846 VCC.n6843 0.00822143
R53643 VCC.n6896 VCC.n6828 0.00822143
R53644 VCC.n6936 VCC.n6786 0.00822143
R53645 VCC.n6968 VCC.n6782 0.00822143
R53646 VCC.n6971 VCC.n6970 0.00822143
R53647 VCC.n7001 VCC.n7000 0.00822143
R53648 VCC.n7062 VCC.n6724 0.00822143
R53649 VCC.n7103 VCC.n6720 0.00822143
R53650 VCC.n7104 VCC.n6716 0.00822143
R53651 VCC.n7144 VCC.n6699 0.00822143
R53652 VCC.n7174 VCC.n6671 0.00822143
R53653 VCC.n7205 VCC.n6653 0.00822143
R53654 VCC.n7397 VCC.n7394 0.00822143
R53655 VCC.n7447 VCC.n7379 0.00822143
R53656 VCC.n7487 VCC.n7337 0.00822143
R53657 VCC.n7519 VCC.n7333 0.00822143
R53658 VCC.n7522 VCC.n7521 0.00822143
R53659 VCC.n7553 VCC.n7552 0.00822143
R53660 VCC.n7614 VCC.n7276 0.00822143
R53661 VCC.n7654 VCC.n7272 0.00822143
R53662 VCC.n7655 VCC.n7268 0.00822143
R53663 VCC.n7687 VCC.n7255 0.00822143
R53664 VCC.n7719 VCC.n7219 0.00822143
R53665 VCC.n7760 VCC.n7208 0.00822143
R53666 VCC.n7955 VCC.n7952 0.00822143
R53667 VCC.n8005 VCC.n7937 0.00822143
R53668 VCC.n8045 VCC.n7895 0.00822143
R53669 VCC.n8077 VCC.n7891 0.00822143
R53670 VCC.n8080 VCC.n8079 0.00822143
R53671 VCC.n8110 VCC.n8109 0.00822143
R53672 VCC.n8171 VCC.n7833 0.00822143
R53673 VCC.n8212 VCC.n7829 0.00822143
R53674 VCC.n8213 VCC.n7825 0.00822143
R53675 VCC.n8253 VCC.n7808 0.00822143
R53676 VCC.n8283 VCC.n7780 0.00822143
R53677 VCC.n8314 VCC.n7762 0.00822143
R53678 VCC.n8631 VCC.n8630 0.00822143
R53679 VCC.n8662 VCC.n8661 0.00822143
R53680 VCC.n8723 VCC.n8385 0.00822143
R53681 VCC.n8763 VCC.n8381 0.00822143
R53682 VCC.n8764 VCC.n8377 0.00822143
R53683 VCC.n8796 VCC.n8364 0.00822143
R53684 VCC.n8828 VCC.n8328 0.00822143
R53685 VCC.n8869 VCC.n8317 0.00822143
R53686 VCC.n9064 VCC.n9061 0.00822143
R53687 VCC.n9114 VCC.n9046 0.00822143
R53688 VCC.n9154 VCC.n9004 0.00822143
R53689 VCC.n9186 VCC.n9000 0.00822143
R53690 VCC.n9189 VCC.n9188 0.00822143
R53691 VCC.n9219 VCC.n9218 0.00822143
R53692 VCC.n9280 VCC.n8942 0.00822143
R53693 VCC.n9321 VCC.n8938 0.00822143
R53694 VCC.n9322 VCC.n8934 0.00822143
R53695 VCC.n9362 VCC.n8917 0.00822143
R53696 VCC.n9392 VCC.n8889 0.00822143
R53697 VCC.n9423 VCC.n8871 0.00822143
R53698 VCC.n9615 VCC.n9612 0.00822143
R53699 VCC.n9665 VCC.n9597 0.00822143
R53700 VCC.n9705 VCC.n9555 0.00822143
R53701 VCC.n9737 VCC.n9551 0.00822143
R53702 VCC.n9740 VCC.n9739 0.00822143
R53703 VCC.n9771 VCC.n9770 0.00822143
R53704 VCC.n9832 VCC.n9494 0.00822143
R53705 VCC.n9872 VCC.n9490 0.00822143
R53706 VCC.n9873 VCC.n9486 0.00822143
R53707 VCC.n9905 VCC.n9473 0.00822143
R53708 VCC.n9937 VCC.n9437 0.00822143
R53709 VCC.n9978 VCC.n9426 0.00822143
R53710 VCC.n10172 VCC.n10169 0.00822143
R53711 VCC.n10222 VCC.n10154 0.00822143
R53712 VCC.n10262 VCC.n10112 0.00822143
R53713 VCC.n10294 VCC.n10108 0.00822143
R53714 VCC.n10297 VCC.n10296 0.00822143
R53715 VCC.n10327 VCC.n10326 0.00822143
R53716 VCC.n10388 VCC.n10050 0.00822143
R53717 VCC.n10429 VCC.n10046 0.00822143
R53718 VCC.n10430 VCC.n10042 0.00822143
R53719 VCC.n10470 VCC.n10025 0.00822143
R53720 VCC.n10500 VCC.n9997 0.00822143
R53721 VCC.n10531 VCC.n9979 0.00822143
R53722 VCC.n10722 VCC.n10719 0.00822143
R53723 VCC.n10772 VCC.n10704 0.00822143
R53724 VCC.n10812 VCC.n10662 0.00822143
R53725 VCC.n10844 VCC.n10658 0.00822143
R53726 VCC.n10847 VCC.n10846 0.00822143
R53727 VCC.n10878 VCC.n10877 0.00822143
R53728 VCC.n10939 VCC.n10601 0.00822143
R53729 VCC.n10979 VCC.n10597 0.00822143
R53730 VCC.n10980 VCC.n10593 0.00822143
R53731 VCC.n11012 VCC.n10580 0.00822143
R53732 VCC.n11044 VCC.n10544 0.00822143
R53733 VCC.n11085 VCC.n10533 0.00822143
R53734 VCC.n11279 VCC.n11276 0.00822143
R53735 VCC.n11329 VCC.n11261 0.00822143
R53736 VCC.n11369 VCC.n11219 0.00822143
R53737 VCC.n11401 VCC.n11215 0.00822143
R53738 VCC.n11404 VCC.n11403 0.00822143
R53739 VCC.n11434 VCC.n11433 0.00822143
R53740 VCC.n11495 VCC.n11157 0.00822143
R53741 VCC.n11536 VCC.n11153 0.00822143
R53742 VCC.n11537 VCC.n11149 0.00822143
R53743 VCC.n11577 VCC.n11132 0.00822143
R53744 VCC.n11607 VCC.n11104 0.00822143
R53745 VCC.n11638 VCC.n11086 0.00822143
R53746 VCC.n11829 VCC.n11826 0.00822143
R53747 VCC.n11879 VCC.n11811 0.00822143
R53748 VCC.n11919 VCC.n11769 0.00822143
R53749 VCC.n11951 VCC.n11765 0.00822143
R53750 VCC.n11954 VCC.n11953 0.00822143
R53751 VCC.n11985 VCC.n11984 0.00822143
R53752 VCC.n12046 VCC.n11708 0.00822143
R53753 VCC.n12086 VCC.n11704 0.00822143
R53754 VCC.n12087 VCC.n11700 0.00822143
R53755 VCC.n12119 VCC.n11687 0.00822143
R53756 VCC.n12151 VCC.n11651 0.00822143
R53757 VCC.n12192 VCC.n11640 0.00822143
R53758 VCC.n12386 VCC.n12383 0.00822143
R53759 VCC.n12436 VCC.n12368 0.00822143
R53760 VCC.n12476 VCC.n12326 0.00822143
R53761 VCC.n12508 VCC.n12322 0.00822143
R53762 VCC.n12511 VCC.n12510 0.00822143
R53763 VCC.n12541 VCC.n12540 0.00822143
R53764 VCC.n12602 VCC.n12264 0.00822143
R53765 VCC.n12643 VCC.n12260 0.00822143
R53766 VCC.n12644 VCC.n12256 0.00822143
R53767 VCC.n12684 VCC.n12239 0.00822143
R53768 VCC.n12714 VCC.n12211 0.00822143
R53769 VCC.n12745 VCC.n12193 0.00822143
R53770 VCC.n12936 VCC.n12933 0.00822143
R53771 VCC.n12986 VCC.n12918 0.00822143
R53772 VCC.n13026 VCC.n12876 0.00822143
R53773 VCC.n13058 VCC.n12872 0.00822143
R53774 VCC.n13061 VCC.n13060 0.00822143
R53775 VCC.n13092 VCC.n13091 0.00822143
R53776 VCC.n13153 VCC.n12815 0.00822143
R53777 VCC.n13193 VCC.n12811 0.00822143
R53778 VCC.n13194 VCC.n12807 0.00822143
R53779 VCC.n13226 VCC.n12794 0.00822143
R53780 VCC.n13258 VCC.n12758 0.00822143
R53781 VCC.n13299 VCC.n12747 0.00822143
R53782 VCC.n13493 VCC.n13490 0.00822143
R53783 VCC.n13543 VCC.n13475 0.00822143
R53784 VCC.n13583 VCC.n13433 0.00822143
R53785 VCC.n13615 VCC.n13429 0.00822143
R53786 VCC.n13618 VCC.n13617 0.00822143
R53787 VCC.n13648 VCC.n13647 0.00822143
R53788 VCC.n13709 VCC.n13371 0.00822143
R53789 VCC.n13750 VCC.n13367 0.00822143
R53790 VCC.n13751 VCC.n13363 0.00822143
R53791 VCC.n13791 VCC.n13346 0.00822143
R53792 VCC.n13821 VCC.n13318 0.00822143
R53793 VCC.n13852 VCC.n13300 0.00822143
R53794 VCC.n14043 VCC.n14040 0.00822143
R53795 VCC.n14093 VCC.n14025 0.00822143
R53796 VCC.n14133 VCC.n13983 0.00822143
R53797 VCC.n14165 VCC.n13979 0.00822143
R53798 VCC.n14168 VCC.n14167 0.00822143
R53799 VCC.n14199 VCC.n14198 0.00822143
R53800 VCC.n14260 VCC.n13922 0.00822143
R53801 VCC.n14300 VCC.n13918 0.00822143
R53802 VCC.n14301 VCC.n13914 0.00822143
R53803 VCC.n14333 VCC.n13901 0.00822143
R53804 VCC.n14365 VCC.n13865 0.00822143
R53805 VCC.n14406 VCC.n13854 0.00822143
R53806 VCC.n14600 VCC.n14597 0.00822143
R53807 VCC.n14650 VCC.n14582 0.00822143
R53808 VCC.n14690 VCC.n14540 0.00822143
R53809 VCC.n14722 VCC.n14536 0.00822143
R53810 VCC.n14725 VCC.n14724 0.00822143
R53811 VCC.n14755 VCC.n14754 0.00822143
R53812 VCC.n14816 VCC.n14478 0.00822143
R53813 VCC.n14857 VCC.n14474 0.00822143
R53814 VCC.n14858 VCC.n14470 0.00822143
R53815 VCC.n14898 VCC.n14453 0.00822143
R53816 VCC.n14928 VCC.n14425 0.00822143
R53817 VCC.n14959 VCC.n14407 0.00822143
R53818 VCC.n15150 VCC.n15147 0.00822143
R53819 VCC.n15200 VCC.n15132 0.00822143
R53820 VCC.n15240 VCC.n15090 0.00822143
R53821 VCC.n15272 VCC.n15086 0.00822143
R53822 VCC.n15275 VCC.n15274 0.00822143
R53823 VCC.n15306 VCC.n15305 0.00822143
R53824 VCC.n15367 VCC.n15029 0.00822143
R53825 VCC.n15407 VCC.n15025 0.00822143
R53826 VCC.n15408 VCC.n15021 0.00822143
R53827 VCC.n15440 VCC.n15008 0.00822143
R53828 VCC.n15472 VCC.n14972 0.00822143
R53829 VCC.n15513 VCC.n14961 0.00822143
R53830 VCC.n15707 VCC.n15704 0.00822143
R53831 VCC.n15757 VCC.n15689 0.00822143
R53832 VCC.n15797 VCC.n15647 0.00822143
R53833 VCC.n15829 VCC.n15643 0.00822143
R53834 VCC.n15832 VCC.n15831 0.00822143
R53835 VCC.n15862 VCC.n15861 0.00822143
R53836 VCC.n15923 VCC.n15585 0.00822143
R53837 VCC.n15964 VCC.n15581 0.00822143
R53838 VCC.n15965 VCC.n15577 0.00822143
R53839 VCC.n16005 VCC.n15560 0.00822143
R53840 VCC.n16035 VCC.n15532 0.00822143
R53841 VCC.n16066 VCC.n15514 0.00822143
R53842 VCC.n16257 VCC.n16254 0.00822143
R53843 VCC.n16307 VCC.n16239 0.00822143
R53844 VCC.n16347 VCC.n16197 0.00822143
R53845 VCC.n16379 VCC.n16193 0.00822143
R53846 VCC.n16382 VCC.n16381 0.00822143
R53847 VCC.n16413 VCC.n16412 0.00822143
R53848 VCC.n16474 VCC.n16136 0.00822143
R53849 VCC.n16514 VCC.n16132 0.00822143
R53850 VCC.n16515 VCC.n16128 0.00822143
R53851 VCC.n16547 VCC.n16115 0.00822143
R53852 VCC.n16579 VCC.n16079 0.00822143
R53853 VCC.n16620 VCC.n16068 0.00822143
R53854 VCC.n16814 VCC.n16811 0.00822143
R53855 VCC.n16864 VCC.n16796 0.00822143
R53856 VCC.n16904 VCC.n16754 0.00822143
R53857 VCC.n16936 VCC.n16750 0.00822143
R53858 VCC.n16939 VCC.n16938 0.00822143
R53859 VCC.n16969 VCC.n16968 0.00822143
R53860 VCC.n17030 VCC.n16692 0.00822143
R53861 VCC.n17071 VCC.n16688 0.00822143
R53862 VCC.n17072 VCC.n16684 0.00822143
R53863 VCC.n17112 VCC.n16667 0.00822143
R53864 VCC.n17142 VCC.n16639 0.00822143
R53865 VCC.n17173 VCC.n16621 0.00822143
R53866 VCC.n17302 VCC.n17301 0.00822143
R53867 VCC.n17333 VCC.n17332 0.00822143
R53868 VCC.n17394 VCC.n17243 0.00822143
R53869 VCC.n17434 VCC.n17239 0.00822143
R53870 VCC.n17435 VCC.n17235 0.00822143
R53871 VCC.n17467 VCC.n17222 0.00822143
R53872 VCC.n17499 VCC.n17186 0.00822143
R53873 VCC.n17540 VCC.n17175 0.00822143
R53874 VCC.n8506 VCC.n8503 0.00816667
R53875 VCC.n8556 VCC.n8488 0.00816667
R53876 VCC.n8596 VCC.n8446 0.00816667
R53877 VCC.n8628 VCC.n8442 0.00816667
R53878 VCC.n221 VCC.n176 0.00764286
R53879 VCC.n236 VCC.n235 0.00764286
R53880 VCC.n276 VCC.n274 0.00764286
R53881 VCC.n273 VCC.n145 0.00764286
R53882 VCC.n284 VCC.n134 0.00764286
R53883 VCC.n192 VCC.n189 0.00764286
R53884 VCC.n234 VCC.n175 0.00764286
R53885 VCC.n244 VCC.n172 0.00764286
R53886 VCC.n260 VCC.n164 0.00764286
R53887 VCC.n279 VCC.n148 0.00764286
R53888 VCC.n275 VCC.n146 0.00764286
R53889 VCC.n117 VCC.n111 0.00764286
R53890 VCC.n404 VCC.n403 0.00764286
R53891 VCC.n400 VCC.n85 0.00764286
R53892 VCC.n411 VCC.n73 0.00764286
R53893 VCC.n354 VCC.n353 0.00764286
R53894 VCC.n368 VCC.n103 0.00764286
R53895 VCC.n369 VCC.n100 0.00764286
R53896 VCC.n374 VCC.n373 0.00764286
R53897 VCC.n402 VCC.n89 0.00764286
R53898 VCC.n447 VCC.n67 0.00764286
R53899 VCC.n477 VCC.n53 0.00764286
R53900 VCC.n516 VCC.n27 0.00764286
R53901 VCC.n450 VCC.n63 0.00764286
R53902 VCC.n480 VCC.n479 0.00764286
R53903 VCC.n487 VCC.n46 0.00764286
R53904 VCC.n483 VCC.n482 0.00764286
R53905 VCC.n506 VCC.n34 0.00764286
R53906 VCC.n520 VCC.n28 0.00764286
R53907 VCC.n773 VCC.n728 0.00764286
R53908 VCC.n788 VCC.n787 0.00764286
R53909 VCC.n828 VCC.n826 0.00764286
R53910 VCC.n825 VCC.n697 0.00764286
R53911 VCC.n836 VCC.n686 0.00764286
R53912 VCC.n744 VCC.n741 0.00764286
R53913 VCC.n786 VCC.n727 0.00764286
R53914 VCC.n796 VCC.n724 0.00764286
R53915 VCC.n812 VCC.n716 0.00764286
R53916 VCC.n831 VCC.n700 0.00764286
R53917 VCC.n827 VCC.n698 0.00764286
R53918 VCC.n669 VCC.n663 0.00764286
R53919 VCC.n956 VCC.n955 0.00764286
R53920 VCC.n952 VCC.n637 0.00764286
R53921 VCC.n963 VCC.n625 0.00764286
R53922 VCC.n906 VCC.n905 0.00764286
R53923 VCC.n920 VCC.n655 0.00764286
R53924 VCC.n921 VCC.n652 0.00764286
R53925 VCC.n926 VCC.n925 0.00764286
R53926 VCC.n954 VCC.n641 0.00764286
R53927 VCC.n999 VCC.n619 0.00764286
R53928 VCC.n1029 VCC.n605 0.00764286
R53929 VCC.n1068 VCC.n579 0.00764286
R53930 VCC.n1002 VCC.n615 0.00764286
R53931 VCC.n1032 VCC.n1031 0.00764286
R53932 VCC.n1039 VCC.n598 0.00764286
R53933 VCC.n1035 VCC.n1034 0.00764286
R53934 VCC.n1058 VCC.n586 0.00764286
R53935 VCC.n1072 VCC.n580 0.00764286
R53936 VCC.n1595 VCC.n1158 0.00764286
R53937 VCC.n1139 VCC.n1138 0.00764286
R53938 VCC.n1560 VCC.n1172 0.00764286
R53939 VCC.n1598 VCC.n1597 0.00764286
R53940 VCC.n1591 VCC.n1590 0.00764286
R53941 VCC.n1602 VCC.n1151 0.00764286
R53942 VCC.n1610 VCC.n1609 0.00764286
R53943 VCC.n1136 VCC.n1132 0.00764286
R53944 VCC.n1226 VCC.n1220 0.00764286
R53945 VCC.n1513 VCC.n1512 0.00764286
R53946 VCC.n1509 VCC.n1194 0.00764286
R53947 VCC.n1520 VCC.n1182 0.00764286
R53948 VCC.n1463 VCC.n1462 0.00764286
R53949 VCC.n1477 VCC.n1212 0.00764286
R53950 VCC.n1478 VCC.n1209 0.00764286
R53951 VCC.n1483 VCC.n1482 0.00764286
R53952 VCC.n1511 VCC.n1198 0.00764286
R53953 VCC.n1557 VCC.n1176 0.00764286
R53954 VCC.n1331 VCC.n1286 0.00764286
R53955 VCC.n1346 VCC.n1345 0.00764286
R53956 VCC.n1386 VCC.n1384 0.00764286
R53957 VCC.n1383 VCC.n1255 0.00764286
R53958 VCC.n1394 VCC.n1244 0.00764286
R53959 VCC.n1302 VCC.n1299 0.00764286
R53960 VCC.n1344 VCC.n1285 0.00764286
R53961 VCC.n1354 VCC.n1282 0.00764286
R53962 VCC.n1370 VCC.n1274 0.00764286
R53963 VCC.n1389 VCC.n1258 0.00764286
R53964 VCC.n1385 VCC.n1256 0.00764286
R53965 VCC.n1882 VCC.n1837 0.00764286
R53966 VCC.n1897 VCC.n1896 0.00764286
R53967 VCC.n1937 VCC.n1935 0.00764286
R53968 VCC.n1934 VCC.n1806 0.00764286
R53969 VCC.n1945 VCC.n1795 0.00764286
R53970 VCC.n1853 VCC.n1850 0.00764286
R53971 VCC.n1895 VCC.n1836 0.00764286
R53972 VCC.n1905 VCC.n1833 0.00764286
R53973 VCC.n1921 VCC.n1825 0.00764286
R53974 VCC.n1940 VCC.n1809 0.00764286
R53975 VCC.n1936 VCC.n1807 0.00764286
R53976 VCC.n1778 VCC.n1772 0.00764286
R53977 VCC.n2065 VCC.n2064 0.00764286
R53978 VCC.n2061 VCC.n1746 0.00764286
R53979 VCC.n2072 VCC.n1734 0.00764286
R53980 VCC.n2015 VCC.n2014 0.00764286
R53981 VCC.n2029 VCC.n1764 0.00764286
R53982 VCC.n2030 VCC.n1761 0.00764286
R53983 VCC.n2035 VCC.n2034 0.00764286
R53984 VCC.n2063 VCC.n1750 0.00764286
R53985 VCC.n2108 VCC.n1728 0.00764286
R53986 VCC.n2138 VCC.n1714 0.00764286
R53987 VCC.n2177 VCC.n1688 0.00764286
R53988 VCC.n2111 VCC.n1724 0.00764286
R53989 VCC.n2141 VCC.n2140 0.00764286
R53990 VCC.n2148 VCC.n1707 0.00764286
R53991 VCC.n2144 VCC.n2143 0.00764286
R53992 VCC.n2167 VCC.n1695 0.00764286
R53993 VCC.n2181 VCC.n1689 0.00764286
R53994 VCC.n2704 VCC.n2267 0.00764286
R53995 VCC.n2248 VCC.n2247 0.00764286
R53996 VCC.n2669 VCC.n2281 0.00764286
R53997 VCC.n2707 VCC.n2706 0.00764286
R53998 VCC.n2700 VCC.n2699 0.00764286
R53999 VCC.n2711 VCC.n2260 0.00764286
R54000 VCC.n2719 VCC.n2718 0.00764286
R54001 VCC.n2245 VCC.n2241 0.00764286
R54002 VCC.n2335 VCC.n2329 0.00764286
R54003 VCC.n2622 VCC.n2621 0.00764286
R54004 VCC.n2618 VCC.n2303 0.00764286
R54005 VCC.n2629 VCC.n2291 0.00764286
R54006 VCC.n2572 VCC.n2571 0.00764286
R54007 VCC.n2586 VCC.n2321 0.00764286
R54008 VCC.n2587 VCC.n2318 0.00764286
R54009 VCC.n2592 VCC.n2591 0.00764286
R54010 VCC.n2620 VCC.n2307 0.00764286
R54011 VCC.n2666 VCC.n2285 0.00764286
R54012 VCC.n2440 VCC.n2395 0.00764286
R54013 VCC.n2455 VCC.n2454 0.00764286
R54014 VCC.n2495 VCC.n2493 0.00764286
R54015 VCC.n2492 VCC.n2364 0.00764286
R54016 VCC.n2503 VCC.n2353 0.00764286
R54017 VCC.n2411 VCC.n2408 0.00764286
R54018 VCC.n2453 VCC.n2394 0.00764286
R54019 VCC.n2463 VCC.n2391 0.00764286
R54020 VCC.n2479 VCC.n2383 0.00764286
R54021 VCC.n2498 VCC.n2367 0.00764286
R54022 VCC.n2494 VCC.n2365 0.00764286
R54023 VCC.n2991 VCC.n2946 0.00764286
R54024 VCC.n3006 VCC.n3005 0.00764286
R54025 VCC.n3046 VCC.n3044 0.00764286
R54026 VCC.n3043 VCC.n2915 0.00764286
R54027 VCC.n3054 VCC.n2904 0.00764286
R54028 VCC.n2962 VCC.n2959 0.00764286
R54029 VCC.n3004 VCC.n2945 0.00764286
R54030 VCC.n3014 VCC.n2942 0.00764286
R54031 VCC.n3030 VCC.n2934 0.00764286
R54032 VCC.n3049 VCC.n2918 0.00764286
R54033 VCC.n3045 VCC.n2916 0.00764286
R54034 VCC.n2887 VCC.n2881 0.00764286
R54035 VCC.n3174 VCC.n3173 0.00764286
R54036 VCC.n3170 VCC.n2855 0.00764286
R54037 VCC.n3181 VCC.n2843 0.00764286
R54038 VCC.n3124 VCC.n3123 0.00764286
R54039 VCC.n3138 VCC.n2873 0.00764286
R54040 VCC.n3139 VCC.n2870 0.00764286
R54041 VCC.n3144 VCC.n3143 0.00764286
R54042 VCC.n3172 VCC.n2859 0.00764286
R54043 VCC.n3217 VCC.n2837 0.00764286
R54044 VCC.n3247 VCC.n2823 0.00764286
R54045 VCC.n3286 VCC.n2797 0.00764286
R54046 VCC.n3220 VCC.n2833 0.00764286
R54047 VCC.n3250 VCC.n3249 0.00764286
R54048 VCC.n3257 VCC.n2816 0.00764286
R54049 VCC.n3253 VCC.n3252 0.00764286
R54050 VCC.n3276 VCC.n2804 0.00764286
R54051 VCC.n3290 VCC.n2798 0.00764286
R54052 VCC.n3813 VCC.n3376 0.00764286
R54053 VCC.n3357 VCC.n3356 0.00764286
R54054 VCC.n3778 VCC.n3390 0.00764286
R54055 VCC.n3816 VCC.n3815 0.00764286
R54056 VCC.n3809 VCC.n3808 0.00764286
R54057 VCC.n3820 VCC.n3369 0.00764286
R54058 VCC.n3828 VCC.n3827 0.00764286
R54059 VCC.n3354 VCC.n3350 0.00764286
R54060 VCC.n3444 VCC.n3438 0.00764286
R54061 VCC.n3731 VCC.n3730 0.00764286
R54062 VCC.n3727 VCC.n3412 0.00764286
R54063 VCC.n3738 VCC.n3400 0.00764286
R54064 VCC.n3681 VCC.n3680 0.00764286
R54065 VCC.n3695 VCC.n3430 0.00764286
R54066 VCC.n3696 VCC.n3427 0.00764286
R54067 VCC.n3701 VCC.n3700 0.00764286
R54068 VCC.n3729 VCC.n3416 0.00764286
R54069 VCC.n3775 VCC.n3394 0.00764286
R54070 VCC.n3549 VCC.n3504 0.00764286
R54071 VCC.n3564 VCC.n3563 0.00764286
R54072 VCC.n3604 VCC.n3602 0.00764286
R54073 VCC.n3601 VCC.n3473 0.00764286
R54074 VCC.n3612 VCC.n3462 0.00764286
R54075 VCC.n3520 VCC.n3517 0.00764286
R54076 VCC.n3562 VCC.n3503 0.00764286
R54077 VCC.n3572 VCC.n3500 0.00764286
R54078 VCC.n3588 VCC.n3492 0.00764286
R54079 VCC.n3607 VCC.n3476 0.00764286
R54080 VCC.n3603 VCC.n3474 0.00764286
R54081 VCC.n4100 VCC.n4055 0.00764286
R54082 VCC.n4115 VCC.n4114 0.00764286
R54083 VCC.n4155 VCC.n4153 0.00764286
R54084 VCC.n4152 VCC.n4024 0.00764286
R54085 VCC.n4163 VCC.n4013 0.00764286
R54086 VCC.n4071 VCC.n4068 0.00764286
R54087 VCC.n4113 VCC.n4054 0.00764286
R54088 VCC.n4123 VCC.n4051 0.00764286
R54089 VCC.n4139 VCC.n4043 0.00764286
R54090 VCC.n4158 VCC.n4027 0.00764286
R54091 VCC.n4154 VCC.n4025 0.00764286
R54092 VCC.n3996 VCC.n3990 0.00764286
R54093 VCC.n4283 VCC.n4282 0.00764286
R54094 VCC.n4279 VCC.n3964 0.00764286
R54095 VCC.n4290 VCC.n3952 0.00764286
R54096 VCC.n4233 VCC.n4232 0.00764286
R54097 VCC.n4247 VCC.n3982 0.00764286
R54098 VCC.n4248 VCC.n3979 0.00764286
R54099 VCC.n4253 VCC.n4252 0.00764286
R54100 VCC.n4281 VCC.n3968 0.00764286
R54101 VCC.n4326 VCC.n3946 0.00764286
R54102 VCC.n4356 VCC.n3932 0.00764286
R54103 VCC.n4395 VCC.n3906 0.00764286
R54104 VCC.n4329 VCC.n3942 0.00764286
R54105 VCC.n4359 VCC.n4358 0.00764286
R54106 VCC.n4366 VCC.n3925 0.00764286
R54107 VCC.n4362 VCC.n4361 0.00764286
R54108 VCC.n4385 VCC.n3913 0.00764286
R54109 VCC.n4399 VCC.n3907 0.00764286
R54110 VCC.n4922 VCC.n4485 0.00764286
R54111 VCC.n4466 VCC.n4465 0.00764286
R54112 VCC.n4887 VCC.n4499 0.00764286
R54113 VCC.n4925 VCC.n4924 0.00764286
R54114 VCC.n4918 VCC.n4917 0.00764286
R54115 VCC.n4929 VCC.n4478 0.00764286
R54116 VCC.n4937 VCC.n4936 0.00764286
R54117 VCC.n4463 VCC.n4459 0.00764286
R54118 VCC.n4553 VCC.n4547 0.00764286
R54119 VCC.n4840 VCC.n4839 0.00764286
R54120 VCC.n4836 VCC.n4521 0.00764286
R54121 VCC.n4847 VCC.n4509 0.00764286
R54122 VCC.n4790 VCC.n4789 0.00764286
R54123 VCC.n4804 VCC.n4539 0.00764286
R54124 VCC.n4805 VCC.n4536 0.00764286
R54125 VCC.n4810 VCC.n4809 0.00764286
R54126 VCC.n4838 VCC.n4525 0.00764286
R54127 VCC.n4884 VCC.n4503 0.00764286
R54128 VCC.n4658 VCC.n4613 0.00764286
R54129 VCC.n4673 VCC.n4672 0.00764286
R54130 VCC.n4713 VCC.n4711 0.00764286
R54131 VCC.n4710 VCC.n4582 0.00764286
R54132 VCC.n4721 VCC.n4571 0.00764286
R54133 VCC.n4629 VCC.n4626 0.00764286
R54134 VCC.n4671 VCC.n4612 0.00764286
R54135 VCC.n4681 VCC.n4609 0.00764286
R54136 VCC.n4697 VCC.n4601 0.00764286
R54137 VCC.n4716 VCC.n4585 0.00764286
R54138 VCC.n4712 VCC.n4583 0.00764286
R54139 VCC.n5209 VCC.n5164 0.00764286
R54140 VCC.n5224 VCC.n5223 0.00764286
R54141 VCC.n5264 VCC.n5262 0.00764286
R54142 VCC.n5261 VCC.n5133 0.00764286
R54143 VCC.n5272 VCC.n5122 0.00764286
R54144 VCC.n5180 VCC.n5177 0.00764286
R54145 VCC.n5222 VCC.n5163 0.00764286
R54146 VCC.n5232 VCC.n5160 0.00764286
R54147 VCC.n5248 VCC.n5152 0.00764286
R54148 VCC.n5267 VCC.n5136 0.00764286
R54149 VCC.n5263 VCC.n5134 0.00764286
R54150 VCC.n5105 VCC.n5099 0.00764286
R54151 VCC.n5392 VCC.n5391 0.00764286
R54152 VCC.n5388 VCC.n5073 0.00764286
R54153 VCC.n5399 VCC.n5061 0.00764286
R54154 VCC.n5342 VCC.n5341 0.00764286
R54155 VCC.n5356 VCC.n5091 0.00764286
R54156 VCC.n5357 VCC.n5088 0.00764286
R54157 VCC.n5362 VCC.n5361 0.00764286
R54158 VCC.n5390 VCC.n5077 0.00764286
R54159 VCC.n5435 VCC.n5055 0.00764286
R54160 VCC.n5465 VCC.n5041 0.00764286
R54161 VCC.n5504 VCC.n5015 0.00764286
R54162 VCC.n5438 VCC.n5051 0.00764286
R54163 VCC.n5468 VCC.n5467 0.00764286
R54164 VCC.n5475 VCC.n5034 0.00764286
R54165 VCC.n5471 VCC.n5470 0.00764286
R54166 VCC.n5494 VCC.n5022 0.00764286
R54167 VCC.n5508 VCC.n5016 0.00764286
R54168 VCC.n6031 VCC.n5594 0.00764286
R54169 VCC.n5575 VCC.n5574 0.00764286
R54170 VCC.n5996 VCC.n5608 0.00764286
R54171 VCC.n6034 VCC.n6033 0.00764286
R54172 VCC.n6027 VCC.n6026 0.00764286
R54173 VCC.n6038 VCC.n5587 0.00764286
R54174 VCC.n6046 VCC.n6045 0.00764286
R54175 VCC.n5572 VCC.n5568 0.00764286
R54176 VCC.n5662 VCC.n5656 0.00764286
R54177 VCC.n5949 VCC.n5948 0.00764286
R54178 VCC.n5945 VCC.n5630 0.00764286
R54179 VCC.n5956 VCC.n5618 0.00764286
R54180 VCC.n5899 VCC.n5898 0.00764286
R54181 VCC.n5913 VCC.n5648 0.00764286
R54182 VCC.n5914 VCC.n5645 0.00764286
R54183 VCC.n5919 VCC.n5918 0.00764286
R54184 VCC.n5947 VCC.n5634 0.00764286
R54185 VCC.n5993 VCC.n5612 0.00764286
R54186 VCC.n5767 VCC.n5722 0.00764286
R54187 VCC.n5782 VCC.n5781 0.00764286
R54188 VCC.n5822 VCC.n5820 0.00764286
R54189 VCC.n5819 VCC.n5691 0.00764286
R54190 VCC.n5830 VCC.n5680 0.00764286
R54191 VCC.n5738 VCC.n5735 0.00764286
R54192 VCC.n5780 VCC.n5721 0.00764286
R54193 VCC.n5790 VCC.n5718 0.00764286
R54194 VCC.n5806 VCC.n5710 0.00764286
R54195 VCC.n5825 VCC.n5694 0.00764286
R54196 VCC.n5821 VCC.n5692 0.00764286
R54197 VCC.n6318 VCC.n6273 0.00764286
R54198 VCC.n6333 VCC.n6332 0.00764286
R54199 VCC.n6373 VCC.n6371 0.00764286
R54200 VCC.n6370 VCC.n6242 0.00764286
R54201 VCC.n6381 VCC.n6231 0.00764286
R54202 VCC.n6289 VCC.n6286 0.00764286
R54203 VCC.n6331 VCC.n6272 0.00764286
R54204 VCC.n6341 VCC.n6269 0.00764286
R54205 VCC.n6357 VCC.n6261 0.00764286
R54206 VCC.n6376 VCC.n6245 0.00764286
R54207 VCC.n6372 VCC.n6243 0.00764286
R54208 VCC.n6214 VCC.n6208 0.00764286
R54209 VCC.n6501 VCC.n6500 0.00764286
R54210 VCC.n6497 VCC.n6182 0.00764286
R54211 VCC.n6508 VCC.n6170 0.00764286
R54212 VCC.n6451 VCC.n6450 0.00764286
R54213 VCC.n6465 VCC.n6200 0.00764286
R54214 VCC.n6466 VCC.n6197 0.00764286
R54215 VCC.n6471 VCC.n6470 0.00764286
R54216 VCC.n6499 VCC.n6186 0.00764286
R54217 VCC.n6544 VCC.n6164 0.00764286
R54218 VCC.n6574 VCC.n6150 0.00764286
R54219 VCC.n6613 VCC.n6124 0.00764286
R54220 VCC.n6547 VCC.n6160 0.00764286
R54221 VCC.n6577 VCC.n6576 0.00764286
R54222 VCC.n6584 VCC.n6143 0.00764286
R54223 VCC.n6580 VCC.n6579 0.00764286
R54224 VCC.n6603 VCC.n6131 0.00764286
R54225 VCC.n6617 VCC.n6125 0.00764286
R54226 VCC.n7140 VCC.n6703 0.00764286
R54227 VCC.n6684 VCC.n6683 0.00764286
R54228 VCC.n7105 VCC.n6717 0.00764286
R54229 VCC.n7143 VCC.n7142 0.00764286
R54230 VCC.n7136 VCC.n7135 0.00764286
R54231 VCC.n7147 VCC.n6696 0.00764286
R54232 VCC.n7155 VCC.n7154 0.00764286
R54233 VCC.n6681 VCC.n6677 0.00764286
R54234 VCC.n6771 VCC.n6765 0.00764286
R54235 VCC.n7058 VCC.n7057 0.00764286
R54236 VCC.n7054 VCC.n6739 0.00764286
R54237 VCC.n7065 VCC.n6727 0.00764286
R54238 VCC.n7008 VCC.n7007 0.00764286
R54239 VCC.n7022 VCC.n6757 0.00764286
R54240 VCC.n7023 VCC.n6754 0.00764286
R54241 VCC.n7028 VCC.n7027 0.00764286
R54242 VCC.n7056 VCC.n6743 0.00764286
R54243 VCC.n7102 VCC.n6721 0.00764286
R54244 VCC.n6876 VCC.n6831 0.00764286
R54245 VCC.n6891 VCC.n6890 0.00764286
R54246 VCC.n6931 VCC.n6929 0.00764286
R54247 VCC.n6928 VCC.n6800 0.00764286
R54248 VCC.n6939 VCC.n6789 0.00764286
R54249 VCC.n6847 VCC.n6844 0.00764286
R54250 VCC.n6889 VCC.n6830 0.00764286
R54251 VCC.n6899 VCC.n6827 0.00764286
R54252 VCC.n6915 VCC.n6819 0.00764286
R54253 VCC.n6934 VCC.n6803 0.00764286
R54254 VCC.n6930 VCC.n6801 0.00764286
R54255 VCC.n7427 VCC.n7382 0.00764286
R54256 VCC.n7442 VCC.n7441 0.00764286
R54257 VCC.n7482 VCC.n7480 0.00764286
R54258 VCC.n7479 VCC.n7351 0.00764286
R54259 VCC.n7490 VCC.n7340 0.00764286
R54260 VCC.n7398 VCC.n7395 0.00764286
R54261 VCC.n7440 VCC.n7381 0.00764286
R54262 VCC.n7450 VCC.n7378 0.00764286
R54263 VCC.n7466 VCC.n7370 0.00764286
R54264 VCC.n7485 VCC.n7354 0.00764286
R54265 VCC.n7481 VCC.n7352 0.00764286
R54266 VCC.n7323 VCC.n7317 0.00764286
R54267 VCC.n7610 VCC.n7609 0.00764286
R54268 VCC.n7606 VCC.n7291 0.00764286
R54269 VCC.n7617 VCC.n7279 0.00764286
R54270 VCC.n7560 VCC.n7559 0.00764286
R54271 VCC.n7574 VCC.n7309 0.00764286
R54272 VCC.n7575 VCC.n7306 0.00764286
R54273 VCC.n7580 VCC.n7579 0.00764286
R54274 VCC.n7608 VCC.n7295 0.00764286
R54275 VCC.n7653 VCC.n7273 0.00764286
R54276 VCC.n7683 VCC.n7259 0.00764286
R54277 VCC.n7722 VCC.n7233 0.00764286
R54278 VCC.n7656 VCC.n7269 0.00764286
R54279 VCC.n7686 VCC.n7685 0.00764286
R54280 VCC.n7693 VCC.n7252 0.00764286
R54281 VCC.n7689 VCC.n7688 0.00764286
R54282 VCC.n7712 VCC.n7240 0.00764286
R54283 VCC.n7726 VCC.n7234 0.00764286
R54284 VCC.n8249 VCC.n7812 0.00764286
R54285 VCC.n7793 VCC.n7792 0.00764286
R54286 VCC.n8214 VCC.n7826 0.00764286
R54287 VCC.n8252 VCC.n8251 0.00764286
R54288 VCC.n8245 VCC.n8244 0.00764286
R54289 VCC.n8256 VCC.n7805 0.00764286
R54290 VCC.n8264 VCC.n8263 0.00764286
R54291 VCC.n7790 VCC.n7786 0.00764286
R54292 VCC.n7880 VCC.n7874 0.00764286
R54293 VCC.n8167 VCC.n8166 0.00764286
R54294 VCC.n8163 VCC.n7848 0.00764286
R54295 VCC.n8174 VCC.n7836 0.00764286
R54296 VCC.n8117 VCC.n8116 0.00764286
R54297 VCC.n8131 VCC.n7866 0.00764286
R54298 VCC.n8132 VCC.n7863 0.00764286
R54299 VCC.n8137 VCC.n8136 0.00764286
R54300 VCC.n8165 VCC.n7852 0.00764286
R54301 VCC.n8211 VCC.n7830 0.00764286
R54302 VCC.n7985 VCC.n7940 0.00764286
R54303 VCC.n8000 VCC.n7999 0.00764286
R54304 VCC.n8040 VCC.n8038 0.00764286
R54305 VCC.n8037 VCC.n7909 0.00764286
R54306 VCC.n8048 VCC.n7898 0.00764286
R54307 VCC.n7956 VCC.n7953 0.00764286
R54308 VCC.n7998 VCC.n7939 0.00764286
R54309 VCC.n8008 VCC.n7936 0.00764286
R54310 VCC.n8024 VCC.n7928 0.00764286
R54311 VCC.n8043 VCC.n7912 0.00764286
R54312 VCC.n8039 VCC.n7910 0.00764286
R54313 VCC.n8432 VCC.n8426 0.00764286
R54314 VCC.n8719 VCC.n8718 0.00764286
R54315 VCC.n8715 VCC.n8400 0.00764286
R54316 VCC.n8726 VCC.n8388 0.00764286
R54317 VCC.n8669 VCC.n8668 0.00764286
R54318 VCC.n8683 VCC.n8418 0.00764286
R54319 VCC.n8684 VCC.n8415 0.00764286
R54320 VCC.n8689 VCC.n8688 0.00764286
R54321 VCC.n8717 VCC.n8404 0.00764286
R54322 VCC.n8762 VCC.n8382 0.00764286
R54323 VCC.n8792 VCC.n8368 0.00764286
R54324 VCC.n8831 VCC.n8342 0.00764286
R54325 VCC.n8765 VCC.n8378 0.00764286
R54326 VCC.n8795 VCC.n8794 0.00764286
R54327 VCC.n8802 VCC.n8361 0.00764286
R54328 VCC.n8798 VCC.n8797 0.00764286
R54329 VCC.n8821 VCC.n8349 0.00764286
R54330 VCC.n8835 VCC.n8343 0.00764286
R54331 VCC.n8536 VCC.n8491 0.00764286
R54332 VCC.n8551 VCC.n8550 0.00764286
R54333 VCC.n8591 VCC.n8589 0.00764286
R54334 VCC.n8588 VCC.n8460 0.00764286
R54335 VCC.n8599 VCC.n8449 0.00764286
R54336 VCC.n8507 VCC.n8504 0.00764286
R54337 VCC.n8549 VCC.n8490 0.00764286
R54338 VCC.n8559 VCC.n8487 0.00764286
R54339 VCC.n8575 VCC.n8479 0.00764286
R54340 VCC.n8594 VCC.n8463 0.00764286
R54341 VCC.n8590 VCC.n8461 0.00764286
R54342 VCC.n9358 VCC.n8921 0.00764286
R54343 VCC.n8902 VCC.n8901 0.00764286
R54344 VCC.n9323 VCC.n8935 0.00764286
R54345 VCC.n9361 VCC.n9360 0.00764286
R54346 VCC.n9354 VCC.n9353 0.00764286
R54347 VCC.n9365 VCC.n8914 0.00764286
R54348 VCC.n9373 VCC.n9372 0.00764286
R54349 VCC.n8899 VCC.n8895 0.00764286
R54350 VCC.n8989 VCC.n8983 0.00764286
R54351 VCC.n9276 VCC.n9275 0.00764286
R54352 VCC.n9272 VCC.n8957 0.00764286
R54353 VCC.n9283 VCC.n8945 0.00764286
R54354 VCC.n9226 VCC.n9225 0.00764286
R54355 VCC.n9240 VCC.n8975 0.00764286
R54356 VCC.n9241 VCC.n8972 0.00764286
R54357 VCC.n9246 VCC.n9245 0.00764286
R54358 VCC.n9274 VCC.n8961 0.00764286
R54359 VCC.n9320 VCC.n8939 0.00764286
R54360 VCC.n9094 VCC.n9049 0.00764286
R54361 VCC.n9109 VCC.n9108 0.00764286
R54362 VCC.n9149 VCC.n9147 0.00764286
R54363 VCC.n9146 VCC.n9018 0.00764286
R54364 VCC.n9157 VCC.n9007 0.00764286
R54365 VCC.n9065 VCC.n9062 0.00764286
R54366 VCC.n9107 VCC.n9048 0.00764286
R54367 VCC.n9117 VCC.n9045 0.00764286
R54368 VCC.n9133 VCC.n9037 0.00764286
R54369 VCC.n9152 VCC.n9021 0.00764286
R54370 VCC.n9148 VCC.n9019 0.00764286
R54371 VCC.n9645 VCC.n9600 0.00764286
R54372 VCC.n9660 VCC.n9659 0.00764286
R54373 VCC.n9700 VCC.n9698 0.00764286
R54374 VCC.n9697 VCC.n9569 0.00764286
R54375 VCC.n9708 VCC.n9558 0.00764286
R54376 VCC.n9616 VCC.n9613 0.00764286
R54377 VCC.n9658 VCC.n9599 0.00764286
R54378 VCC.n9668 VCC.n9596 0.00764286
R54379 VCC.n9684 VCC.n9588 0.00764286
R54380 VCC.n9703 VCC.n9572 0.00764286
R54381 VCC.n9699 VCC.n9570 0.00764286
R54382 VCC.n9541 VCC.n9535 0.00764286
R54383 VCC.n9828 VCC.n9827 0.00764286
R54384 VCC.n9824 VCC.n9509 0.00764286
R54385 VCC.n9835 VCC.n9497 0.00764286
R54386 VCC.n9778 VCC.n9777 0.00764286
R54387 VCC.n9792 VCC.n9527 0.00764286
R54388 VCC.n9793 VCC.n9524 0.00764286
R54389 VCC.n9798 VCC.n9797 0.00764286
R54390 VCC.n9826 VCC.n9513 0.00764286
R54391 VCC.n9871 VCC.n9491 0.00764286
R54392 VCC.n9901 VCC.n9477 0.00764286
R54393 VCC.n9940 VCC.n9451 0.00764286
R54394 VCC.n9874 VCC.n9487 0.00764286
R54395 VCC.n9904 VCC.n9903 0.00764286
R54396 VCC.n9911 VCC.n9470 0.00764286
R54397 VCC.n9907 VCC.n9906 0.00764286
R54398 VCC.n9930 VCC.n9458 0.00764286
R54399 VCC.n9944 VCC.n9452 0.00764286
R54400 VCC.n10466 VCC.n10029 0.00764286
R54401 VCC.n10010 VCC.n10009 0.00764286
R54402 VCC.n10431 VCC.n10043 0.00764286
R54403 VCC.n10469 VCC.n10468 0.00764286
R54404 VCC.n10462 VCC.n10461 0.00764286
R54405 VCC.n10473 VCC.n10022 0.00764286
R54406 VCC.n10481 VCC.n10480 0.00764286
R54407 VCC.n10007 VCC.n10003 0.00764286
R54408 VCC.n10097 VCC.n10091 0.00764286
R54409 VCC.n10384 VCC.n10383 0.00764286
R54410 VCC.n10380 VCC.n10065 0.00764286
R54411 VCC.n10391 VCC.n10053 0.00764286
R54412 VCC.n10334 VCC.n10333 0.00764286
R54413 VCC.n10348 VCC.n10083 0.00764286
R54414 VCC.n10349 VCC.n10080 0.00764286
R54415 VCC.n10354 VCC.n10353 0.00764286
R54416 VCC.n10382 VCC.n10069 0.00764286
R54417 VCC.n10428 VCC.n10047 0.00764286
R54418 VCC.n10202 VCC.n10157 0.00764286
R54419 VCC.n10217 VCC.n10216 0.00764286
R54420 VCC.n10257 VCC.n10255 0.00764286
R54421 VCC.n10254 VCC.n10126 0.00764286
R54422 VCC.n10265 VCC.n10115 0.00764286
R54423 VCC.n10173 VCC.n10170 0.00764286
R54424 VCC.n10215 VCC.n10156 0.00764286
R54425 VCC.n10225 VCC.n10153 0.00764286
R54426 VCC.n10241 VCC.n10145 0.00764286
R54427 VCC.n10260 VCC.n10129 0.00764286
R54428 VCC.n10256 VCC.n10127 0.00764286
R54429 VCC.n10752 VCC.n10707 0.00764286
R54430 VCC.n10767 VCC.n10766 0.00764286
R54431 VCC.n10807 VCC.n10805 0.00764286
R54432 VCC.n10804 VCC.n10676 0.00764286
R54433 VCC.n10815 VCC.n10665 0.00764286
R54434 VCC.n10723 VCC.n10720 0.00764286
R54435 VCC.n10765 VCC.n10706 0.00764286
R54436 VCC.n10775 VCC.n10703 0.00764286
R54437 VCC.n10791 VCC.n10695 0.00764286
R54438 VCC.n10810 VCC.n10679 0.00764286
R54439 VCC.n10806 VCC.n10677 0.00764286
R54440 VCC.n10648 VCC.n10642 0.00764286
R54441 VCC.n10935 VCC.n10934 0.00764286
R54442 VCC.n10931 VCC.n10616 0.00764286
R54443 VCC.n10942 VCC.n10604 0.00764286
R54444 VCC.n10885 VCC.n10884 0.00764286
R54445 VCC.n10899 VCC.n10634 0.00764286
R54446 VCC.n10900 VCC.n10631 0.00764286
R54447 VCC.n10905 VCC.n10904 0.00764286
R54448 VCC.n10933 VCC.n10620 0.00764286
R54449 VCC.n10978 VCC.n10598 0.00764286
R54450 VCC.n11008 VCC.n10584 0.00764286
R54451 VCC.n11047 VCC.n10558 0.00764286
R54452 VCC.n10981 VCC.n10594 0.00764286
R54453 VCC.n11011 VCC.n11010 0.00764286
R54454 VCC.n11018 VCC.n10577 0.00764286
R54455 VCC.n11014 VCC.n11013 0.00764286
R54456 VCC.n11037 VCC.n10565 0.00764286
R54457 VCC.n11051 VCC.n10559 0.00764286
R54458 VCC.n11573 VCC.n11136 0.00764286
R54459 VCC.n11117 VCC.n11116 0.00764286
R54460 VCC.n11538 VCC.n11150 0.00764286
R54461 VCC.n11576 VCC.n11575 0.00764286
R54462 VCC.n11569 VCC.n11568 0.00764286
R54463 VCC.n11580 VCC.n11129 0.00764286
R54464 VCC.n11588 VCC.n11587 0.00764286
R54465 VCC.n11114 VCC.n11110 0.00764286
R54466 VCC.n11204 VCC.n11198 0.00764286
R54467 VCC.n11491 VCC.n11490 0.00764286
R54468 VCC.n11487 VCC.n11172 0.00764286
R54469 VCC.n11498 VCC.n11160 0.00764286
R54470 VCC.n11441 VCC.n11440 0.00764286
R54471 VCC.n11455 VCC.n11190 0.00764286
R54472 VCC.n11456 VCC.n11187 0.00764286
R54473 VCC.n11461 VCC.n11460 0.00764286
R54474 VCC.n11489 VCC.n11176 0.00764286
R54475 VCC.n11535 VCC.n11154 0.00764286
R54476 VCC.n11309 VCC.n11264 0.00764286
R54477 VCC.n11324 VCC.n11323 0.00764286
R54478 VCC.n11364 VCC.n11362 0.00764286
R54479 VCC.n11361 VCC.n11233 0.00764286
R54480 VCC.n11372 VCC.n11222 0.00764286
R54481 VCC.n11280 VCC.n11277 0.00764286
R54482 VCC.n11322 VCC.n11263 0.00764286
R54483 VCC.n11332 VCC.n11260 0.00764286
R54484 VCC.n11348 VCC.n11252 0.00764286
R54485 VCC.n11367 VCC.n11236 0.00764286
R54486 VCC.n11363 VCC.n11234 0.00764286
R54487 VCC.n11859 VCC.n11814 0.00764286
R54488 VCC.n11874 VCC.n11873 0.00764286
R54489 VCC.n11914 VCC.n11912 0.00764286
R54490 VCC.n11911 VCC.n11783 0.00764286
R54491 VCC.n11922 VCC.n11772 0.00764286
R54492 VCC.n11830 VCC.n11827 0.00764286
R54493 VCC.n11872 VCC.n11813 0.00764286
R54494 VCC.n11882 VCC.n11810 0.00764286
R54495 VCC.n11898 VCC.n11802 0.00764286
R54496 VCC.n11917 VCC.n11786 0.00764286
R54497 VCC.n11913 VCC.n11784 0.00764286
R54498 VCC.n11755 VCC.n11749 0.00764286
R54499 VCC.n12042 VCC.n12041 0.00764286
R54500 VCC.n12038 VCC.n11723 0.00764286
R54501 VCC.n12049 VCC.n11711 0.00764286
R54502 VCC.n11992 VCC.n11991 0.00764286
R54503 VCC.n12006 VCC.n11741 0.00764286
R54504 VCC.n12007 VCC.n11738 0.00764286
R54505 VCC.n12012 VCC.n12011 0.00764286
R54506 VCC.n12040 VCC.n11727 0.00764286
R54507 VCC.n12085 VCC.n11705 0.00764286
R54508 VCC.n12115 VCC.n11691 0.00764286
R54509 VCC.n12154 VCC.n11665 0.00764286
R54510 VCC.n12088 VCC.n11701 0.00764286
R54511 VCC.n12118 VCC.n12117 0.00764286
R54512 VCC.n12125 VCC.n11684 0.00764286
R54513 VCC.n12121 VCC.n12120 0.00764286
R54514 VCC.n12144 VCC.n11672 0.00764286
R54515 VCC.n12158 VCC.n11666 0.00764286
R54516 VCC.n12680 VCC.n12243 0.00764286
R54517 VCC.n12224 VCC.n12223 0.00764286
R54518 VCC.n12645 VCC.n12257 0.00764286
R54519 VCC.n12683 VCC.n12682 0.00764286
R54520 VCC.n12676 VCC.n12675 0.00764286
R54521 VCC.n12687 VCC.n12236 0.00764286
R54522 VCC.n12695 VCC.n12694 0.00764286
R54523 VCC.n12221 VCC.n12217 0.00764286
R54524 VCC.n12311 VCC.n12305 0.00764286
R54525 VCC.n12598 VCC.n12597 0.00764286
R54526 VCC.n12594 VCC.n12279 0.00764286
R54527 VCC.n12605 VCC.n12267 0.00764286
R54528 VCC.n12548 VCC.n12547 0.00764286
R54529 VCC.n12562 VCC.n12297 0.00764286
R54530 VCC.n12563 VCC.n12294 0.00764286
R54531 VCC.n12568 VCC.n12567 0.00764286
R54532 VCC.n12596 VCC.n12283 0.00764286
R54533 VCC.n12642 VCC.n12261 0.00764286
R54534 VCC.n12416 VCC.n12371 0.00764286
R54535 VCC.n12431 VCC.n12430 0.00764286
R54536 VCC.n12471 VCC.n12469 0.00764286
R54537 VCC.n12468 VCC.n12340 0.00764286
R54538 VCC.n12479 VCC.n12329 0.00764286
R54539 VCC.n12387 VCC.n12384 0.00764286
R54540 VCC.n12429 VCC.n12370 0.00764286
R54541 VCC.n12439 VCC.n12367 0.00764286
R54542 VCC.n12455 VCC.n12359 0.00764286
R54543 VCC.n12474 VCC.n12343 0.00764286
R54544 VCC.n12470 VCC.n12341 0.00764286
R54545 VCC.n12966 VCC.n12921 0.00764286
R54546 VCC.n12981 VCC.n12980 0.00764286
R54547 VCC.n13021 VCC.n13019 0.00764286
R54548 VCC.n13018 VCC.n12890 0.00764286
R54549 VCC.n13029 VCC.n12879 0.00764286
R54550 VCC.n12937 VCC.n12934 0.00764286
R54551 VCC.n12979 VCC.n12920 0.00764286
R54552 VCC.n12989 VCC.n12917 0.00764286
R54553 VCC.n13005 VCC.n12909 0.00764286
R54554 VCC.n13024 VCC.n12893 0.00764286
R54555 VCC.n13020 VCC.n12891 0.00764286
R54556 VCC.n12862 VCC.n12856 0.00764286
R54557 VCC.n13149 VCC.n13148 0.00764286
R54558 VCC.n13145 VCC.n12830 0.00764286
R54559 VCC.n13156 VCC.n12818 0.00764286
R54560 VCC.n13099 VCC.n13098 0.00764286
R54561 VCC.n13113 VCC.n12848 0.00764286
R54562 VCC.n13114 VCC.n12845 0.00764286
R54563 VCC.n13119 VCC.n13118 0.00764286
R54564 VCC.n13147 VCC.n12834 0.00764286
R54565 VCC.n13192 VCC.n12812 0.00764286
R54566 VCC.n13222 VCC.n12798 0.00764286
R54567 VCC.n13261 VCC.n12772 0.00764286
R54568 VCC.n13195 VCC.n12808 0.00764286
R54569 VCC.n13225 VCC.n13224 0.00764286
R54570 VCC.n13232 VCC.n12791 0.00764286
R54571 VCC.n13228 VCC.n13227 0.00764286
R54572 VCC.n13251 VCC.n12779 0.00764286
R54573 VCC.n13265 VCC.n12773 0.00764286
R54574 VCC.n13787 VCC.n13350 0.00764286
R54575 VCC.n13331 VCC.n13330 0.00764286
R54576 VCC.n13752 VCC.n13364 0.00764286
R54577 VCC.n13790 VCC.n13789 0.00764286
R54578 VCC.n13783 VCC.n13782 0.00764286
R54579 VCC.n13794 VCC.n13343 0.00764286
R54580 VCC.n13802 VCC.n13801 0.00764286
R54581 VCC.n13328 VCC.n13324 0.00764286
R54582 VCC.n13418 VCC.n13412 0.00764286
R54583 VCC.n13705 VCC.n13704 0.00764286
R54584 VCC.n13701 VCC.n13386 0.00764286
R54585 VCC.n13712 VCC.n13374 0.00764286
R54586 VCC.n13655 VCC.n13654 0.00764286
R54587 VCC.n13669 VCC.n13404 0.00764286
R54588 VCC.n13670 VCC.n13401 0.00764286
R54589 VCC.n13675 VCC.n13674 0.00764286
R54590 VCC.n13703 VCC.n13390 0.00764286
R54591 VCC.n13749 VCC.n13368 0.00764286
R54592 VCC.n13523 VCC.n13478 0.00764286
R54593 VCC.n13538 VCC.n13537 0.00764286
R54594 VCC.n13578 VCC.n13576 0.00764286
R54595 VCC.n13575 VCC.n13447 0.00764286
R54596 VCC.n13586 VCC.n13436 0.00764286
R54597 VCC.n13494 VCC.n13491 0.00764286
R54598 VCC.n13536 VCC.n13477 0.00764286
R54599 VCC.n13546 VCC.n13474 0.00764286
R54600 VCC.n13562 VCC.n13466 0.00764286
R54601 VCC.n13581 VCC.n13450 0.00764286
R54602 VCC.n13577 VCC.n13448 0.00764286
R54603 VCC.n14073 VCC.n14028 0.00764286
R54604 VCC.n14088 VCC.n14087 0.00764286
R54605 VCC.n14128 VCC.n14126 0.00764286
R54606 VCC.n14125 VCC.n13997 0.00764286
R54607 VCC.n14136 VCC.n13986 0.00764286
R54608 VCC.n14044 VCC.n14041 0.00764286
R54609 VCC.n14086 VCC.n14027 0.00764286
R54610 VCC.n14096 VCC.n14024 0.00764286
R54611 VCC.n14112 VCC.n14016 0.00764286
R54612 VCC.n14131 VCC.n14000 0.00764286
R54613 VCC.n14127 VCC.n13998 0.00764286
R54614 VCC.n13969 VCC.n13963 0.00764286
R54615 VCC.n14256 VCC.n14255 0.00764286
R54616 VCC.n14252 VCC.n13937 0.00764286
R54617 VCC.n14263 VCC.n13925 0.00764286
R54618 VCC.n14206 VCC.n14205 0.00764286
R54619 VCC.n14220 VCC.n13955 0.00764286
R54620 VCC.n14221 VCC.n13952 0.00764286
R54621 VCC.n14226 VCC.n14225 0.00764286
R54622 VCC.n14254 VCC.n13941 0.00764286
R54623 VCC.n14299 VCC.n13919 0.00764286
R54624 VCC.n14329 VCC.n13905 0.00764286
R54625 VCC.n14368 VCC.n13879 0.00764286
R54626 VCC.n14302 VCC.n13915 0.00764286
R54627 VCC.n14332 VCC.n14331 0.00764286
R54628 VCC.n14339 VCC.n13898 0.00764286
R54629 VCC.n14335 VCC.n14334 0.00764286
R54630 VCC.n14358 VCC.n13886 0.00764286
R54631 VCC.n14372 VCC.n13880 0.00764286
R54632 VCC.n14894 VCC.n14457 0.00764286
R54633 VCC.n14438 VCC.n14437 0.00764286
R54634 VCC.n14859 VCC.n14471 0.00764286
R54635 VCC.n14897 VCC.n14896 0.00764286
R54636 VCC.n14890 VCC.n14889 0.00764286
R54637 VCC.n14901 VCC.n14450 0.00764286
R54638 VCC.n14909 VCC.n14908 0.00764286
R54639 VCC.n14435 VCC.n14431 0.00764286
R54640 VCC.n14525 VCC.n14519 0.00764286
R54641 VCC.n14812 VCC.n14811 0.00764286
R54642 VCC.n14808 VCC.n14493 0.00764286
R54643 VCC.n14819 VCC.n14481 0.00764286
R54644 VCC.n14762 VCC.n14761 0.00764286
R54645 VCC.n14776 VCC.n14511 0.00764286
R54646 VCC.n14777 VCC.n14508 0.00764286
R54647 VCC.n14782 VCC.n14781 0.00764286
R54648 VCC.n14810 VCC.n14497 0.00764286
R54649 VCC.n14856 VCC.n14475 0.00764286
R54650 VCC.n14630 VCC.n14585 0.00764286
R54651 VCC.n14645 VCC.n14644 0.00764286
R54652 VCC.n14685 VCC.n14683 0.00764286
R54653 VCC.n14682 VCC.n14554 0.00764286
R54654 VCC.n14693 VCC.n14543 0.00764286
R54655 VCC.n14601 VCC.n14598 0.00764286
R54656 VCC.n14643 VCC.n14584 0.00764286
R54657 VCC.n14653 VCC.n14581 0.00764286
R54658 VCC.n14669 VCC.n14573 0.00764286
R54659 VCC.n14688 VCC.n14557 0.00764286
R54660 VCC.n14684 VCC.n14555 0.00764286
R54661 VCC.n15180 VCC.n15135 0.00764286
R54662 VCC.n15195 VCC.n15194 0.00764286
R54663 VCC.n15235 VCC.n15233 0.00764286
R54664 VCC.n15232 VCC.n15104 0.00764286
R54665 VCC.n15243 VCC.n15093 0.00764286
R54666 VCC.n15151 VCC.n15148 0.00764286
R54667 VCC.n15193 VCC.n15134 0.00764286
R54668 VCC.n15203 VCC.n15131 0.00764286
R54669 VCC.n15219 VCC.n15123 0.00764286
R54670 VCC.n15238 VCC.n15107 0.00764286
R54671 VCC.n15234 VCC.n15105 0.00764286
R54672 VCC.n15076 VCC.n15070 0.00764286
R54673 VCC.n15363 VCC.n15362 0.00764286
R54674 VCC.n15359 VCC.n15044 0.00764286
R54675 VCC.n15370 VCC.n15032 0.00764286
R54676 VCC.n15313 VCC.n15312 0.00764286
R54677 VCC.n15327 VCC.n15062 0.00764286
R54678 VCC.n15328 VCC.n15059 0.00764286
R54679 VCC.n15333 VCC.n15332 0.00764286
R54680 VCC.n15361 VCC.n15048 0.00764286
R54681 VCC.n15406 VCC.n15026 0.00764286
R54682 VCC.n15436 VCC.n15012 0.00764286
R54683 VCC.n15475 VCC.n14986 0.00764286
R54684 VCC.n15409 VCC.n15022 0.00764286
R54685 VCC.n15439 VCC.n15438 0.00764286
R54686 VCC.n15446 VCC.n15005 0.00764286
R54687 VCC.n15442 VCC.n15441 0.00764286
R54688 VCC.n15465 VCC.n14993 0.00764286
R54689 VCC.n15479 VCC.n14987 0.00764286
R54690 VCC.n16001 VCC.n15564 0.00764286
R54691 VCC.n15545 VCC.n15544 0.00764286
R54692 VCC.n15966 VCC.n15578 0.00764286
R54693 VCC.n16004 VCC.n16003 0.00764286
R54694 VCC.n15997 VCC.n15996 0.00764286
R54695 VCC.n16008 VCC.n15557 0.00764286
R54696 VCC.n16016 VCC.n16015 0.00764286
R54697 VCC.n15542 VCC.n15538 0.00764286
R54698 VCC.n15632 VCC.n15626 0.00764286
R54699 VCC.n15919 VCC.n15918 0.00764286
R54700 VCC.n15915 VCC.n15600 0.00764286
R54701 VCC.n15926 VCC.n15588 0.00764286
R54702 VCC.n15869 VCC.n15868 0.00764286
R54703 VCC.n15883 VCC.n15618 0.00764286
R54704 VCC.n15884 VCC.n15615 0.00764286
R54705 VCC.n15889 VCC.n15888 0.00764286
R54706 VCC.n15917 VCC.n15604 0.00764286
R54707 VCC.n15963 VCC.n15582 0.00764286
R54708 VCC.n15737 VCC.n15692 0.00764286
R54709 VCC.n15752 VCC.n15751 0.00764286
R54710 VCC.n15792 VCC.n15790 0.00764286
R54711 VCC.n15789 VCC.n15661 0.00764286
R54712 VCC.n15800 VCC.n15650 0.00764286
R54713 VCC.n15708 VCC.n15705 0.00764286
R54714 VCC.n15750 VCC.n15691 0.00764286
R54715 VCC.n15760 VCC.n15688 0.00764286
R54716 VCC.n15776 VCC.n15680 0.00764286
R54717 VCC.n15795 VCC.n15664 0.00764286
R54718 VCC.n15791 VCC.n15662 0.00764286
R54719 VCC.n16287 VCC.n16242 0.00764286
R54720 VCC.n16302 VCC.n16301 0.00764286
R54721 VCC.n16342 VCC.n16340 0.00764286
R54722 VCC.n16339 VCC.n16211 0.00764286
R54723 VCC.n16350 VCC.n16200 0.00764286
R54724 VCC.n16258 VCC.n16255 0.00764286
R54725 VCC.n16300 VCC.n16241 0.00764286
R54726 VCC.n16310 VCC.n16238 0.00764286
R54727 VCC.n16326 VCC.n16230 0.00764286
R54728 VCC.n16345 VCC.n16214 0.00764286
R54729 VCC.n16341 VCC.n16212 0.00764286
R54730 VCC.n16183 VCC.n16177 0.00764286
R54731 VCC.n16470 VCC.n16469 0.00764286
R54732 VCC.n16466 VCC.n16151 0.00764286
R54733 VCC.n16477 VCC.n16139 0.00764286
R54734 VCC.n16420 VCC.n16419 0.00764286
R54735 VCC.n16434 VCC.n16169 0.00764286
R54736 VCC.n16435 VCC.n16166 0.00764286
R54737 VCC.n16440 VCC.n16439 0.00764286
R54738 VCC.n16468 VCC.n16155 0.00764286
R54739 VCC.n16513 VCC.n16133 0.00764286
R54740 VCC.n16543 VCC.n16119 0.00764286
R54741 VCC.n16582 VCC.n16093 0.00764286
R54742 VCC.n16516 VCC.n16129 0.00764286
R54743 VCC.n16546 VCC.n16545 0.00764286
R54744 VCC.n16553 VCC.n16112 0.00764286
R54745 VCC.n16549 VCC.n16548 0.00764286
R54746 VCC.n16572 VCC.n16100 0.00764286
R54747 VCC.n16586 VCC.n16094 0.00764286
R54748 VCC.n17108 VCC.n16671 0.00764286
R54749 VCC.n16652 VCC.n16651 0.00764286
R54750 VCC.n17073 VCC.n16685 0.00764286
R54751 VCC.n17111 VCC.n17110 0.00764286
R54752 VCC.n17104 VCC.n17103 0.00764286
R54753 VCC.n17115 VCC.n16664 0.00764286
R54754 VCC.n17123 VCC.n17122 0.00764286
R54755 VCC.n16649 VCC.n16645 0.00764286
R54756 VCC.n16739 VCC.n16733 0.00764286
R54757 VCC.n17026 VCC.n17025 0.00764286
R54758 VCC.n17022 VCC.n16707 0.00764286
R54759 VCC.n17033 VCC.n16695 0.00764286
R54760 VCC.n16976 VCC.n16975 0.00764286
R54761 VCC.n16990 VCC.n16725 0.00764286
R54762 VCC.n16991 VCC.n16722 0.00764286
R54763 VCC.n16996 VCC.n16995 0.00764286
R54764 VCC.n17024 VCC.n16711 0.00764286
R54765 VCC.n17070 VCC.n16689 0.00764286
R54766 VCC.n16844 VCC.n16799 0.00764286
R54767 VCC.n16859 VCC.n16858 0.00764286
R54768 VCC.n16899 VCC.n16897 0.00764286
R54769 VCC.n16896 VCC.n16768 0.00764286
R54770 VCC.n16907 VCC.n16757 0.00764286
R54771 VCC.n16815 VCC.n16812 0.00764286
R54772 VCC.n16857 VCC.n16798 0.00764286
R54773 VCC.n16867 VCC.n16795 0.00764286
R54774 VCC.n16883 VCC.n16787 0.00764286
R54775 VCC.n16902 VCC.n16771 0.00764286
R54776 VCC.n16898 VCC.n16769 0.00764286
R54777 VCC.n17290 VCC.n17284 0.00764286
R54778 VCC.n17390 VCC.n17389 0.00764286
R54779 VCC.n17386 VCC.n17258 0.00764286
R54780 VCC.n17397 VCC.n17246 0.00764286
R54781 VCC.n17340 VCC.n17339 0.00764286
R54782 VCC.n17354 VCC.n17276 0.00764286
R54783 VCC.n17355 VCC.n17273 0.00764286
R54784 VCC.n17360 VCC.n17359 0.00764286
R54785 VCC.n17388 VCC.n17262 0.00764286
R54786 VCC.n17433 VCC.n17240 0.00764286
R54787 VCC.n17463 VCC.n17226 0.00764286
R54788 VCC.n17502 VCC.n17200 0.00764286
R54789 VCC.n17436 VCC.n17236 0.00764286
R54790 VCC.n17466 VCC.n17465 0.00764286
R54791 VCC.n17473 VCC.n17219 0.00764286
R54792 VCC.n17469 VCC.n17468 0.00764286
R54793 VCC.n17492 VCC.n17207 0.00764286
R54794 VCC.n17506 VCC.n17201 0.00764286
R54795 VCC.n203 VCC.n196 0.00675
R54796 VCC.n246 VCC.n170 0.00675
R54797 VCC.n277 VCC.n276 0.00675
R54798 VCC.n298 VCC.n138 0.00675
R54799 VCC.n239 VCC.n175 0.00675
R54800 VCC.n245 VCC.n171 0.00675
R54801 VCC.n275 VCC.n149 0.00675
R54802 VCC.n283 VCC.n132 0.00675
R54803 VCC.n312 VCC.n128 0.00675
R54804 VCC.n352 VCC.n351 0.00675
R54805 VCC.n367 VCC.n104 0.00675
R54806 VCC.n403 VCC.n401 0.00675
R54807 VCC.n433 VCC.n77 0.00675
R54808 VCC.n314 VCC.n126 0.00675
R54809 VCC.n345 VCC.n113 0.00675
R54810 VCC.n353 VCC.n349 0.00675
R54811 VCC.n406 VCC.n88 0.00675
R54812 VCC.n402 VCC.n86 0.00675
R54813 VCC.n53 VCC.n44 0.00675
R54814 VCC.n47 VCC.n45 0.00675
R54815 VCC.n521 VCC.n27 0.00675
R54816 VCC.n51 VCC.n46 0.00675
R54817 VCC.n486 VCC.n48 0.00675
R54818 VCC.n34 VCC.n31 0.00675
R54819 VCC.n520 VCC.n519 0.00675
R54820 VCC.n518 VCC.n514 0.00675
R54821 VCC.n755 VCC.n748 0.00675
R54822 VCC.n798 VCC.n722 0.00675
R54823 VCC.n829 VCC.n828 0.00675
R54824 VCC.n850 VCC.n690 0.00675
R54825 VCC.n791 VCC.n727 0.00675
R54826 VCC.n797 VCC.n723 0.00675
R54827 VCC.n827 VCC.n701 0.00675
R54828 VCC.n835 VCC.n684 0.00675
R54829 VCC.n864 VCC.n680 0.00675
R54830 VCC.n904 VCC.n903 0.00675
R54831 VCC.n919 VCC.n656 0.00675
R54832 VCC.n955 VCC.n953 0.00675
R54833 VCC.n985 VCC.n629 0.00675
R54834 VCC.n866 VCC.n678 0.00675
R54835 VCC.n897 VCC.n665 0.00675
R54836 VCC.n905 VCC.n901 0.00675
R54837 VCC.n958 VCC.n640 0.00675
R54838 VCC.n954 VCC.n638 0.00675
R54839 VCC.n605 VCC.n596 0.00675
R54840 VCC.n599 VCC.n597 0.00675
R54841 VCC.n1073 VCC.n579 0.00675
R54842 VCC.n603 VCC.n598 0.00675
R54843 VCC.n1038 VCC.n600 0.00675
R54844 VCC.n586 VCC.n583 0.00675
R54845 VCC.n1072 VCC.n1071 0.00675
R54846 VCC.n1070 VCC.n1066 0.00675
R54847 VCC.n1592 VCC.n1158 0.00675
R54848 VCC.n1604 VCC.n1152 0.00675
R54849 VCC.n1138 VCC.n1134 0.00675
R54850 VCC.n1591 VCC.n1156 0.00675
R54851 VCC.n1603 VCC.n1153 0.00675
R54852 VCC.n1609 VCC.n1131 0.00675
R54853 VCC.n1137 VCC.n1136 0.00675
R54854 VCC.n1630 VCC.n1129 0.00675
R54855 VCC.n1461 VCC.n1460 0.00675
R54856 VCC.n1476 VCC.n1213 0.00675
R54857 VCC.n1512 VCC.n1510 0.00675
R54858 VCC.n1543 VCC.n1186 0.00675
R54859 VCC.n1424 VCC.n1236 0.00675
R54860 VCC.n1454 VCC.n1222 0.00675
R54861 VCC.n1462 VCC.n1458 0.00675
R54862 VCC.n1515 VCC.n1197 0.00675
R54863 VCC.n1511 VCC.n1195 0.00675
R54864 VCC.n1313 VCC.n1306 0.00675
R54865 VCC.n1356 VCC.n1280 0.00675
R54866 VCC.n1387 VCC.n1386 0.00675
R54867 VCC.n1408 VCC.n1248 0.00675
R54868 VCC.n1349 VCC.n1285 0.00675
R54869 VCC.n1355 VCC.n1281 0.00675
R54870 VCC.n1385 VCC.n1259 0.00675
R54871 VCC.n1393 VCC.n1242 0.00675
R54872 VCC.n1422 VCC.n1238 0.00675
R54873 VCC.n1864 VCC.n1857 0.00675
R54874 VCC.n1907 VCC.n1831 0.00675
R54875 VCC.n1938 VCC.n1937 0.00675
R54876 VCC.n1959 VCC.n1799 0.00675
R54877 VCC.n1900 VCC.n1836 0.00675
R54878 VCC.n1906 VCC.n1832 0.00675
R54879 VCC.n1936 VCC.n1810 0.00675
R54880 VCC.n1944 VCC.n1793 0.00675
R54881 VCC.n1973 VCC.n1789 0.00675
R54882 VCC.n2013 VCC.n2012 0.00675
R54883 VCC.n2028 VCC.n1765 0.00675
R54884 VCC.n2064 VCC.n2062 0.00675
R54885 VCC.n2094 VCC.n1738 0.00675
R54886 VCC.n1975 VCC.n1787 0.00675
R54887 VCC.n2006 VCC.n1774 0.00675
R54888 VCC.n2014 VCC.n2010 0.00675
R54889 VCC.n2067 VCC.n1749 0.00675
R54890 VCC.n2063 VCC.n1747 0.00675
R54891 VCC.n1714 VCC.n1705 0.00675
R54892 VCC.n1708 VCC.n1706 0.00675
R54893 VCC.n2182 VCC.n1688 0.00675
R54894 VCC.n1712 VCC.n1707 0.00675
R54895 VCC.n2147 VCC.n1709 0.00675
R54896 VCC.n1695 VCC.n1692 0.00675
R54897 VCC.n2181 VCC.n2180 0.00675
R54898 VCC.n2179 VCC.n2175 0.00675
R54899 VCC.n2701 VCC.n2267 0.00675
R54900 VCC.n2713 VCC.n2261 0.00675
R54901 VCC.n2247 VCC.n2243 0.00675
R54902 VCC.n2700 VCC.n2265 0.00675
R54903 VCC.n2712 VCC.n2262 0.00675
R54904 VCC.n2718 VCC.n2240 0.00675
R54905 VCC.n2246 VCC.n2245 0.00675
R54906 VCC.n2739 VCC.n2238 0.00675
R54907 VCC.n2570 VCC.n2569 0.00675
R54908 VCC.n2585 VCC.n2322 0.00675
R54909 VCC.n2621 VCC.n2619 0.00675
R54910 VCC.n2652 VCC.n2295 0.00675
R54911 VCC.n2533 VCC.n2345 0.00675
R54912 VCC.n2563 VCC.n2331 0.00675
R54913 VCC.n2571 VCC.n2567 0.00675
R54914 VCC.n2624 VCC.n2306 0.00675
R54915 VCC.n2620 VCC.n2304 0.00675
R54916 VCC.n2422 VCC.n2415 0.00675
R54917 VCC.n2465 VCC.n2389 0.00675
R54918 VCC.n2496 VCC.n2495 0.00675
R54919 VCC.n2517 VCC.n2357 0.00675
R54920 VCC.n2458 VCC.n2394 0.00675
R54921 VCC.n2464 VCC.n2390 0.00675
R54922 VCC.n2494 VCC.n2368 0.00675
R54923 VCC.n2502 VCC.n2351 0.00675
R54924 VCC.n2531 VCC.n2347 0.00675
R54925 VCC.n2973 VCC.n2966 0.00675
R54926 VCC.n3016 VCC.n2940 0.00675
R54927 VCC.n3047 VCC.n3046 0.00675
R54928 VCC.n3068 VCC.n2908 0.00675
R54929 VCC.n3009 VCC.n2945 0.00675
R54930 VCC.n3015 VCC.n2941 0.00675
R54931 VCC.n3045 VCC.n2919 0.00675
R54932 VCC.n3053 VCC.n2902 0.00675
R54933 VCC.n3082 VCC.n2898 0.00675
R54934 VCC.n3122 VCC.n3121 0.00675
R54935 VCC.n3137 VCC.n2874 0.00675
R54936 VCC.n3173 VCC.n3171 0.00675
R54937 VCC.n3203 VCC.n2847 0.00675
R54938 VCC.n3084 VCC.n2896 0.00675
R54939 VCC.n3115 VCC.n2883 0.00675
R54940 VCC.n3123 VCC.n3119 0.00675
R54941 VCC.n3176 VCC.n2858 0.00675
R54942 VCC.n3172 VCC.n2856 0.00675
R54943 VCC.n2823 VCC.n2814 0.00675
R54944 VCC.n2817 VCC.n2815 0.00675
R54945 VCC.n3291 VCC.n2797 0.00675
R54946 VCC.n2821 VCC.n2816 0.00675
R54947 VCC.n3256 VCC.n2818 0.00675
R54948 VCC.n2804 VCC.n2801 0.00675
R54949 VCC.n3290 VCC.n3289 0.00675
R54950 VCC.n3288 VCC.n3284 0.00675
R54951 VCC.n3810 VCC.n3376 0.00675
R54952 VCC.n3822 VCC.n3370 0.00675
R54953 VCC.n3356 VCC.n3352 0.00675
R54954 VCC.n3809 VCC.n3374 0.00675
R54955 VCC.n3821 VCC.n3371 0.00675
R54956 VCC.n3827 VCC.n3349 0.00675
R54957 VCC.n3355 VCC.n3354 0.00675
R54958 VCC.n3848 VCC.n3347 0.00675
R54959 VCC.n3679 VCC.n3678 0.00675
R54960 VCC.n3694 VCC.n3431 0.00675
R54961 VCC.n3730 VCC.n3728 0.00675
R54962 VCC.n3761 VCC.n3404 0.00675
R54963 VCC.n3642 VCC.n3454 0.00675
R54964 VCC.n3672 VCC.n3440 0.00675
R54965 VCC.n3680 VCC.n3676 0.00675
R54966 VCC.n3733 VCC.n3415 0.00675
R54967 VCC.n3729 VCC.n3413 0.00675
R54968 VCC.n3531 VCC.n3524 0.00675
R54969 VCC.n3574 VCC.n3498 0.00675
R54970 VCC.n3605 VCC.n3604 0.00675
R54971 VCC.n3626 VCC.n3466 0.00675
R54972 VCC.n3567 VCC.n3503 0.00675
R54973 VCC.n3573 VCC.n3499 0.00675
R54974 VCC.n3603 VCC.n3477 0.00675
R54975 VCC.n3611 VCC.n3460 0.00675
R54976 VCC.n3640 VCC.n3456 0.00675
R54977 VCC.n4082 VCC.n4075 0.00675
R54978 VCC.n4125 VCC.n4049 0.00675
R54979 VCC.n4156 VCC.n4155 0.00675
R54980 VCC.n4177 VCC.n4017 0.00675
R54981 VCC.n4118 VCC.n4054 0.00675
R54982 VCC.n4124 VCC.n4050 0.00675
R54983 VCC.n4154 VCC.n4028 0.00675
R54984 VCC.n4162 VCC.n4011 0.00675
R54985 VCC.n4191 VCC.n4007 0.00675
R54986 VCC.n4231 VCC.n4230 0.00675
R54987 VCC.n4246 VCC.n3983 0.00675
R54988 VCC.n4282 VCC.n4280 0.00675
R54989 VCC.n4312 VCC.n3956 0.00675
R54990 VCC.n4193 VCC.n4005 0.00675
R54991 VCC.n4224 VCC.n3992 0.00675
R54992 VCC.n4232 VCC.n4228 0.00675
R54993 VCC.n4285 VCC.n3967 0.00675
R54994 VCC.n4281 VCC.n3965 0.00675
R54995 VCC.n3932 VCC.n3923 0.00675
R54996 VCC.n3926 VCC.n3924 0.00675
R54997 VCC.n4400 VCC.n3906 0.00675
R54998 VCC.n3930 VCC.n3925 0.00675
R54999 VCC.n4365 VCC.n3927 0.00675
R55000 VCC.n3913 VCC.n3910 0.00675
R55001 VCC.n4399 VCC.n4398 0.00675
R55002 VCC.n4397 VCC.n4393 0.00675
R55003 VCC.n4919 VCC.n4485 0.00675
R55004 VCC.n4931 VCC.n4479 0.00675
R55005 VCC.n4465 VCC.n4461 0.00675
R55006 VCC.n4918 VCC.n4483 0.00675
R55007 VCC.n4930 VCC.n4480 0.00675
R55008 VCC.n4936 VCC.n4458 0.00675
R55009 VCC.n4464 VCC.n4463 0.00675
R55010 VCC.n4957 VCC.n4456 0.00675
R55011 VCC.n4788 VCC.n4787 0.00675
R55012 VCC.n4803 VCC.n4540 0.00675
R55013 VCC.n4839 VCC.n4837 0.00675
R55014 VCC.n4870 VCC.n4513 0.00675
R55015 VCC.n4751 VCC.n4563 0.00675
R55016 VCC.n4781 VCC.n4549 0.00675
R55017 VCC.n4789 VCC.n4785 0.00675
R55018 VCC.n4842 VCC.n4524 0.00675
R55019 VCC.n4838 VCC.n4522 0.00675
R55020 VCC.n4640 VCC.n4633 0.00675
R55021 VCC.n4683 VCC.n4607 0.00675
R55022 VCC.n4714 VCC.n4713 0.00675
R55023 VCC.n4735 VCC.n4575 0.00675
R55024 VCC.n4676 VCC.n4612 0.00675
R55025 VCC.n4682 VCC.n4608 0.00675
R55026 VCC.n4712 VCC.n4586 0.00675
R55027 VCC.n4720 VCC.n4569 0.00675
R55028 VCC.n4749 VCC.n4565 0.00675
R55029 VCC.n5191 VCC.n5184 0.00675
R55030 VCC.n5234 VCC.n5158 0.00675
R55031 VCC.n5265 VCC.n5264 0.00675
R55032 VCC.n5286 VCC.n5126 0.00675
R55033 VCC.n5227 VCC.n5163 0.00675
R55034 VCC.n5233 VCC.n5159 0.00675
R55035 VCC.n5263 VCC.n5137 0.00675
R55036 VCC.n5271 VCC.n5120 0.00675
R55037 VCC.n5300 VCC.n5116 0.00675
R55038 VCC.n5340 VCC.n5339 0.00675
R55039 VCC.n5355 VCC.n5092 0.00675
R55040 VCC.n5391 VCC.n5389 0.00675
R55041 VCC.n5421 VCC.n5065 0.00675
R55042 VCC.n5302 VCC.n5114 0.00675
R55043 VCC.n5333 VCC.n5101 0.00675
R55044 VCC.n5341 VCC.n5337 0.00675
R55045 VCC.n5394 VCC.n5076 0.00675
R55046 VCC.n5390 VCC.n5074 0.00675
R55047 VCC.n5041 VCC.n5032 0.00675
R55048 VCC.n5035 VCC.n5033 0.00675
R55049 VCC.n5509 VCC.n5015 0.00675
R55050 VCC.n5039 VCC.n5034 0.00675
R55051 VCC.n5474 VCC.n5036 0.00675
R55052 VCC.n5022 VCC.n5019 0.00675
R55053 VCC.n5508 VCC.n5507 0.00675
R55054 VCC.n5506 VCC.n5502 0.00675
R55055 VCC.n6028 VCC.n5594 0.00675
R55056 VCC.n6040 VCC.n5588 0.00675
R55057 VCC.n5574 VCC.n5570 0.00675
R55058 VCC.n6027 VCC.n5592 0.00675
R55059 VCC.n6039 VCC.n5589 0.00675
R55060 VCC.n6045 VCC.n5567 0.00675
R55061 VCC.n5573 VCC.n5572 0.00675
R55062 VCC.n6066 VCC.n5565 0.00675
R55063 VCC.n5897 VCC.n5896 0.00675
R55064 VCC.n5912 VCC.n5649 0.00675
R55065 VCC.n5948 VCC.n5946 0.00675
R55066 VCC.n5979 VCC.n5622 0.00675
R55067 VCC.n5860 VCC.n5672 0.00675
R55068 VCC.n5890 VCC.n5658 0.00675
R55069 VCC.n5898 VCC.n5894 0.00675
R55070 VCC.n5951 VCC.n5633 0.00675
R55071 VCC.n5947 VCC.n5631 0.00675
R55072 VCC.n5749 VCC.n5742 0.00675
R55073 VCC.n5792 VCC.n5716 0.00675
R55074 VCC.n5823 VCC.n5822 0.00675
R55075 VCC.n5844 VCC.n5684 0.00675
R55076 VCC.n5785 VCC.n5721 0.00675
R55077 VCC.n5791 VCC.n5717 0.00675
R55078 VCC.n5821 VCC.n5695 0.00675
R55079 VCC.n5829 VCC.n5678 0.00675
R55080 VCC.n5858 VCC.n5674 0.00675
R55081 VCC.n6300 VCC.n6293 0.00675
R55082 VCC.n6343 VCC.n6267 0.00675
R55083 VCC.n6374 VCC.n6373 0.00675
R55084 VCC.n6395 VCC.n6235 0.00675
R55085 VCC.n6336 VCC.n6272 0.00675
R55086 VCC.n6342 VCC.n6268 0.00675
R55087 VCC.n6372 VCC.n6246 0.00675
R55088 VCC.n6380 VCC.n6229 0.00675
R55089 VCC.n6409 VCC.n6225 0.00675
R55090 VCC.n6449 VCC.n6448 0.00675
R55091 VCC.n6464 VCC.n6201 0.00675
R55092 VCC.n6500 VCC.n6498 0.00675
R55093 VCC.n6530 VCC.n6174 0.00675
R55094 VCC.n6411 VCC.n6223 0.00675
R55095 VCC.n6442 VCC.n6210 0.00675
R55096 VCC.n6450 VCC.n6446 0.00675
R55097 VCC.n6503 VCC.n6185 0.00675
R55098 VCC.n6499 VCC.n6183 0.00675
R55099 VCC.n6150 VCC.n6141 0.00675
R55100 VCC.n6144 VCC.n6142 0.00675
R55101 VCC.n6618 VCC.n6124 0.00675
R55102 VCC.n6148 VCC.n6143 0.00675
R55103 VCC.n6583 VCC.n6145 0.00675
R55104 VCC.n6131 VCC.n6128 0.00675
R55105 VCC.n6617 VCC.n6616 0.00675
R55106 VCC.n6615 VCC.n6611 0.00675
R55107 VCC.n7137 VCC.n6703 0.00675
R55108 VCC.n7149 VCC.n6697 0.00675
R55109 VCC.n6683 VCC.n6679 0.00675
R55110 VCC.n7136 VCC.n6701 0.00675
R55111 VCC.n7148 VCC.n6698 0.00675
R55112 VCC.n7154 VCC.n6676 0.00675
R55113 VCC.n6682 VCC.n6681 0.00675
R55114 VCC.n7175 VCC.n6674 0.00675
R55115 VCC.n7006 VCC.n7005 0.00675
R55116 VCC.n7021 VCC.n6758 0.00675
R55117 VCC.n7057 VCC.n7055 0.00675
R55118 VCC.n7088 VCC.n6731 0.00675
R55119 VCC.n6969 VCC.n6781 0.00675
R55120 VCC.n6999 VCC.n6767 0.00675
R55121 VCC.n7007 VCC.n7003 0.00675
R55122 VCC.n7060 VCC.n6742 0.00675
R55123 VCC.n7056 VCC.n6740 0.00675
R55124 VCC.n6858 VCC.n6851 0.00675
R55125 VCC.n6901 VCC.n6825 0.00675
R55126 VCC.n6932 VCC.n6931 0.00675
R55127 VCC.n6953 VCC.n6793 0.00675
R55128 VCC.n6894 VCC.n6830 0.00675
R55129 VCC.n6900 VCC.n6826 0.00675
R55130 VCC.n6930 VCC.n6804 0.00675
R55131 VCC.n6938 VCC.n6787 0.00675
R55132 VCC.n6967 VCC.n6783 0.00675
R55133 VCC.n7409 VCC.n7402 0.00675
R55134 VCC.n7452 VCC.n7376 0.00675
R55135 VCC.n7483 VCC.n7482 0.00675
R55136 VCC.n7504 VCC.n7344 0.00675
R55137 VCC.n7445 VCC.n7381 0.00675
R55138 VCC.n7451 VCC.n7377 0.00675
R55139 VCC.n7481 VCC.n7355 0.00675
R55140 VCC.n7489 VCC.n7338 0.00675
R55141 VCC.n7518 VCC.n7334 0.00675
R55142 VCC.n7558 VCC.n7557 0.00675
R55143 VCC.n7573 VCC.n7310 0.00675
R55144 VCC.n7609 VCC.n7607 0.00675
R55145 VCC.n7639 VCC.n7283 0.00675
R55146 VCC.n7520 VCC.n7332 0.00675
R55147 VCC.n7551 VCC.n7319 0.00675
R55148 VCC.n7559 VCC.n7555 0.00675
R55149 VCC.n7612 VCC.n7294 0.00675
R55150 VCC.n7608 VCC.n7292 0.00675
R55151 VCC.n7259 VCC.n7250 0.00675
R55152 VCC.n7253 VCC.n7251 0.00675
R55153 VCC.n7727 VCC.n7233 0.00675
R55154 VCC.n7257 VCC.n7252 0.00675
R55155 VCC.n7692 VCC.n7254 0.00675
R55156 VCC.n7240 VCC.n7237 0.00675
R55157 VCC.n7726 VCC.n7725 0.00675
R55158 VCC.n7724 VCC.n7720 0.00675
R55159 VCC.n8246 VCC.n7812 0.00675
R55160 VCC.n8258 VCC.n7806 0.00675
R55161 VCC.n7792 VCC.n7788 0.00675
R55162 VCC.n8245 VCC.n7810 0.00675
R55163 VCC.n8257 VCC.n7807 0.00675
R55164 VCC.n8263 VCC.n7785 0.00675
R55165 VCC.n7791 VCC.n7790 0.00675
R55166 VCC.n8284 VCC.n7783 0.00675
R55167 VCC.n8115 VCC.n8114 0.00675
R55168 VCC.n8130 VCC.n7867 0.00675
R55169 VCC.n8166 VCC.n8164 0.00675
R55170 VCC.n8197 VCC.n7840 0.00675
R55171 VCC.n8078 VCC.n7890 0.00675
R55172 VCC.n8108 VCC.n7876 0.00675
R55173 VCC.n8116 VCC.n8112 0.00675
R55174 VCC.n8169 VCC.n7851 0.00675
R55175 VCC.n8165 VCC.n7849 0.00675
R55176 VCC.n7967 VCC.n7960 0.00675
R55177 VCC.n8010 VCC.n7934 0.00675
R55178 VCC.n8041 VCC.n8040 0.00675
R55179 VCC.n8062 VCC.n7902 0.00675
R55180 VCC.n8003 VCC.n7939 0.00675
R55181 VCC.n8009 VCC.n7935 0.00675
R55182 VCC.n8039 VCC.n7913 0.00675
R55183 VCC.n8047 VCC.n7896 0.00675
R55184 VCC.n8076 VCC.n7892 0.00675
R55185 VCC.n8667 VCC.n8666 0.00675
R55186 VCC.n8682 VCC.n8419 0.00675
R55187 VCC.n8718 VCC.n8716 0.00675
R55188 VCC.n8748 VCC.n8392 0.00675
R55189 VCC.n8629 VCC.n8441 0.00675
R55190 VCC.n8660 VCC.n8428 0.00675
R55191 VCC.n8668 VCC.n8664 0.00675
R55192 VCC.n8721 VCC.n8403 0.00675
R55193 VCC.n8717 VCC.n8401 0.00675
R55194 VCC.n8368 VCC.n8359 0.00675
R55195 VCC.n8362 VCC.n8360 0.00675
R55196 VCC.n8836 VCC.n8342 0.00675
R55197 VCC.n8366 VCC.n8361 0.00675
R55198 VCC.n8801 VCC.n8363 0.00675
R55199 VCC.n8349 VCC.n8346 0.00675
R55200 VCC.n8835 VCC.n8834 0.00675
R55201 VCC.n8833 VCC.n8829 0.00675
R55202 VCC.n8518 VCC.n8511 0.00675
R55203 VCC.n8561 VCC.n8485 0.00675
R55204 VCC.n8592 VCC.n8591 0.00675
R55205 VCC.n8613 VCC.n8453 0.00675
R55206 VCC.n8554 VCC.n8490 0.00675
R55207 VCC.n8560 VCC.n8486 0.00675
R55208 VCC.n8590 VCC.n8464 0.00675
R55209 VCC.n8598 VCC.n8447 0.00675
R55210 VCC.n8627 VCC.n8443 0.00675
R55211 VCC.n9355 VCC.n8921 0.00675
R55212 VCC.n9367 VCC.n8915 0.00675
R55213 VCC.n8901 VCC.n8897 0.00675
R55214 VCC.n9354 VCC.n8919 0.00675
R55215 VCC.n9366 VCC.n8916 0.00675
R55216 VCC.n9372 VCC.n8894 0.00675
R55217 VCC.n8900 VCC.n8899 0.00675
R55218 VCC.n9393 VCC.n8892 0.00675
R55219 VCC.n9224 VCC.n9223 0.00675
R55220 VCC.n9239 VCC.n8976 0.00675
R55221 VCC.n9275 VCC.n9273 0.00675
R55222 VCC.n9306 VCC.n8949 0.00675
R55223 VCC.n9187 VCC.n8999 0.00675
R55224 VCC.n9217 VCC.n8985 0.00675
R55225 VCC.n9225 VCC.n9221 0.00675
R55226 VCC.n9278 VCC.n8960 0.00675
R55227 VCC.n9274 VCC.n8958 0.00675
R55228 VCC.n9076 VCC.n9069 0.00675
R55229 VCC.n9119 VCC.n9043 0.00675
R55230 VCC.n9150 VCC.n9149 0.00675
R55231 VCC.n9171 VCC.n9011 0.00675
R55232 VCC.n9112 VCC.n9048 0.00675
R55233 VCC.n9118 VCC.n9044 0.00675
R55234 VCC.n9148 VCC.n9022 0.00675
R55235 VCC.n9156 VCC.n9005 0.00675
R55236 VCC.n9185 VCC.n9001 0.00675
R55237 VCC.n9627 VCC.n9620 0.00675
R55238 VCC.n9670 VCC.n9594 0.00675
R55239 VCC.n9701 VCC.n9700 0.00675
R55240 VCC.n9722 VCC.n9562 0.00675
R55241 VCC.n9663 VCC.n9599 0.00675
R55242 VCC.n9669 VCC.n9595 0.00675
R55243 VCC.n9699 VCC.n9573 0.00675
R55244 VCC.n9707 VCC.n9556 0.00675
R55245 VCC.n9736 VCC.n9552 0.00675
R55246 VCC.n9776 VCC.n9775 0.00675
R55247 VCC.n9791 VCC.n9528 0.00675
R55248 VCC.n9827 VCC.n9825 0.00675
R55249 VCC.n9857 VCC.n9501 0.00675
R55250 VCC.n9738 VCC.n9550 0.00675
R55251 VCC.n9769 VCC.n9537 0.00675
R55252 VCC.n9777 VCC.n9773 0.00675
R55253 VCC.n9830 VCC.n9512 0.00675
R55254 VCC.n9826 VCC.n9510 0.00675
R55255 VCC.n9477 VCC.n9468 0.00675
R55256 VCC.n9471 VCC.n9469 0.00675
R55257 VCC.n9945 VCC.n9451 0.00675
R55258 VCC.n9475 VCC.n9470 0.00675
R55259 VCC.n9910 VCC.n9472 0.00675
R55260 VCC.n9458 VCC.n9455 0.00675
R55261 VCC.n9944 VCC.n9943 0.00675
R55262 VCC.n9942 VCC.n9938 0.00675
R55263 VCC.n10463 VCC.n10029 0.00675
R55264 VCC.n10475 VCC.n10023 0.00675
R55265 VCC.n10009 VCC.n10005 0.00675
R55266 VCC.n10462 VCC.n10027 0.00675
R55267 VCC.n10474 VCC.n10024 0.00675
R55268 VCC.n10480 VCC.n10002 0.00675
R55269 VCC.n10008 VCC.n10007 0.00675
R55270 VCC.n10501 VCC.n10000 0.00675
R55271 VCC.n10332 VCC.n10331 0.00675
R55272 VCC.n10347 VCC.n10084 0.00675
R55273 VCC.n10383 VCC.n10381 0.00675
R55274 VCC.n10414 VCC.n10057 0.00675
R55275 VCC.n10295 VCC.n10107 0.00675
R55276 VCC.n10325 VCC.n10093 0.00675
R55277 VCC.n10333 VCC.n10329 0.00675
R55278 VCC.n10386 VCC.n10068 0.00675
R55279 VCC.n10382 VCC.n10066 0.00675
R55280 VCC.n10184 VCC.n10177 0.00675
R55281 VCC.n10227 VCC.n10151 0.00675
R55282 VCC.n10258 VCC.n10257 0.00675
R55283 VCC.n10279 VCC.n10119 0.00675
R55284 VCC.n10220 VCC.n10156 0.00675
R55285 VCC.n10226 VCC.n10152 0.00675
R55286 VCC.n10256 VCC.n10130 0.00675
R55287 VCC.n10264 VCC.n10113 0.00675
R55288 VCC.n10293 VCC.n10109 0.00675
R55289 VCC.n10734 VCC.n10727 0.00675
R55290 VCC.n10777 VCC.n10701 0.00675
R55291 VCC.n10808 VCC.n10807 0.00675
R55292 VCC.n10829 VCC.n10669 0.00675
R55293 VCC.n10770 VCC.n10706 0.00675
R55294 VCC.n10776 VCC.n10702 0.00675
R55295 VCC.n10806 VCC.n10680 0.00675
R55296 VCC.n10814 VCC.n10663 0.00675
R55297 VCC.n10843 VCC.n10659 0.00675
R55298 VCC.n10883 VCC.n10882 0.00675
R55299 VCC.n10898 VCC.n10635 0.00675
R55300 VCC.n10934 VCC.n10932 0.00675
R55301 VCC.n10964 VCC.n10608 0.00675
R55302 VCC.n10845 VCC.n10657 0.00675
R55303 VCC.n10876 VCC.n10644 0.00675
R55304 VCC.n10884 VCC.n10880 0.00675
R55305 VCC.n10937 VCC.n10619 0.00675
R55306 VCC.n10933 VCC.n10617 0.00675
R55307 VCC.n10584 VCC.n10575 0.00675
R55308 VCC.n10578 VCC.n10576 0.00675
R55309 VCC.n11052 VCC.n10558 0.00675
R55310 VCC.n10582 VCC.n10577 0.00675
R55311 VCC.n11017 VCC.n10579 0.00675
R55312 VCC.n10565 VCC.n10562 0.00675
R55313 VCC.n11051 VCC.n11050 0.00675
R55314 VCC.n11049 VCC.n11045 0.00675
R55315 VCC.n11570 VCC.n11136 0.00675
R55316 VCC.n11582 VCC.n11130 0.00675
R55317 VCC.n11116 VCC.n11112 0.00675
R55318 VCC.n11569 VCC.n11134 0.00675
R55319 VCC.n11581 VCC.n11131 0.00675
R55320 VCC.n11587 VCC.n11109 0.00675
R55321 VCC.n11115 VCC.n11114 0.00675
R55322 VCC.n11608 VCC.n11107 0.00675
R55323 VCC.n11439 VCC.n11438 0.00675
R55324 VCC.n11454 VCC.n11191 0.00675
R55325 VCC.n11490 VCC.n11488 0.00675
R55326 VCC.n11521 VCC.n11164 0.00675
R55327 VCC.n11402 VCC.n11214 0.00675
R55328 VCC.n11432 VCC.n11200 0.00675
R55329 VCC.n11440 VCC.n11436 0.00675
R55330 VCC.n11493 VCC.n11175 0.00675
R55331 VCC.n11489 VCC.n11173 0.00675
R55332 VCC.n11291 VCC.n11284 0.00675
R55333 VCC.n11334 VCC.n11258 0.00675
R55334 VCC.n11365 VCC.n11364 0.00675
R55335 VCC.n11386 VCC.n11226 0.00675
R55336 VCC.n11327 VCC.n11263 0.00675
R55337 VCC.n11333 VCC.n11259 0.00675
R55338 VCC.n11363 VCC.n11237 0.00675
R55339 VCC.n11371 VCC.n11220 0.00675
R55340 VCC.n11400 VCC.n11216 0.00675
R55341 VCC.n11841 VCC.n11834 0.00675
R55342 VCC.n11884 VCC.n11808 0.00675
R55343 VCC.n11915 VCC.n11914 0.00675
R55344 VCC.n11936 VCC.n11776 0.00675
R55345 VCC.n11877 VCC.n11813 0.00675
R55346 VCC.n11883 VCC.n11809 0.00675
R55347 VCC.n11913 VCC.n11787 0.00675
R55348 VCC.n11921 VCC.n11770 0.00675
R55349 VCC.n11950 VCC.n11766 0.00675
R55350 VCC.n11990 VCC.n11989 0.00675
R55351 VCC.n12005 VCC.n11742 0.00675
R55352 VCC.n12041 VCC.n12039 0.00675
R55353 VCC.n12071 VCC.n11715 0.00675
R55354 VCC.n11952 VCC.n11764 0.00675
R55355 VCC.n11983 VCC.n11751 0.00675
R55356 VCC.n11991 VCC.n11987 0.00675
R55357 VCC.n12044 VCC.n11726 0.00675
R55358 VCC.n12040 VCC.n11724 0.00675
R55359 VCC.n11691 VCC.n11682 0.00675
R55360 VCC.n11685 VCC.n11683 0.00675
R55361 VCC.n12159 VCC.n11665 0.00675
R55362 VCC.n11689 VCC.n11684 0.00675
R55363 VCC.n12124 VCC.n11686 0.00675
R55364 VCC.n11672 VCC.n11669 0.00675
R55365 VCC.n12158 VCC.n12157 0.00675
R55366 VCC.n12156 VCC.n12152 0.00675
R55367 VCC.n12677 VCC.n12243 0.00675
R55368 VCC.n12689 VCC.n12237 0.00675
R55369 VCC.n12223 VCC.n12219 0.00675
R55370 VCC.n12676 VCC.n12241 0.00675
R55371 VCC.n12688 VCC.n12238 0.00675
R55372 VCC.n12694 VCC.n12216 0.00675
R55373 VCC.n12222 VCC.n12221 0.00675
R55374 VCC.n12715 VCC.n12214 0.00675
R55375 VCC.n12546 VCC.n12545 0.00675
R55376 VCC.n12561 VCC.n12298 0.00675
R55377 VCC.n12597 VCC.n12595 0.00675
R55378 VCC.n12628 VCC.n12271 0.00675
R55379 VCC.n12509 VCC.n12321 0.00675
R55380 VCC.n12539 VCC.n12307 0.00675
R55381 VCC.n12547 VCC.n12543 0.00675
R55382 VCC.n12600 VCC.n12282 0.00675
R55383 VCC.n12596 VCC.n12280 0.00675
R55384 VCC.n12398 VCC.n12391 0.00675
R55385 VCC.n12441 VCC.n12365 0.00675
R55386 VCC.n12472 VCC.n12471 0.00675
R55387 VCC.n12493 VCC.n12333 0.00675
R55388 VCC.n12434 VCC.n12370 0.00675
R55389 VCC.n12440 VCC.n12366 0.00675
R55390 VCC.n12470 VCC.n12344 0.00675
R55391 VCC.n12478 VCC.n12327 0.00675
R55392 VCC.n12507 VCC.n12323 0.00675
R55393 VCC.n12948 VCC.n12941 0.00675
R55394 VCC.n12991 VCC.n12915 0.00675
R55395 VCC.n13022 VCC.n13021 0.00675
R55396 VCC.n13043 VCC.n12883 0.00675
R55397 VCC.n12984 VCC.n12920 0.00675
R55398 VCC.n12990 VCC.n12916 0.00675
R55399 VCC.n13020 VCC.n12894 0.00675
R55400 VCC.n13028 VCC.n12877 0.00675
R55401 VCC.n13057 VCC.n12873 0.00675
R55402 VCC.n13097 VCC.n13096 0.00675
R55403 VCC.n13112 VCC.n12849 0.00675
R55404 VCC.n13148 VCC.n13146 0.00675
R55405 VCC.n13178 VCC.n12822 0.00675
R55406 VCC.n13059 VCC.n12871 0.00675
R55407 VCC.n13090 VCC.n12858 0.00675
R55408 VCC.n13098 VCC.n13094 0.00675
R55409 VCC.n13151 VCC.n12833 0.00675
R55410 VCC.n13147 VCC.n12831 0.00675
R55411 VCC.n12798 VCC.n12789 0.00675
R55412 VCC.n12792 VCC.n12790 0.00675
R55413 VCC.n13266 VCC.n12772 0.00675
R55414 VCC.n12796 VCC.n12791 0.00675
R55415 VCC.n13231 VCC.n12793 0.00675
R55416 VCC.n12779 VCC.n12776 0.00675
R55417 VCC.n13265 VCC.n13264 0.00675
R55418 VCC.n13263 VCC.n13259 0.00675
R55419 VCC.n13784 VCC.n13350 0.00675
R55420 VCC.n13796 VCC.n13344 0.00675
R55421 VCC.n13330 VCC.n13326 0.00675
R55422 VCC.n13783 VCC.n13348 0.00675
R55423 VCC.n13795 VCC.n13345 0.00675
R55424 VCC.n13801 VCC.n13323 0.00675
R55425 VCC.n13329 VCC.n13328 0.00675
R55426 VCC.n13822 VCC.n13321 0.00675
R55427 VCC.n13653 VCC.n13652 0.00675
R55428 VCC.n13668 VCC.n13405 0.00675
R55429 VCC.n13704 VCC.n13702 0.00675
R55430 VCC.n13735 VCC.n13378 0.00675
R55431 VCC.n13616 VCC.n13428 0.00675
R55432 VCC.n13646 VCC.n13414 0.00675
R55433 VCC.n13654 VCC.n13650 0.00675
R55434 VCC.n13707 VCC.n13389 0.00675
R55435 VCC.n13703 VCC.n13387 0.00675
R55436 VCC.n13505 VCC.n13498 0.00675
R55437 VCC.n13548 VCC.n13472 0.00675
R55438 VCC.n13579 VCC.n13578 0.00675
R55439 VCC.n13600 VCC.n13440 0.00675
R55440 VCC.n13541 VCC.n13477 0.00675
R55441 VCC.n13547 VCC.n13473 0.00675
R55442 VCC.n13577 VCC.n13451 0.00675
R55443 VCC.n13585 VCC.n13434 0.00675
R55444 VCC.n13614 VCC.n13430 0.00675
R55445 VCC.n14055 VCC.n14048 0.00675
R55446 VCC.n14098 VCC.n14022 0.00675
R55447 VCC.n14129 VCC.n14128 0.00675
R55448 VCC.n14150 VCC.n13990 0.00675
R55449 VCC.n14091 VCC.n14027 0.00675
R55450 VCC.n14097 VCC.n14023 0.00675
R55451 VCC.n14127 VCC.n14001 0.00675
R55452 VCC.n14135 VCC.n13984 0.00675
R55453 VCC.n14164 VCC.n13980 0.00675
R55454 VCC.n14204 VCC.n14203 0.00675
R55455 VCC.n14219 VCC.n13956 0.00675
R55456 VCC.n14255 VCC.n14253 0.00675
R55457 VCC.n14285 VCC.n13929 0.00675
R55458 VCC.n14166 VCC.n13978 0.00675
R55459 VCC.n14197 VCC.n13965 0.00675
R55460 VCC.n14205 VCC.n14201 0.00675
R55461 VCC.n14258 VCC.n13940 0.00675
R55462 VCC.n14254 VCC.n13938 0.00675
R55463 VCC.n13905 VCC.n13896 0.00675
R55464 VCC.n13899 VCC.n13897 0.00675
R55465 VCC.n14373 VCC.n13879 0.00675
R55466 VCC.n13903 VCC.n13898 0.00675
R55467 VCC.n14338 VCC.n13900 0.00675
R55468 VCC.n13886 VCC.n13883 0.00675
R55469 VCC.n14372 VCC.n14371 0.00675
R55470 VCC.n14370 VCC.n14366 0.00675
R55471 VCC.n14891 VCC.n14457 0.00675
R55472 VCC.n14903 VCC.n14451 0.00675
R55473 VCC.n14437 VCC.n14433 0.00675
R55474 VCC.n14890 VCC.n14455 0.00675
R55475 VCC.n14902 VCC.n14452 0.00675
R55476 VCC.n14908 VCC.n14430 0.00675
R55477 VCC.n14436 VCC.n14435 0.00675
R55478 VCC.n14929 VCC.n14428 0.00675
R55479 VCC.n14760 VCC.n14759 0.00675
R55480 VCC.n14775 VCC.n14512 0.00675
R55481 VCC.n14811 VCC.n14809 0.00675
R55482 VCC.n14842 VCC.n14485 0.00675
R55483 VCC.n14723 VCC.n14535 0.00675
R55484 VCC.n14753 VCC.n14521 0.00675
R55485 VCC.n14761 VCC.n14757 0.00675
R55486 VCC.n14814 VCC.n14496 0.00675
R55487 VCC.n14810 VCC.n14494 0.00675
R55488 VCC.n14612 VCC.n14605 0.00675
R55489 VCC.n14655 VCC.n14579 0.00675
R55490 VCC.n14686 VCC.n14685 0.00675
R55491 VCC.n14707 VCC.n14547 0.00675
R55492 VCC.n14648 VCC.n14584 0.00675
R55493 VCC.n14654 VCC.n14580 0.00675
R55494 VCC.n14684 VCC.n14558 0.00675
R55495 VCC.n14692 VCC.n14541 0.00675
R55496 VCC.n14721 VCC.n14537 0.00675
R55497 VCC.n15162 VCC.n15155 0.00675
R55498 VCC.n15205 VCC.n15129 0.00675
R55499 VCC.n15236 VCC.n15235 0.00675
R55500 VCC.n15257 VCC.n15097 0.00675
R55501 VCC.n15198 VCC.n15134 0.00675
R55502 VCC.n15204 VCC.n15130 0.00675
R55503 VCC.n15234 VCC.n15108 0.00675
R55504 VCC.n15242 VCC.n15091 0.00675
R55505 VCC.n15271 VCC.n15087 0.00675
R55506 VCC.n15311 VCC.n15310 0.00675
R55507 VCC.n15326 VCC.n15063 0.00675
R55508 VCC.n15362 VCC.n15360 0.00675
R55509 VCC.n15392 VCC.n15036 0.00675
R55510 VCC.n15273 VCC.n15085 0.00675
R55511 VCC.n15304 VCC.n15072 0.00675
R55512 VCC.n15312 VCC.n15308 0.00675
R55513 VCC.n15365 VCC.n15047 0.00675
R55514 VCC.n15361 VCC.n15045 0.00675
R55515 VCC.n15012 VCC.n15003 0.00675
R55516 VCC.n15006 VCC.n15004 0.00675
R55517 VCC.n15480 VCC.n14986 0.00675
R55518 VCC.n15010 VCC.n15005 0.00675
R55519 VCC.n15445 VCC.n15007 0.00675
R55520 VCC.n14993 VCC.n14990 0.00675
R55521 VCC.n15479 VCC.n15478 0.00675
R55522 VCC.n15477 VCC.n15473 0.00675
R55523 VCC.n15998 VCC.n15564 0.00675
R55524 VCC.n16010 VCC.n15558 0.00675
R55525 VCC.n15544 VCC.n15540 0.00675
R55526 VCC.n15997 VCC.n15562 0.00675
R55527 VCC.n16009 VCC.n15559 0.00675
R55528 VCC.n16015 VCC.n15537 0.00675
R55529 VCC.n15543 VCC.n15542 0.00675
R55530 VCC.n16036 VCC.n15535 0.00675
R55531 VCC.n15867 VCC.n15866 0.00675
R55532 VCC.n15882 VCC.n15619 0.00675
R55533 VCC.n15918 VCC.n15916 0.00675
R55534 VCC.n15949 VCC.n15592 0.00675
R55535 VCC.n15830 VCC.n15642 0.00675
R55536 VCC.n15860 VCC.n15628 0.00675
R55537 VCC.n15868 VCC.n15864 0.00675
R55538 VCC.n15921 VCC.n15603 0.00675
R55539 VCC.n15917 VCC.n15601 0.00675
R55540 VCC.n15719 VCC.n15712 0.00675
R55541 VCC.n15762 VCC.n15686 0.00675
R55542 VCC.n15793 VCC.n15792 0.00675
R55543 VCC.n15814 VCC.n15654 0.00675
R55544 VCC.n15755 VCC.n15691 0.00675
R55545 VCC.n15761 VCC.n15687 0.00675
R55546 VCC.n15791 VCC.n15665 0.00675
R55547 VCC.n15799 VCC.n15648 0.00675
R55548 VCC.n15828 VCC.n15644 0.00675
R55549 VCC.n16269 VCC.n16262 0.00675
R55550 VCC.n16312 VCC.n16236 0.00675
R55551 VCC.n16343 VCC.n16342 0.00675
R55552 VCC.n16364 VCC.n16204 0.00675
R55553 VCC.n16305 VCC.n16241 0.00675
R55554 VCC.n16311 VCC.n16237 0.00675
R55555 VCC.n16341 VCC.n16215 0.00675
R55556 VCC.n16349 VCC.n16198 0.00675
R55557 VCC.n16378 VCC.n16194 0.00675
R55558 VCC.n16418 VCC.n16417 0.00675
R55559 VCC.n16433 VCC.n16170 0.00675
R55560 VCC.n16469 VCC.n16467 0.00675
R55561 VCC.n16499 VCC.n16143 0.00675
R55562 VCC.n16380 VCC.n16192 0.00675
R55563 VCC.n16411 VCC.n16179 0.00675
R55564 VCC.n16419 VCC.n16415 0.00675
R55565 VCC.n16472 VCC.n16154 0.00675
R55566 VCC.n16468 VCC.n16152 0.00675
R55567 VCC.n16119 VCC.n16110 0.00675
R55568 VCC.n16113 VCC.n16111 0.00675
R55569 VCC.n16587 VCC.n16093 0.00675
R55570 VCC.n16117 VCC.n16112 0.00675
R55571 VCC.n16552 VCC.n16114 0.00675
R55572 VCC.n16100 VCC.n16097 0.00675
R55573 VCC.n16586 VCC.n16585 0.00675
R55574 VCC.n16584 VCC.n16580 0.00675
R55575 VCC.n17105 VCC.n16671 0.00675
R55576 VCC.n17117 VCC.n16665 0.00675
R55577 VCC.n16651 VCC.n16647 0.00675
R55578 VCC.n17104 VCC.n16669 0.00675
R55579 VCC.n17116 VCC.n16666 0.00675
R55580 VCC.n17122 VCC.n16644 0.00675
R55581 VCC.n16650 VCC.n16649 0.00675
R55582 VCC.n17143 VCC.n16642 0.00675
R55583 VCC.n16974 VCC.n16973 0.00675
R55584 VCC.n16989 VCC.n16726 0.00675
R55585 VCC.n17025 VCC.n17023 0.00675
R55586 VCC.n17056 VCC.n16699 0.00675
R55587 VCC.n16937 VCC.n16749 0.00675
R55588 VCC.n16967 VCC.n16735 0.00675
R55589 VCC.n16975 VCC.n16971 0.00675
R55590 VCC.n17028 VCC.n16710 0.00675
R55591 VCC.n17024 VCC.n16708 0.00675
R55592 VCC.n16826 VCC.n16819 0.00675
R55593 VCC.n16869 VCC.n16793 0.00675
R55594 VCC.n16900 VCC.n16899 0.00675
R55595 VCC.n16921 VCC.n16761 0.00675
R55596 VCC.n16862 VCC.n16798 0.00675
R55597 VCC.n16868 VCC.n16794 0.00675
R55598 VCC.n16898 VCC.n16772 0.00675
R55599 VCC.n16906 VCC.n16755 0.00675
R55600 VCC.n16935 VCC.n16751 0.00675
R55601 VCC.n17338 VCC.n17337 0.00675
R55602 VCC.n17353 VCC.n17277 0.00675
R55603 VCC.n17389 VCC.n17387 0.00675
R55604 VCC.n17419 VCC.n17250 0.00675
R55605 VCC.n17300 VCC.n17299 0.00675
R55606 VCC.n17331 VCC.n17286 0.00675
R55607 VCC.n17339 VCC.n17335 0.00675
R55608 VCC.n17392 VCC.n17261 0.00675
R55609 VCC.n17388 VCC.n17259 0.00675
R55610 VCC.n17226 VCC.n17217 0.00675
R55611 VCC.n17220 VCC.n17218 0.00675
R55612 VCC.n17507 VCC.n17200 0.00675
R55613 VCC.n17224 VCC.n17219 0.00675
R55614 VCC.n17472 VCC.n17221 0.00675
R55615 VCC.n17207 VCC.n17204 0.00675
R55616 VCC.n17506 VCC.n17505 0.00675
R55617 VCC.n17504 VCC.n17500 0.00675
R55618 VCC.n206 VCC.n196 0.00585714
R55619 VCC.n238 VCC.n237 0.00585714
R55620 VCC.n158 VCC.n150 0.00585714
R55621 VCC.n187 VCC.n174 0.00585714
R55622 VCC.n245 VCC.n244 0.00585714
R55623 VCC.n331 VCC.n320 0.00585714
R55624 VCC.n328 VCC.n320 0.00585714
R55625 VCC.n355 VCC.n112 0.00585714
R55626 VCC.n390 VCC.n90 0.00585714
R55627 VCC.n434 VCC.n433 0.00585714
R55628 VCC.n373 VCC.n88 0.00585714
R55629 VCC.n410 VCC.n71 0.00585714
R55630 VCC.n452 VCC.n58 0.00585714
R55631 VCC.n489 VCC.n488 0.00585714
R55632 VCC.n510 VCC.n509 0.00585714
R55633 VCC.n522 VCC.n26 0.00585714
R55634 VCC.n17 VCC.n8 0.00585714
R55635 VCC.n11 VCC.n9 0.00585714
R55636 VCC.n61 VCC.n50 0.00585714
R55637 VCC.n483 VCC.n48 0.00585714
R55638 VCC.n511 VCC.n31 0.00585714
R55639 VCC.n758 VCC.n748 0.00585714
R55640 VCC.n790 VCC.n789 0.00585714
R55641 VCC.n710 VCC.n702 0.00585714
R55642 VCC.n739 VCC.n726 0.00585714
R55643 VCC.n797 VCC.n796 0.00585714
R55644 VCC.n883 VCC.n872 0.00585714
R55645 VCC.n880 VCC.n872 0.00585714
R55646 VCC.n907 VCC.n664 0.00585714
R55647 VCC.n942 VCC.n642 0.00585714
R55648 VCC.n986 VCC.n985 0.00585714
R55649 VCC.n925 VCC.n640 0.00585714
R55650 VCC.n962 VCC.n623 0.00585714
R55651 VCC.n1004 VCC.n610 0.00585714
R55652 VCC.n1041 VCC.n1040 0.00585714
R55653 VCC.n1062 VCC.n1061 0.00585714
R55654 VCC.n1074 VCC.n578 0.00585714
R55655 VCC.n569 VCC.n562 0.00585714
R55656 VCC.n1091 VCC.n563 0.00585714
R55657 VCC.n613 VCC.n602 0.00585714
R55658 VCC.n1035 VCC.n600 0.00585714
R55659 VCC.n1063 VCC.n583 0.00585714
R55660 VCC.n1562 VCC.n1166 0.00585714
R55661 VCC.n1589 VCC.n1588 0.00585714
R55662 VCC.n1626 VCC.n1133 0.00585714
R55663 VCC.n1625 VCC.n1624 0.00585714
R55664 VCC.n1122 VCC.n1119 0.00585714
R55665 VCC.n1641 VCC.n1640 0.00585714
R55666 VCC.n1170 VCC.n1155 0.00585714
R55667 VCC.n1603 VCC.n1602 0.00585714
R55668 VCC.n1627 VCC.n1131 0.00585714
R55669 VCC.n1430 VCC.n1235 0.00585714
R55670 VCC.n1437 VCC.n1430 0.00585714
R55671 VCC.n1464 VCC.n1221 0.00585714
R55672 VCC.n1499 VCC.n1199 0.00585714
R55673 VCC.n1544 VCC.n1543 0.00585714
R55674 VCC.n1482 VCC.n1197 0.00585714
R55675 VCC.n1519 VCC.n1180 0.00585714
R55676 VCC.n1316 VCC.n1306 0.00585714
R55677 VCC.n1348 VCC.n1347 0.00585714
R55678 VCC.n1268 VCC.n1260 0.00585714
R55679 VCC.n1297 VCC.n1284 0.00585714
R55680 VCC.n1355 VCC.n1354 0.00585714
R55681 VCC.n1867 VCC.n1857 0.00585714
R55682 VCC.n1899 VCC.n1898 0.00585714
R55683 VCC.n1819 VCC.n1811 0.00585714
R55684 VCC.n1848 VCC.n1835 0.00585714
R55685 VCC.n1906 VCC.n1905 0.00585714
R55686 VCC.n1992 VCC.n1981 0.00585714
R55687 VCC.n1989 VCC.n1981 0.00585714
R55688 VCC.n2016 VCC.n1773 0.00585714
R55689 VCC.n2051 VCC.n1751 0.00585714
R55690 VCC.n2095 VCC.n2094 0.00585714
R55691 VCC.n2034 VCC.n1749 0.00585714
R55692 VCC.n2071 VCC.n1732 0.00585714
R55693 VCC.n2113 VCC.n1719 0.00585714
R55694 VCC.n2150 VCC.n2149 0.00585714
R55695 VCC.n2171 VCC.n2170 0.00585714
R55696 VCC.n2183 VCC.n1687 0.00585714
R55697 VCC.n1678 VCC.n1671 0.00585714
R55698 VCC.n2200 VCC.n1672 0.00585714
R55699 VCC.n1722 VCC.n1711 0.00585714
R55700 VCC.n2144 VCC.n1709 0.00585714
R55701 VCC.n2172 VCC.n1692 0.00585714
R55702 VCC.n2671 VCC.n2275 0.00585714
R55703 VCC.n2698 VCC.n2697 0.00585714
R55704 VCC.n2735 VCC.n2242 0.00585714
R55705 VCC.n2734 VCC.n2733 0.00585714
R55706 VCC.n2231 VCC.n2228 0.00585714
R55707 VCC.n2750 VCC.n2749 0.00585714
R55708 VCC.n2279 VCC.n2264 0.00585714
R55709 VCC.n2712 VCC.n2711 0.00585714
R55710 VCC.n2736 VCC.n2240 0.00585714
R55711 VCC.n2539 VCC.n2344 0.00585714
R55712 VCC.n2546 VCC.n2539 0.00585714
R55713 VCC.n2573 VCC.n2330 0.00585714
R55714 VCC.n2608 VCC.n2308 0.00585714
R55715 VCC.n2653 VCC.n2652 0.00585714
R55716 VCC.n2591 VCC.n2306 0.00585714
R55717 VCC.n2628 VCC.n2289 0.00585714
R55718 VCC.n2425 VCC.n2415 0.00585714
R55719 VCC.n2457 VCC.n2456 0.00585714
R55720 VCC.n2377 VCC.n2369 0.00585714
R55721 VCC.n2406 VCC.n2393 0.00585714
R55722 VCC.n2464 VCC.n2463 0.00585714
R55723 VCC.n2976 VCC.n2966 0.00585714
R55724 VCC.n3008 VCC.n3007 0.00585714
R55725 VCC.n2928 VCC.n2920 0.00585714
R55726 VCC.n2957 VCC.n2944 0.00585714
R55727 VCC.n3015 VCC.n3014 0.00585714
R55728 VCC.n3101 VCC.n3090 0.00585714
R55729 VCC.n3098 VCC.n3090 0.00585714
R55730 VCC.n3125 VCC.n2882 0.00585714
R55731 VCC.n3160 VCC.n2860 0.00585714
R55732 VCC.n3204 VCC.n3203 0.00585714
R55733 VCC.n3143 VCC.n2858 0.00585714
R55734 VCC.n3180 VCC.n2841 0.00585714
R55735 VCC.n3222 VCC.n2828 0.00585714
R55736 VCC.n3259 VCC.n3258 0.00585714
R55737 VCC.n3280 VCC.n3279 0.00585714
R55738 VCC.n3292 VCC.n2796 0.00585714
R55739 VCC.n2787 VCC.n2780 0.00585714
R55740 VCC.n3309 VCC.n2781 0.00585714
R55741 VCC.n2831 VCC.n2820 0.00585714
R55742 VCC.n3253 VCC.n2818 0.00585714
R55743 VCC.n3281 VCC.n2801 0.00585714
R55744 VCC.n3780 VCC.n3384 0.00585714
R55745 VCC.n3807 VCC.n3806 0.00585714
R55746 VCC.n3844 VCC.n3351 0.00585714
R55747 VCC.n3843 VCC.n3842 0.00585714
R55748 VCC.n3340 VCC.n3337 0.00585714
R55749 VCC.n3859 VCC.n3858 0.00585714
R55750 VCC.n3388 VCC.n3373 0.00585714
R55751 VCC.n3821 VCC.n3820 0.00585714
R55752 VCC.n3845 VCC.n3349 0.00585714
R55753 VCC.n3648 VCC.n3453 0.00585714
R55754 VCC.n3655 VCC.n3648 0.00585714
R55755 VCC.n3682 VCC.n3439 0.00585714
R55756 VCC.n3717 VCC.n3417 0.00585714
R55757 VCC.n3762 VCC.n3761 0.00585714
R55758 VCC.n3700 VCC.n3415 0.00585714
R55759 VCC.n3737 VCC.n3398 0.00585714
R55760 VCC.n3534 VCC.n3524 0.00585714
R55761 VCC.n3566 VCC.n3565 0.00585714
R55762 VCC.n3486 VCC.n3478 0.00585714
R55763 VCC.n3515 VCC.n3502 0.00585714
R55764 VCC.n3573 VCC.n3572 0.00585714
R55765 VCC.n4085 VCC.n4075 0.00585714
R55766 VCC.n4117 VCC.n4116 0.00585714
R55767 VCC.n4037 VCC.n4029 0.00585714
R55768 VCC.n4066 VCC.n4053 0.00585714
R55769 VCC.n4124 VCC.n4123 0.00585714
R55770 VCC.n4210 VCC.n4199 0.00585714
R55771 VCC.n4207 VCC.n4199 0.00585714
R55772 VCC.n4234 VCC.n3991 0.00585714
R55773 VCC.n4269 VCC.n3969 0.00585714
R55774 VCC.n4313 VCC.n4312 0.00585714
R55775 VCC.n4252 VCC.n3967 0.00585714
R55776 VCC.n4289 VCC.n3950 0.00585714
R55777 VCC.n4331 VCC.n3937 0.00585714
R55778 VCC.n4368 VCC.n4367 0.00585714
R55779 VCC.n4389 VCC.n4388 0.00585714
R55780 VCC.n4401 VCC.n3905 0.00585714
R55781 VCC.n3896 VCC.n3889 0.00585714
R55782 VCC.n4418 VCC.n3890 0.00585714
R55783 VCC.n3940 VCC.n3929 0.00585714
R55784 VCC.n4362 VCC.n3927 0.00585714
R55785 VCC.n4390 VCC.n3910 0.00585714
R55786 VCC.n4889 VCC.n4493 0.00585714
R55787 VCC.n4916 VCC.n4915 0.00585714
R55788 VCC.n4953 VCC.n4460 0.00585714
R55789 VCC.n4952 VCC.n4951 0.00585714
R55790 VCC.n4449 VCC.n4446 0.00585714
R55791 VCC.n4968 VCC.n4967 0.00585714
R55792 VCC.n4497 VCC.n4482 0.00585714
R55793 VCC.n4930 VCC.n4929 0.00585714
R55794 VCC.n4954 VCC.n4458 0.00585714
R55795 VCC.n4757 VCC.n4562 0.00585714
R55796 VCC.n4764 VCC.n4757 0.00585714
R55797 VCC.n4791 VCC.n4548 0.00585714
R55798 VCC.n4826 VCC.n4526 0.00585714
R55799 VCC.n4871 VCC.n4870 0.00585714
R55800 VCC.n4809 VCC.n4524 0.00585714
R55801 VCC.n4846 VCC.n4507 0.00585714
R55802 VCC.n4643 VCC.n4633 0.00585714
R55803 VCC.n4675 VCC.n4674 0.00585714
R55804 VCC.n4595 VCC.n4587 0.00585714
R55805 VCC.n4624 VCC.n4611 0.00585714
R55806 VCC.n4682 VCC.n4681 0.00585714
R55807 VCC.n5194 VCC.n5184 0.00585714
R55808 VCC.n5226 VCC.n5225 0.00585714
R55809 VCC.n5146 VCC.n5138 0.00585714
R55810 VCC.n5175 VCC.n5162 0.00585714
R55811 VCC.n5233 VCC.n5232 0.00585714
R55812 VCC.n5319 VCC.n5308 0.00585714
R55813 VCC.n5316 VCC.n5308 0.00585714
R55814 VCC.n5343 VCC.n5100 0.00585714
R55815 VCC.n5378 VCC.n5078 0.00585714
R55816 VCC.n5422 VCC.n5421 0.00585714
R55817 VCC.n5361 VCC.n5076 0.00585714
R55818 VCC.n5398 VCC.n5059 0.00585714
R55819 VCC.n5440 VCC.n5046 0.00585714
R55820 VCC.n5477 VCC.n5476 0.00585714
R55821 VCC.n5498 VCC.n5497 0.00585714
R55822 VCC.n5510 VCC.n5014 0.00585714
R55823 VCC.n5005 VCC.n4998 0.00585714
R55824 VCC.n5527 VCC.n4999 0.00585714
R55825 VCC.n5049 VCC.n5038 0.00585714
R55826 VCC.n5471 VCC.n5036 0.00585714
R55827 VCC.n5499 VCC.n5019 0.00585714
R55828 VCC.n5998 VCC.n5602 0.00585714
R55829 VCC.n6025 VCC.n6024 0.00585714
R55830 VCC.n6062 VCC.n5569 0.00585714
R55831 VCC.n6061 VCC.n6060 0.00585714
R55832 VCC.n5558 VCC.n5555 0.00585714
R55833 VCC.n6077 VCC.n6076 0.00585714
R55834 VCC.n5606 VCC.n5591 0.00585714
R55835 VCC.n6039 VCC.n6038 0.00585714
R55836 VCC.n6063 VCC.n5567 0.00585714
R55837 VCC.n5866 VCC.n5671 0.00585714
R55838 VCC.n5873 VCC.n5866 0.00585714
R55839 VCC.n5900 VCC.n5657 0.00585714
R55840 VCC.n5935 VCC.n5635 0.00585714
R55841 VCC.n5980 VCC.n5979 0.00585714
R55842 VCC.n5918 VCC.n5633 0.00585714
R55843 VCC.n5955 VCC.n5616 0.00585714
R55844 VCC.n5752 VCC.n5742 0.00585714
R55845 VCC.n5784 VCC.n5783 0.00585714
R55846 VCC.n5704 VCC.n5696 0.00585714
R55847 VCC.n5733 VCC.n5720 0.00585714
R55848 VCC.n5791 VCC.n5790 0.00585714
R55849 VCC.n6303 VCC.n6293 0.00585714
R55850 VCC.n6335 VCC.n6334 0.00585714
R55851 VCC.n6255 VCC.n6247 0.00585714
R55852 VCC.n6284 VCC.n6271 0.00585714
R55853 VCC.n6342 VCC.n6341 0.00585714
R55854 VCC.n6428 VCC.n6417 0.00585714
R55855 VCC.n6425 VCC.n6417 0.00585714
R55856 VCC.n6452 VCC.n6209 0.00585714
R55857 VCC.n6487 VCC.n6187 0.00585714
R55858 VCC.n6531 VCC.n6530 0.00585714
R55859 VCC.n6470 VCC.n6185 0.00585714
R55860 VCC.n6507 VCC.n6168 0.00585714
R55861 VCC.n6549 VCC.n6155 0.00585714
R55862 VCC.n6586 VCC.n6585 0.00585714
R55863 VCC.n6607 VCC.n6606 0.00585714
R55864 VCC.n6619 VCC.n6123 0.00585714
R55865 VCC.n6114 VCC.n6107 0.00585714
R55866 VCC.n6636 VCC.n6108 0.00585714
R55867 VCC.n6158 VCC.n6147 0.00585714
R55868 VCC.n6580 VCC.n6145 0.00585714
R55869 VCC.n6608 VCC.n6128 0.00585714
R55870 VCC.n7107 VCC.n6711 0.00585714
R55871 VCC.n7134 VCC.n7133 0.00585714
R55872 VCC.n7171 VCC.n6678 0.00585714
R55873 VCC.n7170 VCC.n7169 0.00585714
R55874 VCC.n6667 VCC.n6664 0.00585714
R55875 VCC.n7186 VCC.n7185 0.00585714
R55876 VCC.n6715 VCC.n6700 0.00585714
R55877 VCC.n7148 VCC.n7147 0.00585714
R55878 VCC.n7172 VCC.n6676 0.00585714
R55879 VCC.n6975 VCC.n6780 0.00585714
R55880 VCC.n6982 VCC.n6975 0.00585714
R55881 VCC.n7009 VCC.n6766 0.00585714
R55882 VCC.n7044 VCC.n6744 0.00585714
R55883 VCC.n7089 VCC.n7088 0.00585714
R55884 VCC.n7027 VCC.n6742 0.00585714
R55885 VCC.n7064 VCC.n6725 0.00585714
R55886 VCC.n6861 VCC.n6851 0.00585714
R55887 VCC.n6893 VCC.n6892 0.00585714
R55888 VCC.n6813 VCC.n6805 0.00585714
R55889 VCC.n6842 VCC.n6829 0.00585714
R55890 VCC.n6900 VCC.n6899 0.00585714
R55891 VCC.n7412 VCC.n7402 0.00585714
R55892 VCC.n7444 VCC.n7443 0.00585714
R55893 VCC.n7364 VCC.n7356 0.00585714
R55894 VCC.n7393 VCC.n7380 0.00585714
R55895 VCC.n7451 VCC.n7450 0.00585714
R55896 VCC.n7537 VCC.n7526 0.00585714
R55897 VCC.n7534 VCC.n7526 0.00585714
R55898 VCC.n7561 VCC.n7318 0.00585714
R55899 VCC.n7596 VCC.n7296 0.00585714
R55900 VCC.n7640 VCC.n7639 0.00585714
R55901 VCC.n7579 VCC.n7294 0.00585714
R55902 VCC.n7616 VCC.n7277 0.00585714
R55903 VCC.n7658 VCC.n7264 0.00585714
R55904 VCC.n7695 VCC.n7694 0.00585714
R55905 VCC.n7716 VCC.n7715 0.00585714
R55906 VCC.n7728 VCC.n7232 0.00585714
R55907 VCC.n7223 VCC.n7216 0.00585714
R55908 VCC.n7745 VCC.n7217 0.00585714
R55909 VCC.n7267 VCC.n7256 0.00585714
R55910 VCC.n7689 VCC.n7254 0.00585714
R55911 VCC.n7717 VCC.n7237 0.00585714
R55912 VCC.n8216 VCC.n7820 0.00585714
R55913 VCC.n8243 VCC.n8242 0.00585714
R55914 VCC.n8280 VCC.n7787 0.00585714
R55915 VCC.n8279 VCC.n8278 0.00585714
R55916 VCC.n7776 VCC.n7773 0.00585714
R55917 VCC.n8295 VCC.n8294 0.00585714
R55918 VCC.n7824 VCC.n7809 0.00585714
R55919 VCC.n8257 VCC.n8256 0.00585714
R55920 VCC.n8281 VCC.n7785 0.00585714
R55921 VCC.n8084 VCC.n7889 0.00585714
R55922 VCC.n8091 VCC.n8084 0.00585714
R55923 VCC.n8118 VCC.n7875 0.00585714
R55924 VCC.n8153 VCC.n7853 0.00585714
R55925 VCC.n8198 VCC.n8197 0.00585714
R55926 VCC.n8136 VCC.n7851 0.00585714
R55927 VCC.n8173 VCC.n7834 0.00585714
R55928 VCC.n7970 VCC.n7960 0.00585714
R55929 VCC.n8002 VCC.n8001 0.00585714
R55930 VCC.n7922 VCC.n7914 0.00585714
R55931 VCC.n7951 VCC.n7938 0.00585714
R55932 VCC.n8009 VCC.n8008 0.00585714
R55933 VCC.n8646 VCC.n8635 0.00585714
R55934 VCC.n8643 VCC.n8635 0.00585714
R55935 VCC.n8670 VCC.n8427 0.00585714
R55936 VCC.n8705 VCC.n8405 0.00585714
R55937 VCC.n8749 VCC.n8748 0.00585714
R55938 VCC.n8688 VCC.n8403 0.00585714
R55939 VCC.n8725 VCC.n8386 0.00585714
R55940 VCC.n8767 VCC.n8373 0.00585714
R55941 VCC.n8804 VCC.n8803 0.00585714
R55942 VCC.n8825 VCC.n8824 0.00585714
R55943 VCC.n8837 VCC.n8341 0.00585714
R55944 VCC.n8332 VCC.n8325 0.00585714
R55945 VCC.n8854 VCC.n8326 0.00585714
R55946 VCC.n8376 VCC.n8365 0.00585714
R55947 VCC.n8798 VCC.n8363 0.00585714
R55948 VCC.n8826 VCC.n8346 0.00585714
R55949 VCC.n8521 VCC.n8511 0.00585714
R55950 VCC.n8553 VCC.n8552 0.00585714
R55951 VCC.n8473 VCC.n8465 0.00585714
R55952 VCC.n8502 VCC.n8489 0.00585714
R55953 VCC.n8560 VCC.n8559 0.00585714
R55954 VCC.n9325 VCC.n8929 0.00585714
R55955 VCC.n9352 VCC.n9351 0.00585714
R55956 VCC.n9389 VCC.n8896 0.00585714
R55957 VCC.n9388 VCC.n9387 0.00585714
R55958 VCC.n8885 VCC.n8882 0.00585714
R55959 VCC.n9404 VCC.n9403 0.00585714
R55960 VCC.n8933 VCC.n8918 0.00585714
R55961 VCC.n9366 VCC.n9365 0.00585714
R55962 VCC.n9390 VCC.n8894 0.00585714
R55963 VCC.n9193 VCC.n8998 0.00585714
R55964 VCC.n9200 VCC.n9193 0.00585714
R55965 VCC.n9227 VCC.n8984 0.00585714
R55966 VCC.n9262 VCC.n8962 0.00585714
R55967 VCC.n9307 VCC.n9306 0.00585714
R55968 VCC.n9245 VCC.n8960 0.00585714
R55969 VCC.n9282 VCC.n8943 0.00585714
R55970 VCC.n9079 VCC.n9069 0.00585714
R55971 VCC.n9111 VCC.n9110 0.00585714
R55972 VCC.n9031 VCC.n9023 0.00585714
R55973 VCC.n9060 VCC.n9047 0.00585714
R55974 VCC.n9118 VCC.n9117 0.00585714
R55975 VCC.n9630 VCC.n9620 0.00585714
R55976 VCC.n9662 VCC.n9661 0.00585714
R55977 VCC.n9582 VCC.n9574 0.00585714
R55978 VCC.n9611 VCC.n9598 0.00585714
R55979 VCC.n9669 VCC.n9668 0.00585714
R55980 VCC.n9755 VCC.n9744 0.00585714
R55981 VCC.n9752 VCC.n9744 0.00585714
R55982 VCC.n9779 VCC.n9536 0.00585714
R55983 VCC.n9814 VCC.n9514 0.00585714
R55984 VCC.n9858 VCC.n9857 0.00585714
R55985 VCC.n9797 VCC.n9512 0.00585714
R55986 VCC.n9834 VCC.n9495 0.00585714
R55987 VCC.n9876 VCC.n9482 0.00585714
R55988 VCC.n9913 VCC.n9912 0.00585714
R55989 VCC.n9934 VCC.n9933 0.00585714
R55990 VCC.n9946 VCC.n9450 0.00585714
R55991 VCC.n9441 VCC.n9434 0.00585714
R55992 VCC.n9963 VCC.n9435 0.00585714
R55993 VCC.n9485 VCC.n9474 0.00585714
R55994 VCC.n9907 VCC.n9472 0.00585714
R55995 VCC.n9935 VCC.n9455 0.00585714
R55996 VCC.n10433 VCC.n10037 0.00585714
R55997 VCC.n10460 VCC.n10459 0.00585714
R55998 VCC.n10497 VCC.n10004 0.00585714
R55999 VCC.n10496 VCC.n10495 0.00585714
R56000 VCC.n9993 VCC.n9990 0.00585714
R56001 VCC.n10512 VCC.n10511 0.00585714
R56002 VCC.n10041 VCC.n10026 0.00585714
R56003 VCC.n10474 VCC.n10473 0.00585714
R56004 VCC.n10498 VCC.n10002 0.00585714
R56005 VCC.n10301 VCC.n10106 0.00585714
R56006 VCC.n10308 VCC.n10301 0.00585714
R56007 VCC.n10335 VCC.n10092 0.00585714
R56008 VCC.n10370 VCC.n10070 0.00585714
R56009 VCC.n10415 VCC.n10414 0.00585714
R56010 VCC.n10353 VCC.n10068 0.00585714
R56011 VCC.n10390 VCC.n10051 0.00585714
R56012 VCC.n10187 VCC.n10177 0.00585714
R56013 VCC.n10219 VCC.n10218 0.00585714
R56014 VCC.n10139 VCC.n10131 0.00585714
R56015 VCC.n10168 VCC.n10155 0.00585714
R56016 VCC.n10226 VCC.n10225 0.00585714
R56017 VCC.n10737 VCC.n10727 0.00585714
R56018 VCC.n10769 VCC.n10768 0.00585714
R56019 VCC.n10689 VCC.n10681 0.00585714
R56020 VCC.n10718 VCC.n10705 0.00585714
R56021 VCC.n10776 VCC.n10775 0.00585714
R56022 VCC.n10862 VCC.n10851 0.00585714
R56023 VCC.n10859 VCC.n10851 0.00585714
R56024 VCC.n10886 VCC.n10643 0.00585714
R56025 VCC.n10921 VCC.n10621 0.00585714
R56026 VCC.n10965 VCC.n10964 0.00585714
R56027 VCC.n10904 VCC.n10619 0.00585714
R56028 VCC.n10941 VCC.n10602 0.00585714
R56029 VCC.n10983 VCC.n10589 0.00585714
R56030 VCC.n11020 VCC.n11019 0.00585714
R56031 VCC.n11041 VCC.n11040 0.00585714
R56032 VCC.n11053 VCC.n10557 0.00585714
R56033 VCC.n10548 VCC.n10541 0.00585714
R56034 VCC.n11070 VCC.n10542 0.00585714
R56035 VCC.n10592 VCC.n10581 0.00585714
R56036 VCC.n11014 VCC.n10579 0.00585714
R56037 VCC.n11042 VCC.n10562 0.00585714
R56038 VCC.n11540 VCC.n11144 0.00585714
R56039 VCC.n11567 VCC.n11566 0.00585714
R56040 VCC.n11604 VCC.n11111 0.00585714
R56041 VCC.n11603 VCC.n11602 0.00585714
R56042 VCC.n11100 VCC.n11097 0.00585714
R56043 VCC.n11619 VCC.n11618 0.00585714
R56044 VCC.n11148 VCC.n11133 0.00585714
R56045 VCC.n11581 VCC.n11580 0.00585714
R56046 VCC.n11605 VCC.n11109 0.00585714
R56047 VCC.n11408 VCC.n11213 0.00585714
R56048 VCC.n11415 VCC.n11408 0.00585714
R56049 VCC.n11442 VCC.n11199 0.00585714
R56050 VCC.n11477 VCC.n11177 0.00585714
R56051 VCC.n11522 VCC.n11521 0.00585714
R56052 VCC.n11460 VCC.n11175 0.00585714
R56053 VCC.n11497 VCC.n11158 0.00585714
R56054 VCC.n11294 VCC.n11284 0.00585714
R56055 VCC.n11326 VCC.n11325 0.00585714
R56056 VCC.n11246 VCC.n11238 0.00585714
R56057 VCC.n11275 VCC.n11262 0.00585714
R56058 VCC.n11333 VCC.n11332 0.00585714
R56059 VCC.n11844 VCC.n11834 0.00585714
R56060 VCC.n11876 VCC.n11875 0.00585714
R56061 VCC.n11796 VCC.n11788 0.00585714
R56062 VCC.n11825 VCC.n11812 0.00585714
R56063 VCC.n11883 VCC.n11882 0.00585714
R56064 VCC.n11969 VCC.n11958 0.00585714
R56065 VCC.n11966 VCC.n11958 0.00585714
R56066 VCC.n11993 VCC.n11750 0.00585714
R56067 VCC.n12028 VCC.n11728 0.00585714
R56068 VCC.n12072 VCC.n12071 0.00585714
R56069 VCC.n12011 VCC.n11726 0.00585714
R56070 VCC.n12048 VCC.n11709 0.00585714
R56071 VCC.n12090 VCC.n11696 0.00585714
R56072 VCC.n12127 VCC.n12126 0.00585714
R56073 VCC.n12148 VCC.n12147 0.00585714
R56074 VCC.n12160 VCC.n11664 0.00585714
R56075 VCC.n11655 VCC.n11648 0.00585714
R56076 VCC.n12177 VCC.n11649 0.00585714
R56077 VCC.n11699 VCC.n11688 0.00585714
R56078 VCC.n12121 VCC.n11686 0.00585714
R56079 VCC.n12149 VCC.n11669 0.00585714
R56080 VCC.n12647 VCC.n12251 0.00585714
R56081 VCC.n12674 VCC.n12673 0.00585714
R56082 VCC.n12711 VCC.n12218 0.00585714
R56083 VCC.n12710 VCC.n12709 0.00585714
R56084 VCC.n12207 VCC.n12204 0.00585714
R56085 VCC.n12726 VCC.n12725 0.00585714
R56086 VCC.n12255 VCC.n12240 0.00585714
R56087 VCC.n12688 VCC.n12687 0.00585714
R56088 VCC.n12712 VCC.n12216 0.00585714
R56089 VCC.n12515 VCC.n12320 0.00585714
R56090 VCC.n12522 VCC.n12515 0.00585714
R56091 VCC.n12549 VCC.n12306 0.00585714
R56092 VCC.n12584 VCC.n12284 0.00585714
R56093 VCC.n12629 VCC.n12628 0.00585714
R56094 VCC.n12567 VCC.n12282 0.00585714
R56095 VCC.n12604 VCC.n12265 0.00585714
R56096 VCC.n12401 VCC.n12391 0.00585714
R56097 VCC.n12433 VCC.n12432 0.00585714
R56098 VCC.n12353 VCC.n12345 0.00585714
R56099 VCC.n12382 VCC.n12369 0.00585714
R56100 VCC.n12440 VCC.n12439 0.00585714
R56101 VCC.n12951 VCC.n12941 0.00585714
R56102 VCC.n12983 VCC.n12982 0.00585714
R56103 VCC.n12903 VCC.n12895 0.00585714
R56104 VCC.n12932 VCC.n12919 0.00585714
R56105 VCC.n12990 VCC.n12989 0.00585714
R56106 VCC.n13076 VCC.n13065 0.00585714
R56107 VCC.n13073 VCC.n13065 0.00585714
R56108 VCC.n13100 VCC.n12857 0.00585714
R56109 VCC.n13135 VCC.n12835 0.00585714
R56110 VCC.n13179 VCC.n13178 0.00585714
R56111 VCC.n13118 VCC.n12833 0.00585714
R56112 VCC.n13155 VCC.n12816 0.00585714
R56113 VCC.n13197 VCC.n12803 0.00585714
R56114 VCC.n13234 VCC.n13233 0.00585714
R56115 VCC.n13255 VCC.n13254 0.00585714
R56116 VCC.n13267 VCC.n12771 0.00585714
R56117 VCC.n12762 VCC.n12755 0.00585714
R56118 VCC.n13284 VCC.n12756 0.00585714
R56119 VCC.n12806 VCC.n12795 0.00585714
R56120 VCC.n13228 VCC.n12793 0.00585714
R56121 VCC.n13256 VCC.n12776 0.00585714
R56122 VCC.n13754 VCC.n13358 0.00585714
R56123 VCC.n13781 VCC.n13780 0.00585714
R56124 VCC.n13818 VCC.n13325 0.00585714
R56125 VCC.n13817 VCC.n13816 0.00585714
R56126 VCC.n13314 VCC.n13311 0.00585714
R56127 VCC.n13833 VCC.n13832 0.00585714
R56128 VCC.n13362 VCC.n13347 0.00585714
R56129 VCC.n13795 VCC.n13794 0.00585714
R56130 VCC.n13819 VCC.n13323 0.00585714
R56131 VCC.n13622 VCC.n13427 0.00585714
R56132 VCC.n13629 VCC.n13622 0.00585714
R56133 VCC.n13656 VCC.n13413 0.00585714
R56134 VCC.n13691 VCC.n13391 0.00585714
R56135 VCC.n13736 VCC.n13735 0.00585714
R56136 VCC.n13674 VCC.n13389 0.00585714
R56137 VCC.n13711 VCC.n13372 0.00585714
R56138 VCC.n13508 VCC.n13498 0.00585714
R56139 VCC.n13540 VCC.n13539 0.00585714
R56140 VCC.n13460 VCC.n13452 0.00585714
R56141 VCC.n13489 VCC.n13476 0.00585714
R56142 VCC.n13547 VCC.n13546 0.00585714
R56143 VCC.n14058 VCC.n14048 0.00585714
R56144 VCC.n14090 VCC.n14089 0.00585714
R56145 VCC.n14010 VCC.n14002 0.00585714
R56146 VCC.n14039 VCC.n14026 0.00585714
R56147 VCC.n14097 VCC.n14096 0.00585714
R56148 VCC.n14183 VCC.n14172 0.00585714
R56149 VCC.n14180 VCC.n14172 0.00585714
R56150 VCC.n14207 VCC.n13964 0.00585714
R56151 VCC.n14242 VCC.n13942 0.00585714
R56152 VCC.n14286 VCC.n14285 0.00585714
R56153 VCC.n14225 VCC.n13940 0.00585714
R56154 VCC.n14262 VCC.n13923 0.00585714
R56155 VCC.n14304 VCC.n13910 0.00585714
R56156 VCC.n14341 VCC.n14340 0.00585714
R56157 VCC.n14362 VCC.n14361 0.00585714
R56158 VCC.n14374 VCC.n13878 0.00585714
R56159 VCC.n13869 VCC.n13862 0.00585714
R56160 VCC.n14391 VCC.n13863 0.00585714
R56161 VCC.n13913 VCC.n13902 0.00585714
R56162 VCC.n14335 VCC.n13900 0.00585714
R56163 VCC.n14363 VCC.n13883 0.00585714
R56164 VCC.n14861 VCC.n14465 0.00585714
R56165 VCC.n14888 VCC.n14887 0.00585714
R56166 VCC.n14925 VCC.n14432 0.00585714
R56167 VCC.n14924 VCC.n14923 0.00585714
R56168 VCC.n14421 VCC.n14418 0.00585714
R56169 VCC.n14940 VCC.n14939 0.00585714
R56170 VCC.n14469 VCC.n14454 0.00585714
R56171 VCC.n14902 VCC.n14901 0.00585714
R56172 VCC.n14926 VCC.n14430 0.00585714
R56173 VCC.n14729 VCC.n14534 0.00585714
R56174 VCC.n14736 VCC.n14729 0.00585714
R56175 VCC.n14763 VCC.n14520 0.00585714
R56176 VCC.n14798 VCC.n14498 0.00585714
R56177 VCC.n14843 VCC.n14842 0.00585714
R56178 VCC.n14781 VCC.n14496 0.00585714
R56179 VCC.n14818 VCC.n14479 0.00585714
R56180 VCC.n14615 VCC.n14605 0.00585714
R56181 VCC.n14647 VCC.n14646 0.00585714
R56182 VCC.n14567 VCC.n14559 0.00585714
R56183 VCC.n14596 VCC.n14583 0.00585714
R56184 VCC.n14654 VCC.n14653 0.00585714
R56185 VCC.n15165 VCC.n15155 0.00585714
R56186 VCC.n15197 VCC.n15196 0.00585714
R56187 VCC.n15117 VCC.n15109 0.00585714
R56188 VCC.n15146 VCC.n15133 0.00585714
R56189 VCC.n15204 VCC.n15203 0.00585714
R56190 VCC.n15290 VCC.n15279 0.00585714
R56191 VCC.n15287 VCC.n15279 0.00585714
R56192 VCC.n15314 VCC.n15071 0.00585714
R56193 VCC.n15349 VCC.n15049 0.00585714
R56194 VCC.n15393 VCC.n15392 0.00585714
R56195 VCC.n15332 VCC.n15047 0.00585714
R56196 VCC.n15369 VCC.n15030 0.00585714
R56197 VCC.n15411 VCC.n15017 0.00585714
R56198 VCC.n15448 VCC.n15447 0.00585714
R56199 VCC.n15469 VCC.n15468 0.00585714
R56200 VCC.n15481 VCC.n14985 0.00585714
R56201 VCC.n14976 VCC.n14969 0.00585714
R56202 VCC.n15498 VCC.n14970 0.00585714
R56203 VCC.n15020 VCC.n15009 0.00585714
R56204 VCC.n15442 VCC.n15007 0.00585714
R56205 VCC.n15470 VCC.n14990 0.00585714
R56206 VCC.n15968 VCC.n15572 0.00585714
R56207 VCC.n15995 VCC.n15994 0.00585714
R56208 VCC.n16032 VCC.n15539 0.00585714
R56209 VCC.n16031 VCC.n16030 0.00585714
R56210 VCC.n15528 VCC.n15525 0.00585714
R56211 VCC.n16047 VCC.n16046 0.00585714
R56212 VCC.n15576 VCC.n15561 0.00585714
R56213 VCC.n16009 VCC.n16008 0.00585714
R56214 VCC.n16033 VCC.n15537 0.00585714
R56215 VCC.n15836 VCC.n15641 0.00585714
R56216 VCC.n15843 VCC.n15836 0.00585714
R56217 VCC.n15870 VCC.n15627 0.00585714
R56218 VCC.n15905 VCC.n15605 0.00585714
R56219 VCC.n15950 VCC.n15949 0.00585714
R56220 VCC.n15888 VCC.n15603 0.00585714
R56221 VCC.n15925 VCC.n15586 0.00585714
R56222 VCC.n15722 VCC.n15712 0.00585714
R56223 VCC.n15754 VCC.n15753 0.00585714
R56224 VCC.n15674 VCC.n15666 0.00585714
R56225 VCC.n15703 VCC.n15690 0.00585714
R56226 VCC.n15761 VCC.n15760 0.00585714
R56227 VCC.n16272 VCC.n16262 0.00585714
R56228 VCC.n16304 VCC.n16303 0.00585714
R56229 VCC.n16224 VCC.n16216 0.00585714
R56230 VCC.n16253 VCC.n16240 0.00585714
R56231 VCC.n16311 VCC.n16310 0.00585714
R56232 VCC.n16397 VCC.n16386 0.00585714
R56233 VCC.n16394 VCC.n16386 0.00585714
R56234 VCC.n16421 VCC.n16178 0.00585714
R56235 VCC.n16456 VCC.n16156 0.00585714
R56236 VCC.n16500 VCC.n16499 0.00585714
R56237 VCC.n16439 VCC.n16154 0.00585714
R56238 VCC.n16476 VCC.n16137 0.00585714
R56239 VCC.n16518 VCC.n16124 0.00585714
R56240 VCC.n16555 VCC.n16554 0.00585714
R56241 VCC.n16576 VCC.n16575 0.00585714
R56242 VCC.n16588 VCC.n16092 0.00585714
R56243 VCC.n16083 VCC.n16076 0.00585714
R56244 VCC.n16605 VCC.n16077 0.00585714
R56245 VCC.n16127 VCC.n16116 0.00585714
R56246 VCC.n16549 VCC.n16114 0.00585714
R56247 VCC.n16577 VCC.n16097 0.00585714
R56248 VCC.n17075 VCC.n16679 0.00585714
R56249 VCC.n17102 VCC.n17101 0.00585714
R56250 VCC.n17139 VCC.n16646 0.00585714
R56251 VCC.n17138 VCC.n17137 0.00585714
R56252 VCC.n16635 VCC.n16632 0.00585714
R56253 VCC.n17154 VCC.n17153 0.00585714
R56254 VCC.n16683 VCC.n16668 0.00585714
R56255 VCC.n17116 VCC.n17115 0.00585714
R56256 VCC.n17140 VCC.n16644 0.00585714
R56257 VCC.n16943 VCC.n16748 0.00585714
R56258 VCC.n16950 VCC.n16943 0.00585714
R56259 VCC.n16977 VCC.n16734 0.00585714
R56260 VCC.n17012 VCC.n16712 0.00585714
R56261 VCC.n17057 VCC.n17056 0.00585714
R56262 VCC.n16995 VCC.n16710 0.00585714
R56263 VCC.n17032 VCC.n16693 0.00585714
R56264 VCC.n16829 VCC.n16819 0.00585714
R56265 VCC.n16861 VCC.n16860 0.00585714
R56266 VCC.n16781 VCC.n16773 0.00585714
R56267 VCC.n16810 VCC.n16797 0.00585714
R56268 VCC.n16868 VCC.n16867 0.00585714
R56269 VCC.n17317 VCC.n17306 0.00585714
R56270 VCC.n17314 VCC.n17306 0.00585714
R56271 VCC.n17341 VCC.n17285 0.00585714
R56272 VCC.n17376 VCC.n17263 0.00585714
R56273 VCC.n17420 VCC.n17419 0.00585714
R56274 VCC.n17359 VCC.n17261 0.00585714
R56275 VCC.n17396 VCC.n17244 0.00585714
R56276 VCC.n17438 VCC.n17231 0.00585714
R56277 VCC.n17475 VCC.n17474 0.00585714
R56278 VCC.n17496 VCC.n17495 0.00585714
R56279 VCC.n17508 VCC.n17199 0.00585714
R56280 VCC.n17190 VCC.n17183 0.00585714
R56281 VCC.n17525 VCC.n17184 0.00585714
R56282 VCC.n17234 VCC.n17223 0.00585714
R56283 VCC.n17469 VCC.n17221 0.00585714
R56284 VCC.n17497 VCC.n17204 0.00585714
R56285 VCC.n299 VCC.n137 0.00496429
R56286 VCC.n299 VCC.n298 0.00496429
R56287 VCC.n216 VCC.n189 0.00496429
R56288 VCC.n219 VCC.n187 0.00496429
R56289 VCC.n164 VCC.n148 0.00496429
R56290 VCC.n306 VCC.n132 0.00496429
R56291 VCC.n309 VCC.n128 0.00496429
R56292 VCC.n328 VCC.n327 0.00496429
R56293 VCC.n318 VCC.n126 0.00496429
R56294 VCC.n345 VCC.n344 0.00496429
R56295 VCC.n369 VCC.n368 0.00496429
R56296 VCC.n441 VCC.n71 0.00496429
R56297 VCC.n444 VCC.n67 0.00496429
R56298 VCC.n459 VCC.n63 0.00496429
R56299 VCC.n464 VCC.n61 0.00496429
R56300 VCC.n29 VCC.n14 0.00496429
R56301 VCC.n535 VCC.n14 0.00496429
R56302 VCC.n538 VCC.n1 0.00496429
R56303 VCC.n851 VCC.n689 0.00496429
R56304 VCC.n851 VCC.n850 0.00496429
R56305 VCC.n768 VCC.n741 0.00496429
R56306 VCC.n771 VCC.n739 0.00496429
R56307 VCC.n716 VCC.n700 0.00496429
R56308 VCC.n858 VCC.n684 0.00496429
R56309 VCC.n861 VCC.n680 0.00496429
R56310 VCC.n880 VCC.n879 0.00496429
R56311 VCC.n870 VCC.n678 0.00496429
R56312 VCC.n897 VCC.n896 0.00496429
R56313 VCC.n921 VCC.n920 0.00496429
R56314 VCC.n993 VCC.n623 0.00496429
R56315 VCC.n996 VCC.n619 0.00496429
R56316 VCC.n1011 VCC.n615 0.00496429
R56317 VCC.n1016 VCC.n613 0.00496429
R56318 VCC.n581 VCC.n566 0.00496429
R56319 VCC.n1087 VCC.n566 0.00496429
R56320 VCC.n1090 VCC.n555 0.00496429
R56321 VCC.n1570 VCC.n1172 0.00496429
R56322 VCC.n1573 VCC.n1170 0.00496429
R56323 VCC.n1631 VCC.n1127 0.00496429
R56324 VCC.n1634 VCC.n1127 0.00496429
R56325 VCC.n1637 VCC.n1109 0.00496429
R56326 VCC.n1437 VCC.n1436 0.00496429
R56327 VCC.n1428 VCC.n1236 0.00496429
R56328 VCC.n1454 VCC.n1453 0.00496429
R56329 VCC.n1478 VCC.n1477 0.00496429
R56330 VCC.n1551 VCC.n1180 0.00496429
R56331 VCC.n1554 VCC.n1176 0.00496429
R56332 VCC.n1409 VCC.n1247 0.00496429
R56333 VCC.n1409 VCC.n1408 0.00496429
R56334 VCC.n1326 VCC.n1299 0.00496429
R56335 VCC.n1329 VCC.n1297 0.00496429
R56336 VCC.n1274 VCC.n1258 0.00496429
R56337 VCC.n1416 VCC.n1242 0.00496429
R56338 VCC.n1419 VCC.n1238 0.00496429
R56339 VCC.n1960 VCC.n1798 0.00496429
R56340 VCC.n1960 VCC.n1959 0.00496429
R56341 VCC.n1877 VCC.n1850 0.00496429
R56342 VCC.n1880 VCC.n1848 0.00496429
R56343 VCC.n1825 VCC.n1809 0.00496429
R56344 VCC.n1967 VCC.n1793 0.00496429
R56345 VCC.n1970 VCC.n1789 0.00496429
R56346 VCC.n1989 VCC.n1988 0.00496429
R56347 VCC.n1979 VCC.n1787 0.00496429
R56348 VCC.n2006 VCC.n2005 0.00496429
R56349 VCC.n2030 VCC.n2029 0.00496429
R56350 VCC.n2102 VCC.n1732 0.00496429
R56351 VCC.n2105 VCC.n1728 0.00496429
R56352 VCC.n2120 VCC.n1724 0.00496429
R56353 VCC.n2125 VCC.n1722 0.00496429
R56354 VCC.n1690 VCC.n1675 0.00496429
R56355 VCC.n2196 VCC.n1675 0.00496429
R56356 VCC.n2199 VCC.n1664 0.00496429
R56357 VCC.n2679 VCC.n2281 0.00496429
R56358 VCC.n2682 VCC.n2279 0.00496429
R56359 VCC.n2740 VCC.n2236 0.00496429
R56360 VCC.n2743 VCC.n2236 0.00496429
R56361 VCC.n2746 VCC.n2218 0.00496429
R56362 VCC.n2546 VCC.n2545 0.00496429
R56363 VCC.n2537 VCC.n2345 0.00496429
R56364 VCC.n2563 VCC.n2562 0.00496429
R56365 VCC.n2587 VCC.n2586 0.00496429
R56366 VCC.n2660 VCC.n2289 0.00496429
R56367 VCC.n2663 VCC.n2285 0.00496429
R56368 VCC.n2518 VCC.n2356 0.00496429
R56369 VCC.n2518 VCC.n2517 0.00496429
R56370 VCC.n2435 VCC.n2408 0.00496429
R56371 VCC.n2438 VCC.n2406 0.00496429
R56372 VCC.n2383 VCC.n2367 0.00496429
R56373 VCC.n2525 VCC.n2351 0.00496429
R56374 VCC.n2528 VCC.n2347 0.00496429
R56375 VCC.n3069 VCC.n2907 0.00496429
R56376 VCC.n3069 VCC.n3068 0.00496429
R56377 VCC.n2986 VCC.n2959 0.00496429
R56378 VCC.n2989 VCC.n2957 0.00496429
R56379 VCC.n2934 VCC.n2918 0.00496429
R56380 VCC.n3076 VCC.n2902 0.00496429
R56381 VCC.n3079 VCC.n2898 0.00496429
R56382 VCC.n3098 VCC.n3097 0.00496429
R56383 VCC.n3088 VCC.n2896 0.00496429
R56384 VCC.n3115 VCC.n3114 0.00496429
R56385 VCC.n3139 VCC.n3138 0.00496429
R56386 VCC.n3211 VCC.n2841 0.00496429
R56387 VCC.n3214 VCC.n2837 0.00496429
R56388 VCC.n3229 VCC.n2833 0.00496429
R56389 VCC.n3234 VCC.n2831 0.00496429
R56390 VCC.n2799 VCC.n2784 0.00496429
R56391 VCC.n3305 VCC.n2784 0.00496429
R56392 VCC.n3308 VCC.n2773 0.00496429
R56393 VCC.n3788 VCC.n3390 0.00496429
R56394 VCC.n3791 VCC.n3388 0.00496429
R56395 VCC.n3849 VCC.n3345 0.00496429
R56396 VCC.n3852 VCC.n3345 0.00496429
R56397 VCC.n3855 VCC.n3327 0.00496429
R56398 VCC.n3655 VCC.n3654 0.00496429
R56399 VCC.n3646 VCC.n3454 0.00496429
R56400 VCC.n3672 VCC.n3671 0.00496429
R56401 VCC.n3696 VCC.n3695 0.00496429
R56402 VCC.n3769 VCC.n3398 0.00496429
R56403 VCC.n3772 VCC.n3394 0.00496429
R56404 VCC.n3627 VCC.n3465 0.00496429
R56405 VCC.n3627 VCC.n3626 0.00496429
R56406 VCC.n3544 VCC.n3517 0.00496429
R56407 VCC.n3547 VCC.n3515 0.00496429
R56408 VCC.n3492 VCC.n3476 0.00496429
R56409 VCC.n3634 VCC.n3460 0.00496429
R56410 VCC.n3637 VCC.n3456 0.00496429
R56411 VCC.n4178 VCC.n4016 0.00496429
R56412 VCC.n4178 VCC.n4177 0.00496429
R56413 VCC.n4095 VCC.n4068 0.00496429
R56414 VCC.n4098 VCC.n4066 0.00496429
R56415 VCC.n4043 VCC.n4027 0.00496429
R56416 VCC.n4185 VCC.n4011 0.00496429
R56417 VCC.n4188 VCC.n4007 0.00496429
R56418 VCC.n4207 VCC.n4206 0.00496429
R56419 VCC.n4197 VCC.n4005 0.00496429
R56420 VCC.n4224 VCC.n4223 0.00496429
R56421 VCC.n4248 VCC.n4247 0.00496429
R56422 VCC.n4320 VCC.n3950 0.00496429
R56423 VCC.n4323 VCC.n3946 0.00496429
R56424 VCC.n4338 VCC.n3942 0.00496429
R56425 VCC.n4343 VCC.n3940 0.00496429
R56426 VCC.n3908 VCC.n3893 0.00496429
R56427 VCC.n4414 VCC.n3893 0.00496429
R56428 VCC.n4417 VCC.n3882 0.00496429
R56429 VCC.n4897 VCC.n4499 0.00496429
R56430 VCC.n4900 VCC.n4497 0.00496429
R56431 VCC.n4958 VCC.n4454 0.00496429
R56432 VCC.n4961 VCC.n4454 0.00496429
R56433 VCC.n4964 VCC.n4436 0.00496429
R56434 VCC.n4764 VCC.n4763 0.00496429
R56435 VCC.n4755 VCC.n4563 0.00496429
R56436 VCC.n4781 VCC.n4780 0.00496429
R56437 VCC.n4805 VCC.n4804 0.00496429
R56438 VCC.n4878 VCC.n4507 0.00496429
R56439 VCC.n4881 VCC.n4503 0.00496429
R56440 VCC.n4736 VCC.n4574 0.00496429
R56441 VCC.n4736 VCC.n4735 0.00496429
R56442 VCC.n4653 VCC.n4626 0.00496429
R56443 VCC.n4656 VCC.n4624 0.00496429
R56444 VCC.n4601 VCC.n4585 0.00496429
R56445 VCC.n4743 VCC.n4569 0.00496429
R56446 VCC.n4746 VCC.n4565 0.00496429
R56447 VCC.n5287 VCC.n5125 0.00496429
R56448 VCC.n5287 VCC.n5286 0.00496429
R56449 VCC.n5204 VCC.n5177 0.00496429
R56450 VCC.n5207 VCC.n5175 0.00496429
R56451 VCC.n5152 VCC.n5136 0.00496429
R56452 VCC.n5294 VCC.n5120 0.00496429
R56453 VCC.n5297 VCC.n5116 0.00496429
R56454 VCC.n5316 VCC.n5315 0.00496429
R56455 VCC.n5306 VCC.n5114 0.00496429
R56456 VCC.n5333 VCC.n5332 0.00496429
R56457 VCC.n5357 VCC.n5356 0.00496429
R56458 VCC.n5429 VCC.n5059 0.00496429
R56459 VCC.n5432 VCC.n5055 0.00496429
R56460 VCC.n5447 VCC.n5051 0.00496429
R56461 VCC.n5452 VCC.n5049 0.00496429
R56462 VCC.n5017 VCC.n5002 0.00496429
R56463 VCC.n5523 VCC.n5002 0.00496429
R56464 VCC.n5526 VCC.n4991 0.00496429
R56465 VCC.n6006 VCC.n5608 0.00496429
R56466 VCC.n6009 VCC.n5606 0.00496429
R56467 VCC.n6067 VCC.n5563 0.00496429
R56468 VCC.n6070 VCC.n5563 0.00496429
R56469 VCC.n6073 VCC.n5545 0.00496429
R56470 VCC.n5873 VCC.n5872 0.00496429
R56471 VCC.n5864 VCC.n5672 0.00496429
R56472 VCC.n5890 VCC.n5889 0.00496429
R56473 VCC.n5914 VCC.n5913 0.00496429
R56474 VCC.n5987 VCC.n5616 0.00496429
R56475 VCC.n5990 VCC.n5612 0.00496429
R56476 VCC.n5845 VCC.n5683 0.00496429
R56477 VCC.n5845 VCC.n5844 0.00496429
R56478 VCC.n5762 VCC.n5735 0.00496429
R56479 VCC.n5765 VCC.n5733 0.00496429
R56480 VCC.n5710 VCC.n5694 0.00496429
R56481 VCC.n5852 VCC.n5678 0.00496429
R56482 VCC.n5855 VCC.n5674 0.00496429
R56483 VCC.n6396 VCC.n6234 0.00496429
R56484 VCC.n6396 VCC.n6395 0.00496429
R56485 VCC.n6313 VCC.n6286 0.00496429
R56486 VCC.n6316 VCC.n6284 0.00496429
R56487 VCC.n6261 VCC.n6245 0.00496429
R56488 VCC.n6403 VCC.n6229 0.00496429
R56489 VCC.n6406 VCC.n6225 0.00496429
R56490 VCC.n6425 VCC.n6424 0.00496429
R56491 VCC.n6415 VCC.n6223 0.00496429
R56492 VCC.n6442 VCC.n6441 0.00496429
R56493 VCC.n6466 VCC.n6465 0.00496429
R56494 VCC.n6538 VCC.n6168 0.00496429
R56495 VCC.n6541 VCC.n6164 0.00496429
R56496 VCC.n6556 VCC.n6160 0.00496429
R56497 VCC.n6561 VCC.n6158 0.00496429
R56498 VCC.n6126 VCC.n6111 0.00496429
R56499 VCC.n6632 VCC.n6111 0.00496429
R56500 VCC.n6635 VCC.n6100 0.00496429
R56501 VCC.n7115 VCC.n6717 0.00496429
R56502 VCC.n7118 VCC.n6715 0.00496429
R56503 VCC.n7176 VCC.n6672 0.00496429
R56504 VCC.n7179 VCC.n6672 0.00496429
R56505 VCC.n7182 VCC.n6654 0.00496429
R56506 VCC.n6982 VCC.n6981 0.00496429
R56507 VCC.n6973 VCC.n6781 0.00496429
R56508 VCC.n6999 VCC.n6998 0.00496429
R56509 VCC.n7023 VCC.n7022 0.00496429
R56510 VCC.n7096 VCC.n6725 0.00496429
R56511 VCC.n7099 VCC.n6721 0.00496429
R56512 VCC.n6954 VCC.n6792 0.00496429
R56513 VCC.n6954 VCC.n6953 0.00496429
R56514 VCC.n6871 VCC.n6844 0.00496429
R56515 VCC.n6874 VCC.n6842 0.00496429
R56516 VCC.n6819 VCC.n6803 0.00496429
R56517 VCC.n6961 VCC.n6787 0.00496429
R56518 VCC.n6964 VCC.n6783 0.00496429
R56519 VCC.n7505 VCC.n7343 0.00496429
R56520 VCC.n7505 VCC.n7504 0.00496429
R56521 VCC.n7422 VCC.n7395 0.00496429
R56522 VCC.n7425 VCC.n7393 0.00496429
R56523 VCC.n7370 VCC.n7354 0.00496429
R56524 VCC.n7512 VCC.n7338 0.00496429
R56525 VCC.n7515 VCC.n7334 0.00496429
R56526 VCC.n7534 VCC.n7533 0.00496429
R56527 VCC.n7524 VCC.n7332 0.00496429
R56528 VCC.n7551 VCC.n7550 0.00496429
R56529 VCC.n7575 VCC.n7574 0.00496429
R56530 VCC.n7647 VCC.n7277 0.00496429
R56531 VCC.n7650 VCC.n7273 0.00496429
R56532 VCC.n7665 VCC.n7269 0.00496429
R56533 VCC.n7670 VCC.n7267 0.00496429
R56534 VCC.n7235 VCC.n7220 0.00496429
R56535 VCC.n7741 VCC.n7220 0.00496429
R56536 VCC.n7744 VCC.n7209 0.00496429
R56537 VCC.n8224 VCC.n7826 0.00496429
R56538 VCC.n8227 VCC.n7824 0.00496429
R56539 VCC.n8285 VCC.n7781 0.00496429
R56540 VCC.n8288 VCC.n7781 0.00496429
R56541 VCC.n8291 VCC.n7763 0.00496429
R56542 VCC.n8091 VCC.n8090 0.00496429
R56543 VCC.n8082 VCC.n7890 0.00496429
R56544 VCC.n8108 VCC.n8107 0.00496429
R56545 VCC.n8132 VCC.n8131 0.00496429
R56546 VCC.n8205 VCC.n7834 0.00496429
R56547 VCC.n8208 VCC.n7830 0.00496429
R56548 VCC.n8063 VCC.n7901 0.00496429
R56549 VCC.n8063 VCC.n8062 0.00496429
R56550 VCC.n7980 VCC.n7953 0.00496429
R56551 VCC.n7983 VCC.n7951 0.00496429
R56552 VCC.n7928 VCC.n7912 0.00496429
R56553 VCC.n8070 VCC.n7896 0.00496429
R56554 VCC.n8073 VCC.n7892 0.00496429
R56555 VCC.n8643 VCC.n8642 0.00496429
R56556 VCC.n8633 VCC.n8441 0.00496429
R56557 VCC.n8660 VCC.n8659 0.00496429
R56558 VCC.n8684 VCC.n8683 0.00496429
R56559 VCC.n8756 VCC.n8386 0.00496429
R56560 VCC.n8759 VCC.n8382 0.00496429
R56561 VCC.n8774 VCC.n8378 0.00496429
R56562 VCC.n8779 VCC.n8376 0.00496429
R56563 VCC.n8344 VCC.n8329 0.00496429
R56564 VCC.n8850 VCC.n8329 0.00496429
R56565 VCC.n8853 VCC.n8318 0.00496429
R56566 VCC.n8614 VCC.n8452 0.00496429
R56567 VCC.n8614 VCC.n8613 0.00496429
R56568 VCC.n8531 VCC.n8504 0.00496429
R56569 VCC.n8534 VCC.n8502 0.00496429
R56570 VCC.n8479 VCC.n8463 0.00496429
R56571 VCC.n8621 VCC.n8447 0.00496429
R56572 VCC.n8624 VCC.n8443 0.00496429
R56573 VCC.n9333 VCC.n8935 0.00496429
R56574 VCC.n9336 VCC.n8933 0.00496429
R56575 VCC.n9394 VCC.n8890 0.00496429
R56576 VCC.n9397 VCC.n8890 0.00496429
R56577 VCC.n9400 VCC.n8872 0.00496429
R56578 VCC.n9200 VCC.n9199 0.00496429
R56579 VCC.n9191 VCC.n8999 0.00496429
R56580 VCC.n9217 VCC.n9216 0.00496429
R56581 VCC.n9241 VCC.n9240 0.00496429
R56582 VCC.n9314 VCC.n8943 0.00496429
R56583 VCC.n9317 VCC.n8939 0.00496429
R56584 VCC.n9172 VCC.n9010 0.00496429
R56585 VCC.n9172 VCC.n9171 0.00496429
R56586 VCC.n9089 VCC.n9062 0.00496429
R56587 VCC.n9092 VCC.n9060 0.00496429
R56588 VCC.n9037 VCC.n9021 0.00496429
R56589 VCC.n9179 VCC.n9005 0.00496429
R56590 VCC.n9182 VCC.n9001 0.00496429
R56591 VCC.n9723 VCC.n9561 0.00496429
R56592 VCC.n9723 VCC.n9722 0.00496429
R56593 VCC.n9640 VCC.n9613 0.00496429
R56594 VCC.n9643 VCC.n9611 0.00496429
R56595 VCC.n9588 VCC.n9572 0.00496429
R56596 VCC.n9730 VCC.n9556 0.00496429
R56597 VCC.n9733 VCC.n9552 0.00496429
R56598 VCC.n9752 VCC.n9751 0.00496429
R56599 VCC.n9742 VCC.n9550 0.00496429
R56600 VCC.n9769 VCC.n9768 0.00496429
R56601 VCC.n9793 VCC.n9792 0.00496429
R56602 VCC.n9865 VCC.n9495 0.00496429
R56603 VCC.n9868 VCC.n9491 0.00496429
R56604 VCC.n9883 VCC.n9487 0.00496429
R56605 VCC.n9888 VCC.n9485 0.00496429
R56606 VCC.n9453 VCC.n9438 0.00496429
R56607 VCC.n9959 VCC.n9438 0.00496429
R56608 VCC.n9962 VCC.n9427 0.00496429
R56609 VCC.n10441 VCC.n10043 0.00496429
R56610 VCC.n10444 VCC.n10041 0.00496429
R56611 VCC.n10502 VCC.n9998 0.00496429
R56612 VCC.n10505 VCC.n9998 0.00496429
R56613 VCC.n10508 VCC.n9980 0.00496429
R56614 VCC.n10308 VCC.n10307 0.00496429
R56615 VCC.n10299 VCC.n10107 0.00496429
R56616 VCC.n10325 VCC.n10324 0.00496429
R56617 VCC.n10349 VCC.n10348 0.00496429
R56618 VCC.n10422 VCC.n10051 0.00496429
R56619 VCC.n10425 VCC.n10047 0.00496429
R56620 VCC.n10280 VCC.n10118 0.00496429
R56621 VCC.n10280 VCC.n10279 0.00496429
R56622 VCC.n10197 VCC.n10170 0.00496429
R56623 VCC.n10200 VCC.n10168 0.00496429
R56624 VCC.n10145 VCC.n10129 0.00496429
R56625 VCC.n10287 VCC.n10113 0.00496429
R56626 VCC.n10290 VCC.n10109 0.00496429
R56627 VCC.n10830 VCC.n10668 0.00496429
R56628 VCC.n10830 VCC.n10829 0.00496429
R56629 VCC.n10747 VCC.n10720 0.00496429
R56630 VCC.n10750 VCC.n10718 0.00496429
R56631 VCC.n10695 VCC.n10679 0.00496429
R56632 VCC.n10837 VCC.n10663 0.00496429
R56633 VCC.n10840 VCC.n10659 0.00496429
R56634 VCC.n10859 VCC.n10858 0.00496429
R56635 VCC.n10849 VCC.n10657 0.00496429
R56636 VCC.n10876 VCC.n10875 0.00496429
R56637 VCC.n10900 VCC.n10899 0.00496429
R56638 VCC.n10972 VCC.n10602 0.00496429
R56639 VCC.n10975 VCC.n10598 0.00496429
R56640 VCC.n10990 VCC.n10594 0.00496429
R56641 VCC.n10995 VCC.n10592 0.00496429
R56642 VCC.n10560 VCC.n10545 0.00496429
R56643 VCC.n11066 VCC.n10545 0.00496429
R56644 VCC.n11069 VCC.n10534 0.00496429
R56645 VCC.n11548 VCC.n11150 0.00496429
R56646 VCC.n11551 VCC.n11148 0.00496429
R56647 VCC.n11609 VCC.n11105 0.00496429
R56648 VCC.n11612 VCC.n11105 0.00496429
R56649 VCC.n11615 VCC.n11087 0.00496429
R56650 VCC.n11415 VCC.n11414 0.00496429
R56651 VCC.n11406 VCC.n11214 0.00496429
R56652 VCC.n11432 VCC.n11431 0.00496429
R56653 VCC.n11456 VCC.n11455 0.00496429
R56654 VCC.n11529 VCC.n11158 0.00496429
R56655 VCC.n11532 VCC.n11154 0.00496429
R56656 VCC.n11387 VCC.n11225 0.00496429
R56657 VCC.n11387 VCC.n11386 0.00496429
R56658 VCC.n11304 VCC.n11277 0.00496429
R56659 VCC.n11307 VCC.n11275 0.00496429
R56660 VCC.n11252 VCC.n11236 0.00496429
R56661 VCC.n11394 VCC.n11220 0.00496429
R56662 VCC.n11397 VCC.n11216 0.00496429
R56663 VCC.n11937 VCC.n11775 0.00496429
R56664 VCC.n11937 VCC.n11936 0.00496429
R56665 VCC.n11854 VCC.n11827 0.00496429
R56666 VCC.n11857 VCC.n11825 0.00496429
R56667 VCC.n11802 VCC.n11786 0.00496429
R56668 VCC.n11944 VCC.n11770 0.00496429
R56669 VCC.n11947 VCC.n11766 0.00496429
R56670 VCC.n11966 VCC.n11965 0.00496429
R56671 VCC.n11956 VCC.n11764 0.00496429
R56672 VCC.n11983 VCC.n11982 0.00496429
R56673 VCC.n12007 VCC.n12006 0.00496429
R56674 VCC.n12079 VCC.n11709 0.00496429
R56675 VCC.n12082 VCC.n11705 0.00496429
R56676 VCC.n12097 VCC.n11701 0.00496429
R56677 VCC.n12102 VCC.n11699 0.00496429
R56678 VCC.n11667 VCC.n11652 0.00496429
R56679 VCC.n12173 VCC.n11652 0.00496429
R56680 VCC.n12176 VCC.n11641 0.00496429
R56681 VCC.n12655 VCC.n12257 0.00496429
R56682 VCC.n12658 VCC.n12255 0.00496429
R56683 VCC.n12716 VCC.n12212 0.00496429
R56684 VCC.n12719 VCC.n12212 0.00496429
R56685 VCC.n12722 VCC.n12194 0.00496429
R56686 VCC.n12522 VCC.n12521 0.00496429
R56687 VCC.n12513 VCC.n12321 0.00496429
R56688 VCC.n12539 VCC.n12538 0.00496429
R56689 VCC.n12563 VCC.n12562 0.00496429
R56690 VCC.n12636 VCC.n12265 0.00496429
R56691 VCC.n12639 VCC.n12261 0.00496429
R56692 VCC.n12494 VCC.n12332 0.00496429
R56693 VCC.n12494 VCC.n12493 0.00496429
R56694 VCC.n12411 VCC.n12384 0.00496429
R56695 VCC.n12414 VCC.n12382 0.00496429
R56696 VCC.n12359 VCC.n12343 0.00496429
R56697 VCC.n12501 VCC.n12327 0.00496429
R56698 VCC.n12504 VCC.n12323 0.00496429
R56699 VCC.n13044 VCC.n12882 0.00496429
R56700 VCC.n13044 VCC.n13043 0.00496429
R56701 VCC.n12961 VCC.n12934 0.00496429
R56702 VCC.n12964 VCC.n12932 0.00496429
R56703 VCC.n12909 VCC.n12893 0.00496429
R56704 VCC.n13051 VCC.n12877 0.00496429
R56705 VCC.n13054 VCC.n12873 0.00496429
R56706 VCC.n13073 VCC.n13072 0.00496429
R56707 VCC.n13063 VCC.n12871 0.00496429
R56708 VCC.n13090 VCC.n13089 0.00496429
R56709 VCC.n13114 VCC.n13113 0.00496429
R56710 VCC.n13186 VCC.n12816 0.00496429
R56711 VCC.n13189 VCC.n12812 0.00496429
R56712 VCC.n13204 VCC.n12808 0.00496429
R56713 VCC.n13209 VCC.n12806 0.00496429
R56714 VCC.n12774 VCC.n12759 0.00496429
R56715 VCC.n13280 VCC.n12759 0.00496429
R56716 VCC.n13283 VCC.n12748 0.00496429
R56717 VCC.n13762 VCC.n13364 0.00496429
R56718 VCC.n13765 VCC.n13362 0.00496429
R56719 VCC.n13823 VCC.n13319 0.00496429
R56720 VCC.n13826 VCC.n13319 0.00496429
R56721 VCC.n13829 VCC.n13301 0.00496429
R56722 VCC.n13629 VCC.n13628 0.00496429
R56723 VCC.n13620 VCC.n13428 0.00496429
R56724 VCC.n13646 VCC.n13645 0.00496429
R56725 VCC.n13670 VCC.n13669 0.00496429
R56726 VCC.n13743 VCC.n13372 0.00496429
R56727 VCC.n13746 VCC.n13368 0.00496429
R56728 VCC.n13601 VCC.n13439 0.00496429
R56729 VCC.n13601 VCC.n13600 0.00496429
R56730 VCC.n13518 VCC.n13491 0.00496429
R56731 VCC.n13521 VCC.n13489 0.00496429
R56732 VCC.n13466 VCC.n13450 0.00496429
R56733 VCC.n13608 VCC.n13434 0.00496429
R56734 VCC.n13611 VCC.n13430 0.00496429
R56735 VCC.n14151 VCC.n13989 0.00496429
R56736 VCC.n14151 VCC.n14150 0.00496429
R56737 VCC.n14068 VCC.n14041 0.00496429
R56738 VCC.n14071 VCC.n14039 0.00496429
R56739 VCC.n14016 VCC.n14000 0.00496429
R56740 VCC.n14158 VCC.n13984 0.00496429
R56741 VCC.n14161 VCC.n13980 0.00496429
R56742 VCC.n14180 VCC.n14179 0.00496429
R56743 VCC.n14170 VCC.n13978 0.00496429
R56744 VCC.n14197 VCC.n14196 0.00496429
R56745 VCC.n14221 VCC.n14220 0.00496429
R56746 VCC.n14293 VCC.n13923 0.00496429
R56747 VCC.n14296 VCC.n13919 0.00496429
R56748 VCC.n14311 VCC.n13915 0.00496429
R56749 VCC.n14316 VCC.n13913 0.00496429
R56750 VCC.n13881 VCC.n13866 0.00496429
R56751 VCC.n14387 VCC.n13866 0.00496429
R56752 VCC.n14390 VCC.n13855 0.00496429
R56753 VCC.n14869 VCC.n14471 0.00496429
R56754 VCC.n14872 VCC.n14469 0.00496429
R56755 VCC.n14930 VCC.n14426 0.00496429
R56756 VCC.n14933 VCC.n14426 0.00496429
R56757 VCC.n14936 VCC.n14408 0.00496429
R56758 VCC.n14736 VCC.n14735 0.00496429
R56759 VCC.n14727 VCC.n14535 0.00496429
R56760 VCC.n14753 VCC.n14752 0.00496429
R56761 VCC.n14777 VCC.n14776 0.00496429
R56762 VCC.n14850 VCC.n14479 0.00496429
R56763 VCC.n14853 VCC.n14475 0.00496429
R56764 VCC.n14708 VCC.n14546 0.00496429
R56765 VCC.n14708 VCC.n14707 0.00496429
R56766 VCC.n14625 VCC.n14598 0.00496429
R56767 VCC.n14628 VCC.n14596 0.00496429
R56768 VCC.n14573 VCC.n14557 0.00496429
R56769 VCC.n14715 VCC.n14541 0.00496429
R56770 VCC.n14718 VCC.n14537 0.00496429
R56771 VCC.n15258 VCC.n15096 0.00496429
R56772 VCC.n15258 VCC.n15257 0.00496429
R56773 VCC.n15175 VCC.n15148 0.00496429
R56774 VCC.n15178 VCC.n15146 0.00496429
R56775 VCC.n15123 VCC.n15107 0.00496429
R56776 VCC.n15265 VCC.n15091 0.00496429
R56777 VCC.n15268 VCC.n15087 0.00496429
R56778 VCC.n15287 VCC.n15286 0.00496429
R56779 VCC.n15277 VCC.n15085 0.00496429
R56780 VCC.n15304 VCC.n15303 0.00496429
R56781 VCC.n15328 VCC.n15327 0.00496429
R56782 VCC.n15400 VCC.n15030 0.00496429
R56783 VCC.n15403 VCC.n15026 0.00496429
R56784 VCC.n15418 VCC.n15022 0.00496429
R56785 VCC.n15423 VCC.n15020 0.00496429
R56786 VCC.n14988 VCC.n14973 0.00496429
R56787 VCC.n15494 VCC.n14973 0.00496429
R56788 VCC.n15497 VCC.n14962 0.00496429
R56789 VCC.n15976 VCC.n15578 0.00496429
R56790 VCC.n15979 VCC.n15576 0.00496429
R56791 VCC.n16037 VCC.n15533 0.00496429
R56792 VCC.n16040 VCC.n15533 0.00496429
R56793 VCC.n16043 VCC.n15515 0.00496429
R56794 VCC.n15843 VCC.n15842 0.00496429
R56795 VCC.n15834 VCC.n15642 0.00496429
R56796 VCC.n15860 VCC.n15859 0.00496429
R56797 VCC.n15884 VCC.n15883 0.00496429
R56798 VCC.n15957 VCC.n15586 0.00496429
R56799 VCC.n15960 VCC.n15582 0.00496429
R56800 VCC.n15815 VCC.n15653 0.00496429
R56801 VCC.n15815 VCC.n15814 0.00496429
R56802 VCC.n15732 VCC.n15705 0.00496429
R56803 VCC.n15735 VCC.n15703 0.00496429
R56804 VCC.n15680 VCC.n15664 0.00496429
R56805 VCC.n15822 VCC.n15648 0.00496429
R56806 VCC.n15825 VCC.n15644 0.00496429
R56807 VCC.n16365 VCC.n16203 0.00496429
R56808 VCC.n16365 VCC.n16364 0.00496429
R56809 VCC.n16282 VCC.n16255 0.00496429
R56810 VCC.n16285 VCC.n16253 0.00496429
R56811 VCC.n16230 VCC.n16214 0.00496429
R56812 VCC.n16372 VCC.n16198 0.00496429
R56813 VCC.n16375 VCC.n16194 0.00496429
R56814 VCC.n16394 VCC.n16393 0.00496429
R56815 VCC.n16384 VCC.n16192 0.00496429
R56816 VCC.n16411 VCC.n16410 0.00496429
R56817 VCC.n16435 VCC.n16434 0.00496429
R56818 VCC.n16507 VCC.n16137 0.00496429
R56819 VCC.n16510 VCC.n16133 0.00496429
R56820 VCC.n16525 VCC.n16129 0.00496429
R56821 VCC.n16530 VCC.n16127 0.00496429
R56822 VCC.n16095 VCC.n16080 0.00496429
R56823 VCC.n16601 VCC.n16080 0.00496429
R56824 VCC.n16604 VCC.n16069 0.00496429
R56825 VCC.n17083 VCC.n16685 0.00496429
R56826 VCC.n17086 VCC.n16683 0.00496429
R56827 VCC.n17144 VCC.n16640 0.00496429
R56828 VCC.n17147 VCC.n16640 0.00496429
R56829 VCC.n17150 VCC.n16622 0.00496429
R56830 VCC.n16950 VCC.n16949 0.00496429
R56831 VCC.n16941 VCC.n16749 0.00496429
R56832 VCC.n16967 VCC.n16966 0.00496429
R56833 VCC.n16991 VCC.n16990 0.00496429
R56834 VCC.n17064 VCC.n16693 0.00496429
R56835 VCC.n17067 VCC.n16689 0.00496429
R56836 VCC.n16922 VCC.n16760 0.00496429
R56837 VCC.n16922 VCC.n16921 0.00496429
R56838 VCC.n16839 VCC.n16812 0.00496429
R56839 VCC.n16842 VCC.n16810 0.00496429
R56840 VCC.n16787 VCC.n16771 0.00496429
R56841 VCC.n16929 VCC.n16755 0.00496429
R56842 VCC.n16932 VCC.n16751 0.00496429
R56843 VCC.n17314 VCC.n17313 0.00496429
R56844 VCC.n17304 VCC.n17299 0.00496429
R56845 VCC.n17331 VCC.n17330 0.00496429
R56846 VCC.n17355 VCC.n17354 0.00496429
R56847 VCC.n17427 VCC.n17244 0.00496429
R56848 VCC.n17430 VCC.n17240 0.00496429
R56849 VCC.n17445 VCC.n17236 0.00496429
R56850 VCC.n17450 VCC.n17234 0.00496429
R56851 VCC.n17202 VCC.n17187 0.00496429
R56852 VCC.n17521 VCC.n17187 0.00496429
R56853 VCC.n17524 VCC.n17176 0.00496429
R56854 VCC.n243 VCC.n242 0.00486429
R56855 VCC.n257 VCC.n165 0.00486429
R56856 VCC.n259 VCC.n258 0.00486429
R56857 VCC.n280 VCC.n147 0.00486429
R56858 VCC.n370 VCC.n102 0.00486429
R56859 VCC.n380 VCC.n371 0.00486429
R56860 VCC.n379 VCC.n372 0.00486429
R56861 VCC.n407 VCC.n87 0.00486429
R56862 VCC.n485 VCC.n484 0.00486429
R56863 VCC.n503 VCC.n35 0.00486429
R56864 VCC.n505 VCC.n504 0.00486429
R56865 VCC.n512 VCC.n30 0.00486429
R56866 VCC.n795 VCC.n794 0.00486429
R56867 VCC.n809 VCC.n717 0.00486429
R56868 VCC.n811 VCC.n810 0.00486429
R56869 VCC.n832 VCC.n699 0.00486429
R56870 VCC.n922 VCC.n654 0.00486429
R56871 VCC.n932 VCC.n923 0.00486429
R56872 VCC.n931 VCC.n924 0.00486429
R56873 VCC.n959 VCC.n639 0.00486429
R56874 VCC.n1037 VCC.n1036 0.00486429
R56875 VCC.n1055 VCC.n587 0.00486429
R56876 VCC.n1057 VCC.n1056 0.00486429
R56877 VCC.n1064 VCC.n582 0.00486429
R56878 VCC.n1353 VCC.n1352 0.00486429
R56879 VCC.n1367 VCC.n1275 0.00486429
R56880 VCC.n1369 VCC.n1368 0.00486429
R56881 VCC.n1390 VCC.n1257 0.00486429
R56882 VCC.n1479 VCC.n1211 0.00486429
R56883 VCC.n1489 VCC.n1480 0.00486429
R56884 VCC.n1488 VCC.n1481 0.00486429
R56885 VCC.n1516 VCC.n1196 0.00486429
R56886 VCC.n1601 VCC.n1600 0.00486429
R56887 VCC.n1608 VCC.n1150 0.00486429
R56888 VCC.n1612 VCC.n1611 0.00486429
R56889 VCC.n1628 VCC.n1130 0.00486429
R56890 VCC.n1904 VCC.n1903 0.00486429
R56891 VCC.n1918 VCC.n1826 0.00486429
R56892 VCC.n1920 VCC.n1919 0.00486429
R56893 VCC.n1941 VCC.n1808 0.00486429
R56894 VCC.n2031 VCC.n1763 0.00486429
R56895 VCC.n2041 VCC.n2032 0.00486429
R56896 VCC.n2040 VCC.n2033 0.00486429
R56897 VCC.n2068 VCC.n1748 0.00486429
R56898 VCC.n2146 VCC.n2145 0.00486429
R56899 VCC.n2164 VCC.n1696 0.00486429
R56900 VCC.n2166 VCC.n2165 0.00486429
R56901 VCC.n2173 VCC.n1691 0.00486429
R56902 VCC.n2462 VCC.n2461 0.00486429
R56903 VCC.n2476 VCC.n2384 0.00486429
R56904 VCC.n2478 VCC.n2477 0.00486429
R56905 VCC.n2499 VCC.n2366 0.00486429
R56906 VCC.n2588 VCC.n2320 0.00486429
R56907 VCC.n2598 VCC.n2589 0.00486429
R56908 VCC.n2597 VCC.n2590 0.00486429
R56909 VCC.n2625 VCC.n2305 0.00486429
R56910 VCC.n2710 VCC.n2709 0.00486429
R56911 VCC.n2717 VCC.n2259 0.00486429
R56912 VCC.n2721 VCC.n2720 0.00486429
R56913 VCC.n2737 VCC.n2239 0.00486429
R56914 VCC.n3013 VCC.n3012 0.00486429
R56915 VCC.n3027 VCC.n2935 0.00486429
R56916 VCC.n3029 VCC.n3028 0.00486429
R56917 VCC.n3050 VCC.n2917 0.00486429
R56918 VCC.n3140 VCC.n2872 0.00486429
R56919 VCC.n3150 VCC.n3141 0.00486429
R56920 VCC.n3149 VCC.n3142 0.00486429
R56921 VCC.n3177 VCC.n2857 0.00486429
R56922 VCC.n3255 VCC.n3254 0.00486429
R56923 VCC.n3273 VCC.n2805 0.00486429
R56924 VCC.n3275 VCC.n3274 0.00486429
R56925 VCC.n3282 VCC.n2800 0.00486429
R56926 VCC.n3571 VCC.n3570 0.00486429
R56927 VCC.n3585 VCC.n3493 0.00486429
R56928 VCC.n3587 VCC.n3586 0.00486429
R56929 VCC.n3608 VCC.n3475 0.00486429
R56930 VCC.n3697 VCC.n3429 0.00486429
R56931 VCC.n3707 VCC.n3698 0.00486429
R56932 VCC.n3706 VCC.n3699 0.00486429
R56933 VCC.n3734 VCC.n3414 0.00486429
R56934 VCC.n3819 VCC.n3818 0.00486429
R56935 VCC.n3826 VCC.n3368 0.00486429
R56936 VCC.n3830 VCC.n3829 0.00486429
R56937 VCC.n3846 VCC.n3348 0.00486429
R56938 VCC.n4122 VCC.n4121 0.00486429
R56939 VCC.n4136 VCC.n4044 0.00486429
R56940 VCC.n4138 VCC.n4137 0.00486429
R56941 VCC.n4159 VCC.n4026 0.00486429
R56942 VCC.n4249 VCC.n3981 0.00486429
R56943 VCC.n4259 VCC.n4250 0.00486429
R56944 VCC.n4258 VCC.n4251 0.00486429
R56945 VCC.n4286 VCC.n3966 0.00486429
R56946 VCC.n4364 VCC.n4363 0.00486429
R56947 VCC.n4382 VCC.n3914 0.00486429
R56948 VCC.n4384 VCC.n4383 0.00486429
R56949 VCC.n4391 VCC.n3909 0.00486429
R56950 VCC.n4680 VCC.n4679 0.00486429
R56951 VCC.n4694 VCC.n4602 0.00486429
R56952 VCC.n4696 VCC.n4695 0.00486429
R56953 VCC.n4717 VCC.n4584 0.00486429
R56954 VCC.n4806 VCC.n4538 0.00486429
R56955 VCC.n4816 VCC.n4807 0.00486429
R56956 VCC.n4815 VCC.n4808 0.00486429
R56957 VCC.n4843 VCC.n4523 0.00486429
R56958 VCC.n4928 VCC.n4927 0.00486429
R56959 VCC.n4935 VCC.n4477 0.00486429
R56960 VCC.n4939 VCC.n4938 0.00486429
R56961 VCC.n4955 VCC.n4457 0.00486429
R56962 VCC.n5231 VCC.n5230 0.00486429
R56963 VCC.n5245 VCC.n5153 0.00486429
R56964 VCC.n5247 VCC.n5246 0.00486429
R56965 VCC.n5268 VCC.n5135 0.00486429
R56966 VCC.n5358 VCC.n5090 0.00486429
R56967 VCC.n5368 VCC.n5359 0.00486429
R56968 VCC.n5367 VCC.n5360 0.00486429
R56969 VCC.n5395 VCC.n5075 0.00486429
R56970 VCC.n5473 VCC.n5472 0.00486429
R56971 VCC.n5491 VCC.n5023 0.00486429
R56972 VCC.n5493 VCC.n5492 0.00486429
R56973 VCC.n5500 VCC.n5018 0.00486429
R56974 VCC.n5789 VCC.n5788 0.00486429
R56975 VCC.n5803 VCC.n5711 0.00486429
R56976 VCC.n5805 VCC.n5804 0.00486429
R56977 VCC.n5826 VCC.n5693 0.00486429
R56978 VCC.n5915 VCC.n5647 0.00486429
R56979 VCC.n5925 VCC.n5916 0.00486429
R56980 VCC.n5924 VCC.n5917 0.00486429
R56981 VCC.n5952 VCC.n5632 0.00486429
R56982 VCC.n6037 VCC.n6036 0.00486429
R56983 VCC.n6044 VCC.n5586 0.00486429
R56984 VCC.n6048 VCC.n6047 0.00486429
R56985 VCC.n6064 VCC.n5566 0.00486429
R56986 VCC.n6340 VCC.n6339 0.00486429
R56987 VCC.n6354 VCC.n6262 0.00486429
R56988 VCC.n6356 VCC.n6355 0.00486429
R56989 VCC.n6377 VCC.n6244 0.00486429
R56990 VCC.n6467 VCC.n6199 0.00486429
R56991 VCC.n6477 VCC.n6468 0.00486429
R56992 VCC.n6476 VCC.n6469 0.00486429
R56993 VCC.n6504 VCC.n6184 0.00486429
R56994 VCC.n6582 VCC.n6581 0.00486429
R56995 VCC.n6600 VCC.n6132 0.00486429
R56996 VCC.n6602 VCC.n6601 0.00486429
R56997 VCC.n6609 VCC.n6127 0.00486429
R56998 VCC.n6898 VCC.n6897 0.00486429
R56999 VCC.n6912 VCC.n6820 0.00486429
R57000 VCC.n6914 VCC.n6913 0.00486429
R57001 VCC.n6935 VCC.n6802 0.00486429
R57002 VCC.n7024 VCC.n6756 0.00486429
R57003 VCC.n7034 VCC.n7025 0.00486429
R57004 VCC.n7033 VCC.n7026 0.00486429
R57005 VCC.n7061 VCC.n6741 0.00486429
R57006 VCC.n7146 VCC.n7145 0.00486429
R57007 VCC.n7153 VCC.n6695 0.00486429
R57008 VCC.n7157 VCC.n7156 0.00486429
R57009 VCC.n7173 VCC.n6675 0.00486429
R57010 VCC.n7449 VCC.n7448 0.00486429
R57011 VCC.n7463 VCC.n7371 0.00486429
R57012 VCC.n7465 VCC.n7464 0.00486429
R57013 VCC.n7486 VCC.n7353 0.00486429
R57014 VCC.n7576 VCC.n7308 0.00486429
R57015 VCC.n7586 VCC.n7577 0.00486429
R57016 VCC.n7585 VCC.n7578 0.00486429
R57017 VCC.n7613 VCC.n7293 0.00486429
R57018 VCC.n7691 VCC.n7690 0.00486429
R57019 VCC.n7709 VCC.n7241 0.00486429
R57020 VCC.n7711 VCC.n7710 0.00486429
R57021 VCC.n7718 VCC.n7236 0.00486429
R57022 VCC.n8007 VCC.n8006 0.00486429
R57023 VCC.n8021 VCC.n7929 0.00486429
R57024 VCC.n8023 VCC.n8022 0.00486429
R57025 VCC.n8044 VCC.n7911 0.00486429
R57026 VCC.n8133 VCC.n7865 0.00486429
R57027 VCC.n8143 VCC.n8134 0.00486429
R57028 VCC.n8142 VCC.n8135 0.00486429
R57029 VCC.n8170 VCC.n7850 0.00486429
R57030 VCC.n8255 VCC.n8254 0.00486429
R57031 VCC.n8262 VCC.n7804 0.00486429
R57032 VCC.n8266 VCC.n8265 0.00486429
R57033 VCC.n8282 VCC.n7784 0.00486429
R57034 VCC.n8685 VCC.n8417 0.00486429
R57035 VCC.n8695 VCC.n8686 0.00486429
R57036 VCC.n8694 VCC.n8687 0.00486429
R57037 VCC.n8722 VCC.n8402 0.00486429
R57038 VCC.n8800 VCC.n8799 0.00486429
R57039 VCC.n8818 VCC.n8350 0.00486429
R57040 VCC.n8820 VCC.n8819 0.00486429
R57041 VCC.n8827 VCC.n8345 0.00486429
R57042 VCC.n9116 VCC.n9115 0.00486429
R57043 VCC.n9130 VCC.n9038 0.00486429
R57044 VCC.n9132 VCC.n9131 0.00486429
R57045 VCC.n9153 VCC.n9020 0.00486429
R57046 VCC.n9242 VCC.n8974 0.00486429
R57047 VCC.n9252 VCC.n9243 0.00486429
R57048 VCC.n9251 VCC.n9244 0.00486429
R57049 VCC.n9279 VCC.n8959 0.00486429
R57050 VCC.n9364 VCC.n9363 0.00486429
R57051 VCC.n9371 VCC.n8913 0.00486429
R57052 VCC.n9375 VCC.n9374 0.00486429
R57053 VCC.n9391 VCC.n8893 0.00486429
R57054 VCC.n9667 VCC.n9666 0.00486429
R57055 VCC.n9681 VCC.n9589 0.00486429
R57056 VCC.n9683 VCC.n9682 0.00486429
R57057 VCC.n9704 VCC.n9571 0.00486429
R57058 VCC.n9794 VCC.n9526 0.00486429
R57059 VCC.n9804 VCC.n9795 0.00486429
R57060 VCC.n9803 VCC.n9796 0.00486429
R57061 VCC.n9831 VCC.n9511 0.00486429
R57062 VCC.n9909 VCC.n9908 0.00486429
R57063 VCC.n9927 VCC.n9459 0.00486429
R57064 VCC.n9929 VCC.n9928 0.00486429
R57065 VCC.n9936 VCC.n9454 0.00486429
R57066 VCC.n10224 VCC.n10223 0.00486429
R57067 VCC.n10238 VCC.n10146 0.00486429
R57068 VCC.n10240 VCC.n10239 0.00486429
R57069 VCC.n10261 VCC.n10128 0.00486429
R57070 VCC.n10350 VCC.n10082 0.00486429
R57071 VCC.n10360 VCC.n10351 0.00486429
R57072 VCC.n10359 VCC.n10352 0.00486429
R57073 VCC.n10387 VCC.n10067 0.00486429
R57074 VCC.n10472 VCC.n10471 0.00486429
R57075 VCC.n10479 VCC.n10021 0.00486429
R57076 VCC.n10483 VCC.n10482 0.00486429
R57077 VCC.n10499 VCC.n10001 0.00486429
R57078 VCC.n10774 VCC.n10773 0.00486429
R57079 VCC.n10788 VCC.n10696 0.00486429
R57080 VCC.n10790 VCC.n10789 0.00486429
R57081 VCC.n10811 VCC.n10678 0.00486429
R57082 VCC.n10901 VCC.n10633 0.00486429
R57083 VCC.n10911 VCC.n10902 0.00486429
R57084 VCC.n10910 VCC.n10903 0.00486429
R57085 VCC.n10938 VCC.n10618 0.00486429
R57086 VCC.n11016 VCC.n11015 0.00486429
R57087 VCC.n11034 VCC.n10566 0.00486429
R57088 VCC.n11036 VCC.n11035 0.00486429
R57089 VCC.n11043 VCC.n10561 0.00486429
R57090 VCC.n11331 VCC.n11330 0.00486429
R57091 VCC.n11345 VCC.n11253 0.00486429
R57092 VCC.n11347 VCC.n11346 0.00486429
R57093 VCC.n11368 VCC.n11235 0.00486429
R57094 VCC.n11457 VCC.n11189 0.00486429
R57095 VCC.n11467 VCC.n11458 0.00486429
R57096 VCC.n11466 VCC.n11459 0.00486429
R57097 VCC.n11494 VCC.n11174 0.00486429
R57098 VCC.n11579 VCC.n11578 0.00486429
R57099 VCC.n11586 VCC.n11128 0.00486429
R57100 VCC.n11590 VCC.n11589 0.00486429
R57101 VCC.n11606 VCC.n11108 0.00486429
R57102 VCC.n11881 VCC.n11880 0.00486429
R57103 VCC.n11895 VCC.n11803 0.00486429
R57104 VCC.n11897 VCC.n11896 0.00486429
R57105 VCC.n11918 VCC.n11785 0.00486429
R57106 VCC.n12008 VCC.n11740 0.00486429
R57107 VCC.n12018 VCC.n12009 0.00486429
R57108 VCC.n12017 VCC.n12010 0.00486429
R57109 VCC.n12045 VCC.n11725 0.00486429
R57110 VCC.n12123 VCC.n12122 0.00486429
R57111 VCC.n12141 VCC.n11673 0.00486429
R57112 VCC.n12143 VCC.n12142 0.00486429
R57113 VCC.n12150 VCC.n11668 0.00486429
R57114 VCC.n12438 VCC.n12437 0.00486429
R57115 VCC.n12452 VCC.n12360 0.00486429
R57116 VCC.n12454 VCC.n12453 0.00486429
R57117 VCC.n12475 VCC.n12342 0.00486429
R57118 VCC.n12564 VCC.n12296 0.00486429
R57119 VCC.n12574 VCC.n12565 0.00486429
R57120 VCC.n12573 VCC.n12566 0.00486429
R57121 VCC.n12601 VCC.n12281 0.00486429
R57122 VCC.n12686 VCC.n12685 0.00486429
R57123 VCC.n12693 VCC.n12235 0.00486429
R57124 VCC.n12697 VCC.n12696 0.00486429
R57125 VCC.n12713 VCC.n12215 0.00486429
R57126 VCC.n12988 VCC.n12987 0.00486429
R57127 VCC.n13002 VCC.n12910 0.00486429
R57128 VCC.n13004 VCC.n13003 0.00486429
R57129 VCC.n13025 VCC.n12892 0.00486429
R57130 VCC.n13115 VCC.n12847 0.00486429
R57131 VCC.n13125 VCC.n13116 0.00486429
R57132 VCC.n13124 VCC.n13117 0.00486429
R57133 VCC.n13152 VCC.n12832 0.00486429
R57134 VCC.n13230 VCC.n13229 0.00486429
R57135 VCC.n13248 VCC.n12780 0.00486429
R57136 VCC.n13250 VCC.n13249 0.00486429
R57137 VCC.n13257 VCC.n12775 0.00486429
R57138 VCC.n13545 VCC.n13544 0.00486429
R57139 VCC.n13559 VCC.n13467 0.00486429
R57140 VCC.n13561 VCC.n13560 0.00486429
R57141 VCC.n13582 VCC.n13449 0.00486429
R57142 VCC.n13671 VCC.n13403 0.00486429
R57143 VCC.n13681 VCC.n13672 0.00486429
R57144 VCC.n13680 VCC.n13673 0.00486429
R57145 VCC.n13708 VCC.n13388 0.00486429
R57146 VCC.n13793 VCC.n13792 0.00486429
R57147 VCC.n13800 VCC.n13342 0.00486429
R57148 VCC.n13804 VCC.n13803 0.00486429
R57149 VCC.n13820 VCC.n13322 0.00486429
R57150 VCC.n14095 VCC.n14094 0.00486429
R57151 VCC.n14109 VCC.n14017 0.00486429
R57152 VCC.n14111 VCC.n14110 0.00486429
R57153 VCC.n14132 VCC.n13999 0.00486429
R57154 VCC.n14222 VCC.n13954 0.00486429
R57155 VCC.n14232 VCC.n14223 0.00486429
R57156 VCC.n14231 VCC.n14224 0.00486429
R57157 VCC.n14259 VCC.n13939 0.00486429
R57158 VCC.n14337 VCC.n14336 0.00486429
R57159 VCC.n14355 VCC.n13887 0.00486429
R57160 VCC.n14357 VCC.n14356 0.00486429
R57161 VCC.n14364 VCC.n13882 0.00486429
R57162 VCC.n14652 VCC.n14651 0.00486429
R57163 VCC.n14666 VCC.n14574 0.00486429
R57164 VCC.n14668 VCC.n14667 0.00486429
R57165 VCC.n14689 VCC.n14556 0.00486429
R57166 VCC.n14778 VCC.n14510 0.00486429
R57167 VCC.n14788 VCC.n14779 0.00486429
R57168 VCC.n14787 VCC.n14780 0.00486429
R57169 VCC.n14815 VCC.n14495 0.00486429
R57170 VCC.n14900 VCC.n14899 0.00486429
R57171 VCC.n14907 VCC.n14449 0.00486429
R57172 VCC.n14911 VCC.n14910 0.00486429
R57173 VCC.n14927 VCC.n14429 0.00486429
R57174 VCC.n15202 VCC.n15201 0.00486429
R57175 VCC.n15216 VCC.n15124 0.00486429
R57176 VCC.n15218 VCC.n15217 0.00486429
R57177 VCC.n15239 VCC.n15106 0.00486429
R57178 VCC.n15329 VCC.n15061 0.00486429
R57179 VCC.n15339 VCC.n15330 0.00486429
R57180 VCC.n15338 VCC.n15331 0.00486429
R57181 VCC.n15366 VCC.n15046 0.00486429
R57182 VCC.n15444 VCC.n15443 0.00486429
R57183 VCC.n15462 VCC.n14994 0.00486429
R57184 VCC.n15464 VCC.n15463 0.00486429
R57185 VCC.n15471 VCC.n14989 0.00486429
R57186 VCC.n15759 VCC.n15758 0.00486429
R57187 VCC.n15773 VCC.n15681 0.00486429
R57188 VCC.n15775 VCC.n15774 0.00486429
R57189 VCC.n15796 VCC.n15663 0.00486429
R57190 VCC.n15885 VCC.n15617 0.00486429
R57191 VCC.n15895 VCC.n15886 0.00486429
R57192 VCC.n15894 VCC.n15887 0.00486429
R57193 VCC.n15922 VCC.n15602 0.00486429
R57194 VCC.n16007 VCC.n16006 0.00486429
R57195 VCC.n16014 VCC.n15556 0.00486429
R57196 VCC.n16018 VCC.n16017 0.00486429
R57197 VCC.n16034 VCC.n15536 0.00486429
R57198 VCC.n16309 VCC.n16308 0.00486429
R57199 VCC.n16323 VCC.n16231 0.00486429
R57200 VCC.n16325 VCC.n16324 0.00486429
R57201 VCC.n16346 VCC.n16213 0.00486429
R57202 VCC.n16436 VCC.n16168 0.00486429
R57203 VCC.n16446 VCC.n16437 0.00486429
R57204 VCC.n16445 VCC.n16438 0.00486429
R57205 VCC.n16473 VCC.n16153 0.00486429
R57206 VCC.n16551 VCC.n16550 0.00486429
R57207 VCC.n16569 VCC.n16101 0.00486429
R57208 VCC.n16571 VCC.n16570 0.00486429
R57209 VCC.n16578 VCC.n16096 0.00486429
R57210 VCC.n16866 VCC.n16865 0.00486429
R57211 VCC.n16880 VCC.n16788 0.00486429
R57212 VCC.n16882 VCC.n16881 0.00486429
R57213 VCC.n16903 VCC.n16770 0.00486429
R57214 VCC.n16992 VCC.n16724 0.00486429
R57215 VCC.n17002 VCC.n16993 0.00486429
R57216 VCC.n17001 VCC.n16994 0.00486429
R57217 VCC.n17029 VCC.n16709 0.00486429
R57218 VCC.n17114 VCC.n17113 0.00486429
R57219 VCC.n17121 VCC.n16663 0.00486429
R57220 VCC.n17125 VCC.n17124 0.00486429
R57221 VCC.n17141 VCC.n16643 0.00486429
R57222 VCC.n17356 VCC.n17275 0.00486429
R57223 VCC.n17366 VCC.n17357 0.00486429
R57224 VCC.n17365 VCC.n17358 0.00486429
R57225 VCC.n17393 VCC.n17260 0.00486429
R57226 VCC.n17471 VCC.n17470 0.00486429
R57227 VCC.n17489 VCC.n17208 0.00486429
R57228 VCC.n17491 VCC.n17490 0.00486429
R57229 VCC.n17498 VCC.n17203 0.00486429
R57230 VCC.n8558 VCC.n8557 0.00483333
R57231 VCC.n8572 VCC.n8480 0.00483333
R57232 VCC.n8574 VCC.n8573 0.00483333
R57233 VCC.n8595 VCC.n8462 0.00483333
R57234 VCC.n203 VCC.n202 0.00407143
R57235 VCC.n250 VCC.n168 0.00407143
R57236 VCC.n255 VCC.n251 0.00407143
R57237 VCC.n305 VCC.n134 0.00407143
R57238 VCC.n256 VCC.n166 0.00407143
R57239 VCC.n377 VCC.n96 0.00407143
R57240 VCC.n434 VCC.n76 0.00407143
R57241 VCC.n378 VCC.n375 0.00407143
R57242 VCC.n755 VCC.n754 0.00407143
R57243 VCC.n802 VCC.n720 0.00407143
R57244 VCC.n807 VCC.n803 0.00407143
R57245 VCC.n857 VCC.n686 0.00407143
R57246 VCC.n808 VCC.n718 0.00407143
R57247 VCC.n929 VCC.n648 0.00407143
R57248 VCC.n986 VCC.n628 0.00407143
R57249 VCC.n930 VCC.n927 0.00407143
R57250 VCC.n1486 VCC.n1205 0.00407143
R57251 VCC.n1544 VCC.n1185 0.00407143
R57252 VCC.n1487 VCC.n1484 0.00407143
R57253 VCC.n1313 VCC.n1312 0.00407143
R57254 VCC.n1360 VCC.n1278 0.00407143
R57255 VCC.n1365 VCC.n1361 0.00407143
R57256 VCC.n1415 VCC.n1244 0.00407143
R57257 VCC.n1366 VCC.n1276 0.00407143
R57258 VCC.n1864 VCC.n1863 0.00407143
R57259 VCC.n1911 VCC.n1829 0.00407143
R57260 VCC.n1916 VCC.n1912 0.00407143
R57261 VCC.n1966 VCC.n1795 0.00407143
R57262 VCC.n1917 VCC.n1827 0.00407143
R57263 VCC.n2038 VCC.n1757 0.00407143
R57264 VCC.n2095 VCC.n1737 0.00407143
R57265 VCC.n2039 VCC.n2036 0.00407143
R57266 VCC.n2595 VCC.n2314 0.00407143
R57267 VCC.n2653 VCC.n2294 0.00407143
R57268 VCC.n2596 VCC.n2593 0.00407143
R57269 VCC.n2422 VCC.n2421 0.00407143
R57270 VCC.n2469 VCC.n2387 0.00407143
R57271 VCC.n2474 VCC.n2470 0.00407143
R57272 VCC.n2524 VCC.n2353 0.00407143
R57273 VCC.n2475 VCC.n2385 0.00407143
R57274 VCC.n2973 VCC.n2972 0.00407143
R57275 VCC.n3020 VCC.n2938 0.00407143
R57276 VCC.n3025 VCC.n3021 0.00407143
R57277 VCC.n3075 VCC.n2904 0.00407143
R57278 VCC.n3026 VCC.n2936 0.00407143
R57279 VCC.n3147 VCC.n2866 0.00407143
R57280 VCC.n3204 VCC.n2846 0.00407143
R57281 VCC.n3148 VCC.n3145 0.00407143
R57282 VCC.n3704 VCC.n3423 0.00407143
R57283 VCC.n3762 VCC.n3403 0.00407143
R57284 VCC.n3705 VCC.n3702 0.00407143
R57285 VCC.n3531 VCC.n3530 0.00407143
R57286 VCC.n3578 VCC.n3496 0.00407143
R57287 VCC.n3583 VCC.n3579 0.00407143
R57288 VCC.n3633 VCC.n3462 0.00407143
R57289 VCC.n3584 VCC.n3494 0.00407143
R57290 VCC.n4082 VCC.n4081 0.00407143
R57291 VCC.n4129 VCC.n4047 0.00407143
R57292 VCC.n4134 VCC.n4130 0.00407143
R57293 VCC.n4184 VCC.n4013 0.00407143
R57294 VCC.n4135 VCC.n4045 0.00407143
R57295 VCC.n4256 VCC.n3975 0.00407143
R57296 VCC.n4313 VCC.n3955 0.00407143
R57297 VCC.n4257 VCC.n4254 0.00407143
R57298 VCC.n4813 VCC.n4532 0.00407143
R57299 VCC.n4871 VCC.n4512 0.00407143
R57300 VCC.n4814 VCC.n4811 0.00407143
R57301 VCC.n4640 VCC.n4639 0.00407143
R57302 VCC.n4687 VCC.n4605 0.00407143
R57303 VCC.n4692 VCC.n4688 0.00407143
R57304 VCC.n4742 VCC.n4571 0.00407143
R57305 VCC.n4693 VCC.n4603 0.00407143
R57306 VCC.n5191 VCC.n5190 0.00407143
R57307 VCC.n5238 VCC.n5156 0.00407143
R57308 VCC.n5243 VCC.n5239 0.00407143
R57309 VCC.n5293 VCC.n5122 0.00407143
R57310 VCC.n5244 VCC.n5154 0.00407143
R57311 VCC.n5365 VCC.n5084 0.00407143
R57312 VCC.n5422 VCC.n5064 0.00407143
R57313 VCC.n5366 VCC.n5363 0.00407143
R57314 VCC.n5922 VCC.n5641 0.00407143
R57315 VCC.n5980 VCC.n5621 0.00407143
R57316 VCC.n5923 VCC.n5920 0.00407143
R57317 VCC.n5749 VCC.n5748 0.00407143
R57318 VCC.n5796 VCC.n5714 0.00407143
R57319 VCC.n5801 VCC.n5797 0.00407143
R57320 VCC.n5851 VCC.n5680 0.00407143
R57321 VCC.n5802 VCC.n5712 0.00407143
R57322 VCC.n6300 VCC.n6299 0.00407143
R57323 VCC.n6347 VCC.n6265 0.00407143
R57324 VCC.n6352 VCC.n6348 0.00407143
R57325 VCC.n6402 VCC.n6231 0.00407143
R57326 VCC.n6353 VCC.n6263 0.00407143
R57327 VCC.n6474 VCC.n6193 0.00407143
R57328 VCC.n6531 VCC.n6173 0.00407143
R57329 VCC.n6475 VCC.n6472 0.00407143
R57330 VCC.n7031 VCC.n6750 0.00407143
R57331 VCC.n7089 VCC.n6730 0.00407143
R57332 VCC.n7032 VCC.n7029 0.00407143
R57333 VCC.n6858 VCC.n6857 0.00407143
R57334 VCC.n6905 VCC.n6823 0.00407143
R57335 VCC.n6910 VCC.n6906 0.00407143
R57336 VCC.n6960 VCC.n6789 0.00407143
R57337 VCC.n6911 VCC.n6821 0.00407143
R57338 VCC.n7409 VCC.n7408 0.00407143
R57339 VCC.n7456 VCC.n7374 0.00407143
R57340 VCC.n7461 VCC.n7457 0.00407143
R57341 VCC.n7511 VCC.n7340 0.00407143
R57342 VCC.n7462 VCC.n7372 0.00407143
R57343 VCC.n7583 VCC.n7302 0.00407143
R57344 VCC.n7640 VCC.n7282 0.00407143
R57345 VCC.n7584 VCC.n7581 0.00407143
R57346 VCC.n8140 VCC.n7859 0.00407143
R57347 VCC.n8198 VCC.n7839 0.00407143
R57348 VCC.n8141 VCC.n8138 0.00407143
R57349 VCC.n7967 VCC.n7966 0.00407143
R57350 VCC.n8014 VCC.n7932 0.00407143
R57351 VCC.n8019 VCC.n8015 0.00407143
R57352 VCC.n8069 VCC.n7898 0.00407143
R57353 VCC.n8020 VCC.n7930 0.00407143
R57354 VCC.n8692 VCC.n8411 0.00407143
R57355 VCC.n8749 VCC.n8391 0.00407143
R57356 VCC.n8693 VCC.n8690 0.00407143
R57357 VCC.n8518 VCC.n8517 0.00407143
R57358 VCC.n8565 VCC.n8483 0.00407143
R57359 VCC.n8570 VCC.n8566 0.00407143
R57360 VCC.n8620 VCC.n8449 0.00407143
R57361 VCC.n8571 VCC.n8481 0.00407143
R57362 VCC.n9249 VCC.n8968 0.00407143
R57363 VCC.n9307 VCC.n8948 0.00407143
R57364 VCC.n9250 VCC.n9247 0.00407143
R57365 VCC.n9076 VCC.n9075 0.00407143
R57366 VCC.n9123 VCC.n9041 0.00407143
R57367 VCC.n9128 VCC.n9124 0.00407143
R57368 VCC.n9178 VCC.n9007 0.00407143
R57369 VCC.n9129 VCC.n9039 0.00407143
R57370 VCC.n9627 VCC.n9626 0.00407143
R57371 VCC.n9674 VCC.n9592 0.00407143
R57372 VCC.n9679 VCC.n9675 0.00407143
R57373 VCC.n9729 VCC.n9558 0.00407143
R57374 VCC.n9680 VCC.n9590 0.00407143
R57375 VCC.n9801 VCC.n9520 0.00407143
R57376 VCC.n9858 VCC.n9500 0.00407143
R57377 VCC.n9802 VCC.n9799 0.00407143
R57378 VCC.n10357 VCC.n10076 0.00407143
R57379 VCC.n10415 VCC.n10056 0.00407143
R57380 VCC.n10358 VCC.n10355 0.00407143
R57381 VCC.n10184 VCC.n10183 0.00407143
R57382 VCC.n10231 VCC.n10149 0.00407143
R57383 VCC.n10236 VCC.n10232 0.00407143
R57384 VCC.n10286 VCC.n10115 0.00407143
R57385 VCC.n10237 VCC.n10147 0.00407143
R57386 VCC.n10734 VCC.n10733 0.00407143
R57387 VCC.n10781 VCC.n10699 0.00407143
R57388 VCC.n10786 VCC.n10782 0.00407143
R57389 VCC.n10836 VCC.n10665 0.00407143
R57390 VCC.n10787 VCC.n10697 0.00407143
R57391 VCC.n10908 VCC.n10627 0.00407143
R57392 VCC.n10965 VCC.n10607 0.00407143
R57393 VCC.n10909 VCC.n10906 0.00407143
R57394 VCC.n11464 VCC.n11183 0.00407143
R57395 VCC.n11522 VCC.n11163 0.00407143
R57396 VCC.n11465 VCC.n11462 0.00407143
R57397 VCC.n11291 VCC.n11290 0.00407143
R57398 VCC.n11338 VCC.n11256 0.00407143
R57399 VCC.n11343 VCC.n11339 0.00407143
R57400 VCC.n11393 VCC.n11222 0.00407143
R57401 VCC.n11344 VCC.n11254 0.00407143
R57402 VCC.n11841 VCC.n11840 0.00407143
R57403 VCC.n11888 VCC.n11806 0.00407143
R57404 VCC.n11893 VCC.n11889 0.00407143
R57405 VCC.n11943 VCC.n11772 0.00407143
R57406 VCC.n11894 VCC.n11804 0.00407143
R57407 VCC.n12015 VCC.n11734 0.00407143
R57408 VCC.n12072 VCC.n11714 0.00407143
R57409 VCC.n12016 VCC.n12013 0.00407143
R57410 VCC.n12571 VCC.n12290 0.00407143
R57411 VCC.n12629 VCC.n12270 0.00407143
R57412 VCC.n12572 VCC.n12569 0.00407143
R57413 VCC.n12398 VCC.n12397 0.00407143
R57414 VCC.n12445 VCC.n12363 0.00407143
R57415 VCC.n12450 VCC.n12446 0.00407143
R57416 VCC.n12500 VCC.n12329 0.00407143
R57417 VCC.n12451 VCC.n12361 0.00407143
R57418 VCC.n12948 VCC.n12947 0.00407143
R57419 VCC.n12995 VCC.n12913 0.00407143
R57420 VCC.n13000 VCC.n12996 0.00407143
R57421 VCC.n13050 VCC.n12879 0.00407143
R57422 VCC.n13001 VCC.n12911 0.00407143
R57423 VCC.n13122 VCC.n12841 0.00407143
R57424 VCC.n13179 VCC.n12821 0.00407143
R57425 VCC.n13123 VCC.n13120 0.00407143
R57426 VCC.n13678 VCC.n13397 0.00407143
R57427 VCC.n13736 VCC.n13377 0.00407143
R57428 VCC.n13679 VCC.n13676 0.00407143
R57429 VCC.n13505 VCC.n13504 0.00407143
R57430 VCC.n13552 VCC.n13470 0.00407143
R57431 VCC.n13557 VCC.n13553 0.00407143
R57432 VCC.n13607 VCC.n13436 0.00407143
R57433 VCC.n13558 VCC.n13468 0.00407143
R57434 VCC.n14055 VCC.n14054 0.00407143
R57435 VCC.n14102 VCC.n14020 0.00407143
R57436 VCC.n14107 VCC.n14103 0.00407143
R57437 VCC.n14157 VCC.n13986 0.00407143
R57438 VCC.n14108 VCC.n14018 0.00407143
R57439 VCC.n14229 VCC.n13948 0.00407143
R57440 VCC.n14286 VCC.n13928 0.00407143
R57441 VCC.n14230 VCC.n14227 0.00407143
R57442 VCC.n14785 VCC.n14504 0.00407143
R57443 VCC.n14843 VCC.n14484 0.00407143
R57444 VCC.n14786 VCC.n14783 0.00407143
R57445 VCC.n14612 VCC.n14611 0.00407143
R57446 VCC.n14659 VCC.n14577 0.00407143
R57447 VCC.n14664 VCC.n14660 0.00407143
R57448 VCC.n14714 VCC.n14543 0.00407143
R57449 VCC.n14665 VCC.n14575 0.00407143
R57450 VCC.n15162 VCC.n15161 0.00407143
R57451 VCC.n15209 VCC.n15127 0.00407143
R57452 VCC.n15214 VCC.n15210 0.00407143
R57453 VCC.n15264 VCC.n15093 0.00407143
R57454 VCC.n15215 VCC.n15125 0.00407143
R57455 VCC.n15336 VCC.n15055 0.00407143
R57456 VCC.n15393 VCC.n15035 0.00407143
R57457 VCC.n15337 VCC.n15334 0.00407143
R57458 VCC.n15892 VCC.n15611 0.00407143
R57459 VCC.n15950 VCC.n15591 0.00407143
R57460 VCC.n15893 VCC.n15890 0.00407143
R57461 VCC.n15719 VCC.n15718 0.00407143
R57462 VCC.n15766 VCC.n15684 0.00407143
R57463 VCC.n15771 VCC.n15767 0.00407143
R57464 VCC.n15821 VCC.n15650 0.00407143
R57465 VCC.n15772 VCC.n15682 0.00407143
R57466 VCC.n16269 VCC.n16268 0.00407143
R57467 VCC.n16316 VCC.n16234 0.00407143
R57468 VCC.n16321 VCC.n16317 0.00407143
R57469 VCC.n16371 VCC.n16200 0.00407143
R57470 VCC.n16322 VCC.n16232 0.00407143
R57471 VCC.n16443 VCC.n16162 0.00407143
R57472 VCC.n16500 VCC.n16142 0.00407143
R57473 VCC.n16444 VCC.n16441 0.00407143
R57474 VCC.n16999 VCC.n16718 0.00407143
R57475 VCC.n17057 VCC.n16698 0.00407143
R57476 VCC.n17000 VCC.n16997 0.00407143
R57477 VCC.n16826 VCC.n16825 0.00407143
R57478 VCC.n16873 VCC.n16791 0.00407143
R57479 VCC.n16878 VCC.n16874 0.00407143
R57480 VCC.n16928 VCC.n16757 0.00407143
R57481 VCC.n16879 VCC.n16789 0.00407143
R57482 VCC.n17363 VCC.n17269 0.00407143
R57483 VCC.n17420 VCC.n17249 0.00407143
R57484 VCC.n17364 VCC.n17361 0.00407143
R57485 VCC.n243 VCC.n165 0.00318571
R57486 VCC.n259 VCC.n147 0.00318571
R57487 VCC.n371 VCC.n370 0.00318571
R57488 VCC.n372 VCC.n87 0.00318571
R57489 VCC.n484 VCC.n35 0.00318571
R57490 VCC.n505 VCC.n30 0.00318571
R57491 VCC.n795 VCC.n717 0.00318571
R57492 VCC.n811 VCC.n699 0.00318571
R57493 VCC.n923 VCC.n922 0.00318571
R57494 VCC.n924 VCC.n639 0.00318571
R57495 VCC.n1036 VCC.n587 0.00318571
R57496 VCC.n1057 VCC.n582 0.00318571
R57497 VCC.n1353 VCC.n1275 0.00318571
R57498 VCC.n1369 VCC.n1257 0.00318571
R57499 VCC.n1480 VCC.n1479 0.00318571
R57500 VCC.n1481 VCC.n1196 0.00318571
R57501 VCC.n1601 VCC.n1150 0.00318571
R57502 VCC.n1611 VCC.n1130 0.00318571
R57503 VCC.n1904 VCC.n1826 0.00318571
R57504 VCC.n1920 VCC.n1808 0.00318571
R57505 VCC.n2032 VCC.n2031 0.00318571
R57506 VCC.n2033 VCC.n1748 0.00318571
R57507 VCC.n2145 VCC.n1696 0.00318571
R57508 VCC.n2166 VCC.n1691 0.00318571
R57509 VCC.n2462 VCC.n2384 0.00318571
R57510 VCC.n2478 VCC.n2366 0.00318571
R57511 VCC.n2589 VCC.n2588 0.00318571
R57512 VCC.n2590 VCC.n2305 0.00318571
R57513 VCC.n2710 VCC.n2259 0.00318571
R57514 VCC.n2720 VCC.n2239 0.00318571
R57515 VCC.n3013 VCC.n2935 0.00318571
R57516 VCC.n3029 VCC.n2917 0.00318571
R57517 VCC.n3141 VCC.n3140 0.00318571
R57518 VCC.n3142 VCC.n2857 0.00318571
R57519 VCC.n3254 VCC.n2805 0.00318571
R57520 VCC.n3275 VCC.n2800 0.00318571
R57521 VCC.n3571 VCC.n3493 0.00318571
R57522 VCC.n3587 VCC.n3475 0.00318571
R57523 VCC.n3698 VCC.n3697 0.00318571
R57524 VCC.n3699 VCC.n3414 0.00318571
R57525 VCC.n3819 VCC.n3368 0.00318571
R57526 VCC.n3829 VCC.n3348 0.00318571
R57527 VCC.n4122 VCC.n4044 0.00318571
R57528 VCC.n4138 VCC.n4026 0.00318571
R57529 VCC.n4250 VCC.n4249 0.00318571
R57530 VCC.n4251 VCC.n3966 0.00318571
R57531 VCC.n4363 VCC.n3914 0.00318571
R57532 VCC.n4384 VCC.n3909 0.00318571
R57533 VCC.n4680 VCC.n4602 0.00318571
R57534 VCC.n4696 VCC.n4584 0.00318571
R57535 VCC.n4807 VCC.n4806 0.00318571
R57536 VCC.n4808 VCC.n4523 0.00318571
R57537 VCC.n4928 VCC.n4477 0.00318571
R57538 VCC.n4938 VCC.n4457 0.00318571
R57539 VCC.n5231 VCC.n5153 0.00318571
R57540 VCC.n5247 VCC.n5135 0.00318571
R57541 VCC.n5359 VCC.n5358 0.00318571
R57542 VCC.n5360 VCC.n5075 0.00318571
R57543 VCC.n5472 VCC.n5023 0.00318571
R57544 VCC.n5493 VCC.n5018 0.00318571
R57545 VCC.n5789 VCC.n5711 0.00318571
R57546 VCC.n5805 VCC.n5693 0.00318571
R57547 VCC.n5916 VCC.n5915 0.00318571
R57548 VCC.n5917 VCC.n5632 0.00318571
R57549 VCC.n6037 VCC.n5586 0.00318571
R57550 VCC.n6047 VCC.n5566 0.00318571
R57551 VCC.n6340 VCC.n6262 0.00318571
R57552 VCC.n6356 VCC.n6244 0.00318571
R57553 VCC.n6468 VCC.n6467 0.00318571
R57554 VCC.n6469 VCC.n6184 0.00318571
R57555 VCC.n6581 VCC.n6132 0.00318571
R57556 VCC.n6602 VCC.n6127 0.00318571
R57557 VCC.n6898 VCC.n6820 0.00318571
R57558 VCC.n6914 VCC.n6802 0.00318571
R57559 VCC.n7025 VCC.n7024 0.00318571
R57560 VCC.n7026 VCC.n6741 0.00318571
R57561 VCC.n7146 VCC.n6695 0.00318571
R57562 VCC.n7156 VCC.n6675 0.00318571
R57563 VCC.n7449 VCC.n7371 0.00318571
R57564 VCC.n7465 VCC.n7353 0.00318571
R57565 VCC.n7577 VCC.n7576 0.00318571
R57566 VCC.n7578 VCC.n7293 0.00318571
R57567 VCC.n7690 VCC.n7241 0.00318571
R57568 VCC.n7711 VCC.n7236 0.00318571
R57569 VCC.n8007 VCC.n7929 0.00318571
R57570 VCC.n8023 VCC.n7911 0.00318571
R57571 VCC.n8134 VCC.n8133 0.00318571
R57572 VCC.n8135 VCC.n7850 0.00318571
R57573 VCC.n8255 VCC.n7804 0.00318571
R57574 VCC.n8265 VCC.n7784 0.00318571
R57575 VCC.n8686 VCC.n8685 0.00318571
R57576 VCC.n8687 VCC.n8402 0.00318571
R57577 VCC.n8799 VCC.n8350 0.00318571
R57578 VCC.n8820 VCC.n8345 0.00318571
R57579 VCC.n9116 VCC.n9038 0.00318571
R57580 VCC.n9132 VCC.n9020 0.00318571
R57581 VCC.n9243 VCC.n9242 0.00318571
R57582 VCC.n9244 VCC.n8959 0.00318571
R57583 VCC.n9364 VCC.n8913 0.00318571
R57584 VCC.n9374 VCC.n8893 0.00318571
R57585 VCC.n9667 VCC.n9589 0.00318571
R57586 VCC.n9683 VCC.n9571 0.00318571
R57587 VCC.n9795 VCC.n9794 0.00318571
R57588 VCC.n9796 VCC.n9511 0.00318571
R57589 VCC.n9908 VCC.n9459 0.00318571
R57590 VCC.n9929 VCC.n9454 0.00318571
R57591 VCC.n10224 VCC.n10146 0.00318571
R57592 VCC.n10240 VCC.n10128 0.00318571
R57593 VCC.n10351 VCC.n10350 0.00318571
R57594 VCC.n10352 VCC.n10067 0.00318571
R57595 VCC.n10472 VCC.n10021 0.00318571
R57596 VCC.n10482 VCC.n10001 0.00318571
R57597 VCC.n10774 VCC.n10696 0.00318571
R57598 VCC.n10790 VCC.n10678 0.00318571
R57599 VCC.n10902 VCC.n10901 0.00318571
R57600 VCC.n10903 VCC.n10618 0.00318571
R57601 VCC.n11015 VCC.n10566 0.00318571
R57602 VCC.n11036 VCC.n10561 0.00318571
R57603 VCC.n11331 VCC.n11253 0.00318571
R57604 VCC.n11347 VCC.n11235 0.00318571
R57605 VCC.n11458 VCC.n11457 0.00318571
R57606 VCC.n11459 VCC.n11174 0.00318571
R57607 VCC.n11579 VCC.n11128 0.00318571
R57608 VCC.n11589 VCC.n11108 0.00318571
R57609 VCC.n11881 VCC.n11803 0.00318571
R57610 VCC.n11897 VCC.n11785 0.00318571
R57611 VCC.n12009 VCC.n12008 0.00318571
R57612 VCC.n12010 VCC.n11725 0.00318571
R57613 VCC.n12122 VCC.n11673 0.00318571
R57614 VCC.n12143 VCC.n11668 0.00318571
R57615 VCC.n12438 VCC.n12360 0.00318571
R57616 VCC.n12454 VCC.n12342 0.00318571
R57617 VCC.n12565 VCC.n12564 0.00318571
R57618 VCC.n12566 VCC.n12281 0.00318571
R57619 VCC.n12686 VCC.n12235 0.00318571
R57620 VCC.n12696 VCC.n12215 0.00318571
R57621 VCC.n12988 VCC.n12910 0.00318571
R57622 VCC.n13004 VCC.n12892 0.00318571
R57623 VCC.n13116 VCC.n13115 0.00318571
R57624 VCC.n13117 VCC.n12832 0.00318571
R57625 VCC.n13229 VCC.n12780 0.00318571
R57626 VCC.n13250 VCC.n12775 0.00318571
R57627 VCC.n13545 VCC.n13467 0.00318571
R57628 VCC.n13561 VCC.n13449 0.00318571
R57629 VCC.n13672 VCC.n13671 0.00318571
R57630 VCC.n13673 VCC.n13388 0.00318571
R57631 VCC.n13793 VCC.n13342 0.00318571
R57632 VCC.n13803 VCC.n13322 0.00318571
R57633 VCC.n14095 VCC.n14017 0.00318571
R57634 VCC.n14111 VCC.n13999 0.00318571
R57635 VCC.n14223 VCC.n14222 0.00318571
R57636 VCC.n14224 VCC.n13939 0.00318571
R57637 VCC.n14336 VCC.n13887 0.00318571
R57638 VCC.n14357 VCC.n13882 0.00318571
R57639 VCC.n14652 VCC.n14574 0.00318571
R57640 VCC.n14668 VCC.n14556 0.00318571
R57641 VCC.n14779 VCC.n14778 0.00318571
R57642 VCC.n14780 VCC.n14495 0.00318571
R57643 VCC.n14900 VCC.n14449 0.00318571
R57644 VCC.n14910 VCC.n14429 0.00318571
R57645 VCC.n15202 VCC.n15124 0.00318571
R57646 VCC.n15218 VCC.n15106 0.00318571
R57647 VCC.n15330 VCC.n15329 0.00318571
R57648 VCC.n15331 VCC.n15046 0.00318571
R57649 VCC.n15443 VCC.n14994 0.00318571
R57650 VCC.n15464 VCC.n14989 0.00318571
R57651 VCC.n15759 VCC.n15681 0.00318571
R57652 VCC.n15775 VCC.n15663 0.00318571
R57653 VCC.n15886 VCC.n15885 0.00318571
R57654 VCC.n15887 VCC.n15602 0.00318571
R57655 VCC.n16007 VCC.n15556 0.00318571
R57656 VCC.n16017 VCC.n15536 0.00318571
R57657 VCC.n16309 VCC.n16231 0.00318571
R57658 VCC.n16325 VCC.n16213 0.00318571
R57659 VCC.n16437 VCC.n16436 0.00318571
R57660 VCC.n16438 VCC.n16153 0.00318571
R57661 VCC.n16550 VCC.n16101 0.00318571
R57662 VCC.n16571 VCC.n16096 0.00318571
R57663 VCC.n16866 VCC.n16788 0.00318571
R57664 VCC.n16882 VCC.n16770 0.00318571
R57665 VCC.n16993 VCC.n16992 0.00318571
R57666 VCC.n16994 VCC.n16709 0.00318571
R57667 VCC.n17114 VCC.n16663 0.00318571
R57668 VCC.n17124 VCC.n16643 0.00318571
R57669 VCC.n17357 VCC.n17356 0.00318571
R57670 VCC.n17358 VCC.n17260 0.00318571
R57671 VCC.n17470 VCC.n17208 0.00318571
R57672 VCC.n17491 VCC.n17203 0.00318571
R57673 VCC.n220 VCC.n185 0.00317857
R57674 VCC.n262 VCC.n157 0.00317857
R57675 VCC.n305 VCC.n304 0.00317857
R57676 VCC.n310 VCC.n129 0.00317857
R57677 VCC.n216 VCC.n190 0.00317857
R57678 VCC.n219 VCC.n186 0.00317857
R57679 VCC.n261 VCC.n163 0.00317857
R57680 VCC.n306 VCC.n133 0.00317857
R57681 VCC.n309 VCC.n130 0.00317857
R57682 VCC.n332 VCC.n125 0.00317857
R57683 VCC.n343 VCC.n116 0.00317857
R57684 VCC.n343 VCC.n342 0.00317857
R57685 VCC.n105 VCC.n98 0.00317857
R57686 VCC.n383 VCC.n99 0.00317857
R57687 VCC.n389 VCC.n388 0.00317857
R57688 VCC.n440 VCC.n73 0.00317857
R57689 VCC.n440 VCC.n439 0.00317857
R57690 VCC.n445 VCC.n68 0.00317857
R57691 VCC.n319 VCC.n318 0.00317857
R57692 VCC.n344 VCC.n115 0.00317857
R57693 VCC.n382 VCC.n381 0.00317857
R57694 VCC.n441 VCC.n72 0.00317857
R57695 VCC.n444 VCC.n69 0.00317857
R57696 VCC.n458 VCC.n457 0.00317857
R57697 VCC.n463 VCC.n59 0.00317857
R57698 VCC.n508 VCC.n32 0.00317857
R57699 VCC.n517 VCC.n516 0.00317857
R57700 VCC.n534 VCC.n533 0.00317857
R57701 VCC.n12 VCC.n11 0.00317857
R57702 VCC.n12 VCC.n2 0.00317857
R57703 VCC.n459 VCC.n64 0.00317857
R57704 VCC.n465 VCC.n464 0.00317857
R57705 VCC.n507 VCC.n33 0.00317857
R57706 VCC.n535 VCC.n15 0.00317857
R57707 VCC.n539 VCC.n538 0.00317857
R57708 VCC.n772 VCC.n737 0.00317857
R57709 VCC.n814 VCC.n709 0.00317857
R57710 VCC.n857 VCC.n856 0.00317857
R57711 VCC.n862 VCC.n681 0.00317857
R57712 VCC.n768 VCC.n742 0.00317857
R57713 VCC.n771 VCC.n738 0.00317857
R57714 VCC.n813 VCC.n715 0.00317857
R57715 VCC.n858 VCC.n685 0.00317857
R57716 VCC.n861 VCC.n682 0.00317857
R57717 VCC.n884 VCC.n677 0.00317857
R57718 VCC.n895 VCC.n668 0.00317857
R57719 VCC.n895 VCC.n894 0.00317857
R57720 VCC.n657 VCC.n650 0.00317857
R57721 VCC.n935 VCC.n651 0.00317857
R57722 VCC.n941 VCC.n940 0.00317857
R57723 VCC.n992 VCC.n625 0.00317857
R57724 VCC.n992 VCC.n991 0.00317857
R57725 VCC.n997 VCC.n620 0.00317857
R57726 VCC.n871 VCC.n870 0.00317857
R57727 VCC.n896 VCC.n667 0.00317857
R57728 VCC.n934 VCC.n933 0.00317857
R57729 VCC.n993 VCC.n624 0.00317857
R57730 VCC.n996 VCC.n621 0.00317857
R57731 VCC.n1010 VCC.n1009 0.00317857
R57732 VCC.n1015 VCC.n611 0.00317857
R57733 VCC.n1060 VCC.n584 0.00317857
R57734 VCC.n1069 VCC.n1068 0.00317857
R57735 VCC.n1086 VCC.n1085 0.00317857
R57736 VCC.n1092 VCC.n1091 0.00317857
R57737 VCC.n1092 VCC.n556 0.00317857
R57738 VCC.n1011 VCC.n616 0.00317857
R57739 VCC.n1017 VCC.n1016 0.00317857
R57740 VCC.n1059 VCC.n585 0.00317857
R57741 VCC.n1087 VCC.n567 0.00317857
R57742 VCC.n1093 VCC.n1090 0.00317857
R57743 VCC.n1569 VCC.n1568 0.00317857
R57744 VCC.n1575 VCC.n1169 0.00317857
R57745 VCC.n1614 VCC.n1148 0.00317857
R57746 VCC.n1139 VCC.n1128 0.00317857
R57747 VCC.n1633 VCC.n1118 0.00317857
R57748 VCC.n1640 VCC.n1639 0.00317857
R57749 VCC.n1639 VCC.n1110 0.00317857
R57750 VCC.n1570 VCC.n1173 0.00317857
R57751 VCC.n1574 VCC.n1573 0.00317857
R57752 VCC.n1613 VCC.n1149 0.00317857
R57753 VCC.n1634 VCC.n1120 0.00317857
R57754 VCC.n1638 VCC.n1637 0.00317857
R57755 VCC.n1441 VCC.n1234 0.00317857
R57756 VCC.n1452 VCC.n1225 0.00317857
R57757 VCC.n1452 VCC.n1451 0.00317857
R57758 VCC.n1214 VCC.n1207 0.00317857
R57759 VCC.n1492 VCC.n1208 0.00317857
R57760 VCC.n1498 VCC.n1497 0.00317857
R57761 VCC.n1550 VCC.n1182 0.00317857
R57762 VCC.n1550 VCC.n1549 0.00317857
R57763 VCC.n1555 VCC.n1177 0.00317857
R57764 VCC.n1440 VCC.n1428 0.00317857
R57765 VCC.n1453 VCC.n1224 0.00317857
R57766 VCC.n1491 VCC.n1490 0.00317857
R57767 VCC.n1551 VCC.n1181 0.00317857
R57768 VCC.n1554 VCC.n1178 0.00317857
R57769 VCC.n1330 VCC.n1295 0.00317857
R57770 VCC.n1372 VCC.n1267 0.00317857
R57771 VCC.n1415 VCC.n1414 0.00317857
R57772 VCC.n1420 VCC.n1239 0.00317857
R57773 VCC.n1326 VCC.n1300 0.00317857
R57774 VCC.n1329 VCC.n1296 0.00317857
R57775 VCC.n1371 VCC.n1273 0.00317857
R57776 VCC.n1416 VCC.n1243 0.00317857
R57777 VCC.n1419 VCC.n1240 0.00317857
R57778 VCC.n1881 VCC.n1846 0.00317857
R57779 VCC.n1923 VCC.n1818 0.00317857
R57780 VCC.n1966 VCC.n1965 0.00317857
R57781 VCC.n1971 VCC.n1790 0.00317857
R57782 VCC.n1877 VCC.n1851 0.00317857
R57783 VCC.n1880 VCC.n1847 0.00317857
R57784 VCC.n1922 VCC.n1824 0.00317857
R57785 VCC.n1967 VCC.n1794 0.00317857
R57786 VCC.n1970 VCC.n1791 0.00317857
R57787 VCC.n1993 VCC.n1786 0.00317857
R57788 VCC.n2004 VCC.n1777 0.00317857
R57789 VCC.n2004 VCC.n2003 0.00317857
R57790 VCC.n1766 VCC.n1759 0.00317857
R57791 VCC.n2044 VCC.n1760 0.00317857
R57792 VCC.n2050 VCC.n2049 0.00317857
R57793 VCC.n2101 VCC.n1734 0.00317857
R57794 VCC.n2101 VCC.n2100 0.00317857
R57795 VCC.n2106 VCC.n1729 0.00317857
R57796 VCC.n1980 VCC.n1979 0.00317857
R57797 VCC.n2005 VCC.n1776 0.00317857
R57798 VCC.n2043 VCC.n2042 0.00317857
R57799 VCC.n2102 VCC.n1733 0.00317857
R57800 VCC.n2105 VCC.n1730 0.00317857
R57801 VCC.n2119 VCC.n2118 0.00317857
R57802 VCC.n2124 VCC.n1720 0.00317857
R57803 VCC.n2169 VCC.n1693 0.00317857
R57804 VCC.n2178 VCC.n2177 0.00317857
R57805 VCC.n2195 VCC.n2194 0.00317857
R57806 VCC.n2201 VCC.n2200 0.00317857
R57807 VCC.n2201 VCC.n1665 0.00317857
R57808 VCC.n2120 VCC.n1725 0.00317857
R57809 VCC.n2126 VCC.n2125 0.00317857
R57810 VCC.n2168 VCC.n1694 0.00317857
R57811 VCC.n2196 VCC.n1676 0.00317857
R57812 VCC.n2202 VCC.n2199 0.00317857
R57813 VCC.n2678 VCC.n2677 0.00317857
R57814 VCC.n2684 VCC.n2278 0.00317857
R57815 VCC.n2723 VCC.n2257 0.00317857
R57816 VCC.n2248 VCC.n2237 0.00317857
R57817 VCC.n2742 VCC.n2227 0.00317857
R57818 VCC.n2749 VCC.n2748 0.00317857
R57819 VCC.n2748 VCC.n2219 0.00317857
R57820 VCC.n2679 VCC.n2282 0.00317857
R57821 VCC.n2683 VCC.n2682 0.00317857
R57822 VCC.n2722 VCC.n2258 0.00317857
R57823 VCC.n2743 VCC.n2229 0.00317857
R57824 VCC.n2747 VCC.n2746 0.00317857
R57825 VCC.n2550 VCC.n2343 0.00317857
R57826 VCC.n2561 VCC.n2334 0.00317857
R57827 VCC.n2561 VCC.n2560 0.00317857
R57828 VCC.n2323 VCC.n2316 0.00317857
R57829 VCC.n2601 VCC.n2317 0.00317857
R57830 VCC.n2607 VCC.n2606 0.00317857
R57831 VCC.n2659 VCC.n2291 0.00317857
R57832 VCC.n2659 VCC.n2658 0.00317857
R57833 VCC.n2664 VCC.n2286 0.00317857
R57834 VCC.n2549 VCC.n2537 0.00317857
R57835 VCC.n2562 VCC.n2333 0.00317857
R57836 VCC.n2600 VCC.n2599 0.00317857
R57837 VCC.n2660 VCC.n2290 0.00317857
R57838 VCC.n2663 VCC.n2287 0.00317857
R57839 VCC.n2439 VCC.n2404 0.00317857
R57840 VCC.n2481 VCC.n2376 0.00317857
R57841 VCC.n2524 VCC.n2523 0.00317857
R57842 VCC.n2529 VCC.n2348 0.00317857
R57843 VCC.n2435 VCC.n2409 0.00317857
R57844 VCC.n2438 VCC.n2405 0.00317857
R57845 VCC.n2480 VCC.n2382 0.00317857
R57846 VCC.n2525 VCC.n2352 0.00317857
R57847 VCC.n2528 VCC.n2349 0.00317857
R57848 VCC.n2990 VCC.n2955 0.00317857
R57849 VCC.n3032 VCC.n2927 0.00317857
R57850 VCC.n3075 VCC.n3074 0.00317857
R57851 VCC.n3080 VCC.n2899 0.00317857
R57852 VCC.n2986 VCC.n2960 0.00317857
R57853 VCC.n2989 VCC.n2956 0.00317857
R57854 VCC.n3031 VCC.n2933 0.00317857
R57855 VCC.n3076 VCC.n2903 0.00317857
R57856 VCC.n3079 VCC.n2900 0.00317857
R57857 VCC.n3102 VCC.n2895 0.00317857
R57858 VCC.n3113 VCC.n2886 0.00317857
R57859 VCC.n3113 VCC.n3112 0.00317857
R57860 VCC.n2875 VCC.n2868 0.00317857
R57861 VCC.n3153 VCC.n2869 0.00317857
R57862 VCC.n3159 VCC.n3158 0.00317857
R57863 VCC.n3210 VCC.n2843 0.00317857
R57864 VCC.n3210 VCC.n3209 0.00317857
R57865 VCC.n3215 VCC.n2838 0.00317857
R57866 VCC.n3089 VCC.n3088 0.00317857
R57867 VCC.n3114 VCC.n2885 0.00317857
R57868 VCC.n3152 VCC.n3151 0.00317857
R57869 VCC.n3211 VCC.n2842 0.00317857
R57870 VCC.n3214 VCC.n2839 0.00317857
R57871 VCC.n3228 VCC.n3227 0.00317857
R57872 VCC.n3233 VCC.n2829 0.00317857
R57873 VCC.n3278 VCC.n2802 0.00317857
R57874 VCC.n3287 VCC.n3286 0.00317857
R57875 VCC.n3304 VCC.n3303 0.00317857
R57876 VCC.n3310 VCC.n3309 0.00317857
R57877 VCC.n3310 VCC.n2774 0.00317857
R57878 VCC.n3229 VCC.n2834 0.00317857
R57879 VCC.n3235 VCC.n3234 0.00317857
R57880 VCC.n3277 VCC.n2803 0.00317857
R57881 VCC.n3305 VCC.n2785 0.00317857
R57882 VCC.n3311 VCC.n3308 0.00317857
R57883 VCC.n3787 VCC.n3786 0.00317857
R57884 VCC.n3793 VCC.n3387 0.00317857
R57885 VCC.n3832 VCC.n3366 0.00317857
R57886 VCC.n3357 VCC.n3346 0.00317857
R57887 VCC.n3851 VCC.n3336 0.00317857
R57888 VCC.n3858 VCC.n3857 0.00317857
R57889 VCC.n3857 VCC.n3328 0.00317857
R57890 VCC.n3788 VCC.n3391 0.00317857
R57891 VCC.n3792 VCC.n3791 0.00317857
R57892 VCC.n3831 VCC.n3367 0.00317857
R57893 VCC.n3852 VCC.n3338 0.00317857
R57894 VCC.n3856 VCC.n3855 0.00317857
R57895 VCC.n3659 VCC.n3452 0.00317857
R57896 VCC.n3670 VCC.n3443 0.00317857
R57897 VCC.n3670 VCC.n3669 0.00317857
R57898 VCC.n3432 VCC.n3425 0.00317857
R57899 VCC.n3710 VCC.n3426 0.00317857
R57900 VCC.n3716 VCC.n3715 0.00317857
R57901 VCC.n3768 VCC.n3400 0.00317857
R57902 VCC.n3768 VCC.n3767 0.00317857
R57903 VCC.n3773 VCC.n3395 0.00317857
R57904 VCC.n3658 VCC.n3646 0.00317857
R57905 VCC.n3671 VCC.n3442 0.00317857
R57906 VCC.n3709 VCC.n3708 0.00317857
R57907 VCC.n3769 VCC.n3399 0.00317857
R57908 VCC.n3772 VCC.n3396 0.00317857
R57909 VCC.n3548 VCC.n3513 0.00317857
R57910 VCC.n3590 VCC.n3485 0.00317857
R57911 VCC.n3633 VCC.n3632 0.00317857
R57912 VCC.n3638 VCC.n3457 0.00317857
R57913 VCC.n3544 VCC.n3518 0.00317857
R57914 VCC.n3547 VCC.n3514 0.00317857
R57915 VCC.n3589 VCC.n3491 0.00317857
R57916 VCC.n3634 VCC.n3461 0.00317857
R57917 VCC.n3637 VCC.n3458 0.00317857
R57918 VCC.n4099 VCC.n4064 0.00317857
R57919 VCC.n4141 VCC.n4036 0.00317857
R57920 VCC.n4184 VCC.n4183 0.00317857
R57921 VCC.n4189 VCC.n4008 0.00317857
R57922 VCC.n4095 VCC.n4069 0.00317857
R57923 VCC.n4098 VCC.n4065 0.00317857
R57924 VCC.n4140 VCC.n4042 0.00317857
R57925 VCC.n4185 VCC.n4012 0.00317857
R57926 VCC.n4188 VCC.n4009 0.00317857
R57927 VCC.n4211 VCC.n4004 0.00317857
R57928 VCC.n4222 VCC.n3995 0.00317857
R57929 VCC.n4222 VCC.n4221 0.00317857
R57930 VCC.n3984 VCC.n3977 0.00317857
R57931 VCC.n4262 VCC.n3978 0.00317857
R57932 VCC.n4268 VCC.n4267 0.00317857
R57933 VCC.n4319 VCC.n3952 0.00317857
R57934 VCC.n4319 VCC.n4318 0.00317857
R57935 VCC.n4324 VCC.n3947 0.00317857
R57936 VCC.n4198 VCC.n4197 0.00317857
R57937 VCC.n4223 VCC.n3994 0.00317857
R57938 VCC.n4261 VCC.n4260 0.00317857
R57939 VCC.n4320 VCC.n3951 0.00317857
R57940 VCC.n4323 VCC.n3948 0.00317857
R57941 VCC.n4337 VCC.n4336 0.00317857
R57942 VCC.n4342 VCC.n3938 0.00317857
R57943 VCC.n4387 VCC.n3911 0.00317857
R57944 VCC.n4396 VCC.n4395 0.00317857
R57945 VCC.n4413 VCC.n4412 0.00317857
R57946 VCC.n4419 VCC.n4418 0.00317857
R57947 VCC.n4419 VCC.n3883 0.00317857
R57948 VCC.n4338 VCC.n3943 0.00317857
R57949 VCC.n4344 VCC.n4343 0.00317857
R57950 VCC.n4386 VCC.n3912 0.00317857
R57951 VCC.n4414 VCC.n3894 0.00317857
R57952 VCC.n4420 VCC.n4417 0.00317857
R57953 VCC.n4896 VCC.n4895 0.00317857
R57954 VCC.n4902 VCC.n4496 0.00317857
R57955 VCC.n4941 VCC.n4475 0.00317857
R57956 VCC.n4466 VCC.n4455 0.00317857
R57957 VCC.n4960 VCC.n4445 0.00317857
R57958 VCC.n4967 VCC.n4966 0.00317857
R57959 VCC.n4966 VCC.n4437 0.00317857
R57960 VCC.n4897 VCC.n4500 0.00317857
R57961 VCC.n4901 VCC.n4900 0.00317857
R57962 VCC.n4940 VCC.n4476 0.00317857
R57963 VCC.n4961 VCC.n4447 0.00317857
R57964 VCC.n4965 VCC.n4964 0.00317857
R57965 VCC.n4768 VCC.n4561 0.00317857
R57966 VCC.n4779 VCC.n4552 0.00317857
R57967 VCC.n4779 VCC.n4778 0.00317857
R57968 VCC.n4541 VCC.n4534 0.00317857
R57969 VCC.n4819 VCC.n4535 0.00317857
R57970 VCC.n4825 VCC.n4824 0.00317857
R57971 VCC.n4877 VCC.n4509 0.00317857
R57972 VCC.n4877 VCC.n4876 0.00317857
R57973 VCC.n4882 VCC.n4504 0.00317857
R57974 VCC.n4767 VCC.n4755 0.00317857
R57975 VCC.n4780 VCC.n4551 0.00317857
R57976 VCC.n4818 VCC.n4817 0.00317857
R57977 VCC.n4878 VCC.n4508 0.00317857
R57978 VCC.n4881 VCC.n4505 0.00317857
R57979 VCC.n4657 VCC.n4622 0.00317857
R57980 VCC.n4699 VCC.n4594 0.00317857
R57981 VCC.n4742 VCC.n4741 0.00317857
R57982 VCC.n4747 VCC.n4566 0.00317857
R57983 VCC.n4653 VCC.n4627 0.00317857
R57984 VCC.n4656 VCC.n4623 0.00317857
R57985 VCC.n4698 VCC.n4600 0.00317857
R57986 VCC.n4743 VCC.n4570 0.00317857
R57987 VCC.n4746 VCC.n4567 0.00317857
R57988 VCC.n5208 VCC.n5173 0.00317857
R57989 VCC.n5250 VCC.n5145 0.00317857
R57990 VCC.n5293 VCC.n5292 0.00317857
R57991 VCC.n5298 VCC.n5117 0.00317857
R57992 VCC.n5204 VCC.n5178 0.00317857
R57993 VCC.n5207 VCC.n5174 0.00317857
R57994 VCC.n5249 VCC.n5151 0.00317857
R57995 VCC.n5294 VCC.n5121 0.00317857
R57996 VCC.n5297 VCC.n5118 0.00317857
R57997 VCC.n5320 VCC.n5113 0.00317857
R57998 VCC.n5331 VCC.n5104 0.00317857
R57999 VCC.n5331 VCC.n5330 0.00317857
R58000 VCC.n5093 VCC.n5086 0.00317857
R58001 VCC.n5371 VCC.n5087 0.00317857
R58002 VCC.n5377 VCC.n5376 0.00317857
R58003 VCC.n5428 VCC.n5061 0.00317857
R58004 VCC.n5428 VCC.n5427 0.00317857
R58005 VCC.n5433 VCC.n5056 0.00317857
R58006 VCC.n5307 VCC.n5306 0.00317857
R58007 VCC.n5332 VCC.n5103 0.00317857
R58008 VCC.n5370 VCC.n5369 0.00317857
R58009 VCC.n5429 VCC.n5060 0.00317857
R58010 VCC.n5432 VCC.n5057 0.00317857
R58011 VCC.n5446 VCC.n5445 0.00317857
R58012 VCC.n5451 VCC.n5047 0.00317857
R58013 VCC.n5496 VCC.n5020 0.00317857
R58014 VCC.n5505 VCC.n5504 0.00317857
R58015 VCC.n5522 VCC.n5521 0.00317857
R58016 VCC.n5528 VCC.n5527 0.00317857
R58017 VCC.n5528 VCC.n4992 0.00317857
R58018 VCC.n5447 VCC.n5052 0.00317857
R58019 VCC.n5453 VCC.n5452 0.00317857
R58020 VCC.n5495 VCC.n5021 0.00317857
R58021 VCC.n5523 VCC.n5003 0.00317857
R58022 VCC.n5529 VCC.n5526 0.00317857
R58023 VCC.n6005 VCC.n6004 0.00317857
R58024 VCC.n6011 VCC.n5605 0.00317857
R58025 VCC.n6050 VCC.n5584 0.00317857
R58026 VCC.n5575 VCC.n5564 0.00317857
R58027 VCC.n6069 VCC.n5554 0.00317857
R58028 VCC.n6076 VCC.n6075 0.00317857
R58029 VCC.n6075 VCC.n5546 0.00317857
R58030 VCC.n6006 VCC.n5609 0.00317857
R58031 VCC.n6010 VCC.n6009 0.00317857
R58032 VCC.n6049 VCC.n5585 0.00317857
R58033 VCC.n6070 VCC.n5556 0.00317857
R58034 VCC.n6074 VCC.n6073 0.00317857
R58035 VCC.n5877 VCC.n5670 0.00317857
R58036 VCC.n5888 VCC.n5661 0.00317857
R58037 VCC.n5888 VCC.n5887 0.00317857
R58038 VCC.n5650 VCC.n5643 0.00317857
R58039 VCC.n5928 VCC.n5644 0.00317857
R58040 VCC.n5934 VCC.n5933 0.00317857
R58041 VCC.n5986 VCC.n5618 0.00317857
R58042 VCC.n5986 VCC.n5985 0.00317857
R58043 VCC.n5991 VCC.n5613 0.00317857
R58044 VCC.n5876 VCC.n5864 0.00317857
R58045 VCC.n5889 VCC.n5660 0.00317857
R58046 VCC.n5927 VCC.n5926 0.00317857
R58047 VCC.n5987 VCC.n5617 0.00317857
R58048 VCC.n5990 VCC.n5614 0.00317857
R58049 VCC.n5766 VCC.n5731 0.00317857
R58050 VCC.n5808 VCC.n5703 0.00317857
R58051 VCC.n5851 VCC.n5850 0.00317857
R58052 VCC.n5856 VCC.n5675 0.00317857
R58053 VCC.n5762 VCC.n5736 0.00317857
R58054 VCC.n5765 VCC.n5732 0.00317857
R58055 VCC.n5807 VCC.n5709 0.00317857
R58056 VCC.n5852 VCC.n5679 0.00317857
R58057 VCC.n5855 VCC.n5676 0.00317857
R58058 VCC.n6317 VCC.n6282 0.00317857
R58059 VCC.n6359 VCC.n6254 0.00317857
R58060 VCC.n6402 VCC.n6401 0.00317857
R58061 VCC.n6407 VCC.n6226 0.00317857
R58062 VCC.n6313 VCC.n6287 0.00317857
R58063 VCC.n6316 VCC.n6283 0.00317857
R58064 VCC.n6358 VCC.n6260 0.00317857
R58065 VCC.n6403 VCC.n6230 0.00317857
R58066 VCC.n6406 VCC.n6227 0.00317857
R58067 VCC.n6429 VCC.n6222 0.00317857
R58068 VCC.n6440 VCC.n6213 0.00317857
R58069 VCC.n6440 VCC.n6439 0.00317857
R58070 VCC.n6202 VCC.n6195 0.00317857
R58071 VCC.n6480 VCC.n6196 0.00317857
R58072 VCC.n6486 VCC.n6485 0.00317857
R58073 VCC.n6537 VCC.n6170 0.00317857
R58074 VCC.n6537 VCC.n6536 0.00317857
R58075 VCC.n6542 VCC.n6165 0.00317857
R58076 VCC.n6416 VCC.n6415 0.00317857
R58077 VCC.n6441 VCC.n6212 0.00317857
R58078 VCC.n6479 VCC.n6478 0.00317857
R58079 VCC.n6538 VCC.n6169 0.00317857
R58080 VCC.n6541 VCC.n6166 0.00317857
R58081 VCC.n6555 VCC.n6554 0.00317857
R58082 VCC.n6560 VCC.n6156 0.00317857
R58083 VCC.n6605 VCC.n6129 0.00317857
R58084 VCC.n6614 VCC.n6613 0.00317857
R58085 VCC.n6631 VCC.n6630 0.00317857
R58086 VCC.n6637 VCC.n6636 0.00317857
R58087 VCC.n6637 VCC.n6101 0.00317857
R58088 VCC.n6556 VCC.n6161 0.00317857
R58089 VCC.n6562 VCC.n6561 0.00317857
R58090 VCC.n6604 VCC.n6130 0.00317857
R58091 VCC.n6632 VCC.n6112 0.00317857
R58092 VCC.n6638 VCC.n6635 0.00317857
R58093 VCC.n7114 VCC.n7113 0.00317857
R58094 VCC.n7120 VCC.n6714 0.00317857
R58095 VCC.n7159 VCC.n6693 0.00317857
R58096 VCC.n6684 VCC.n6673 0.00317857
R58097 VCC.n7178 VCC.n6663 0.00317857
R58098 VCC.n7185 VCC.n7184 0.00317857
R58099 VCC.n7184 VCC.n6655 0.00317857
R58100 VCC.n7115 VCC.n6718 0.00317857
R58101 VCC.n7119 VCC.n7118 0.00317857
R58102 VCC.n7158 VCC.n6694 0.00317857
R58103 VCC.n7179 VCC.n6665 0.00317857
R58104 VCC.n7183 VCC.n7182 0.00317857
R58105 VCC.n6986 VCC.n6779 0.00317857
R58106 VCC.n6997 VCC.n6770 0.00317857
R58107 VCC.n6997 VCC.n6996 0.00317857
R58108 VCC.n6759 VCC.n6752 0.00317857
R58109 VCC.n7037 VCC.n6753 0.00317857
R58110 VCC.n7043 VCC.n7042 0.00317857
R58111 VCC.n7095 VCC.n6727 0.00317857
R58112 VCC.n7095 VCC.n7094 0.00317857
R58113 VCC.n7100 VCC.n6722 0.00317857
R58114 VCC.n6985 VCC.n6973 0.00317857
R58115 VCC.n6998 VCC.n6769 0.00317857
R58116 VCC.n7036 VCC.n7035 0.00317857
R58117 VCC.n7096 VCC.n6726 0.00317857
R58118 VCC.n7099 VCC.n6723 0.00317857
R58119 VCC.n6875 VCC.n6840 0.00317857
R58120 VCC.n6917 VCC.n6812 0.00317857
R58121 VCC.n6960 VCC.n6959 0.00317857
R58122 VCC.n6965 VCC.n6784 0.00317857
R58123 VCC.n6871 VCC.n6845 0.00317857
R58124 VCC.n6874 VCC.n6841 0.00317857
R58125 VCC.n6916 VCC.n6818 0.00317857
R58126 VCC.n6961 VCC.n6788 0.00317857
R58127 VCC.n6964 VCC.n6785 0.00317857
R58128 VCC.n7426 VCC.n7391 0.00317857
R58129 VCC.n7468 VCC.n7363 0.00317857
R58130 VCC.n7511 VCC.n7510 0.00317857
R58131 VCC.n7516 VCC.n7335 0.00317857
R58132 VCC.n7422 VCC.n7396 0.00317857
R58133 VCC.n7425 VCC.n7392 0.00317857
R58134 VCC.n7467 VCC.n7369 0.00317857
R58135 VCC.n7512 VCC.n7339 0.00317857
R58136 VCC.n7515 VCC.n7336 0.00317857
R58137 VCC.n7538 VCC.n7331 0.00317857
R58138 VCC.n7549 VCC.n7322 0.00317857
R58139 VCC.n7549 VCC.n7548 0.00317857
R58140 VCC.n7311 VCC.n7304 0.00317857
R58141 VCC.n7589 VCC.n7305 0.00317857
R58142 VCC.n7595 VCC.n7594 0.00317857
R58143 VCC.n7646 VCC.n7279 0.00317857
R58144 VCC.n7646 VCC.n7645 0.00317857
R58145 VCC.n7651 VCC.n7274 0.00317857
R58146 VCC.n7525 VCC.n7524 0.00317857
R58147 VCC.n7550 VCC.n7321 0.00317857
R58148 VCC.n7588 VCC.n7587 0.00317857
R58149 VCC.n7647 VCC.n7278 0.00317857
R58150 VCC.n7650 VCC.n7275 0.00317857
R58151 VCC.n7664 VCC.n7663 0.00317857
R58152 VCC.n7669 VCC.n7265 0.00317857
R58153 VCC.n7714 VCC.n7238 0.00317857
R58154 VCC.n7723 VCC.n7722 0.00317857
R58155 VCC.n7740 VCC.n7739 0.00317857
R58156 VCC.n7746 VCC.n7745 0.00317857
R58157 VCC.n7746 VCC.n7210 0.00317857
R58158 VCC.n7665 VCC.n7270 0.00317857
R58159 VCC.n7671 VCC.n7670 0.00317857
R58160 VCC.n7713 VCC.n7239 0.00317857
R58161 VCC.n7741 VCC.n7221 0.00317857
R58162 VCC.n7747 VCC.n7744 0.00317857
R58163 VCC.n8223 VCC.n8222 0.00317857
R58164 VCC.n8229 VCC.n7823 0.00317857
R58165 VCC.n8268 VCC.n7802 0.00317857
R58166 VCC.n7793 VCC.n7782 0.00317857
R58167 VCC.n8287 VCC.n7772 0.00317857
R58168 VCC.n8294 VCC.n8293 0.00317857
R58169 VCC.n8293 VCC.n7764 0.00317857
R58170 VCC.n8224 VCC.n7827 0.00317857
R58171 VCC.n8228 VCC.n8227 0.00317857
R58172 VCC.n8267 VCC.n7803 0.00317857
R58173 VCC.n8288 VCC.n7774 0.00317857
R58174 VCC.n8292 VCC.n8291 0.00317857
R58175 VCC.n8095 VCC.n7888 0.00317857
R58176 VCC.n8106 VCC.n7879 0.00317857
R58177 VCC.n8106 VCC.n8105 0.00317857
R58178 VCC.n7868 VCC.n7861 0.00317857
R58179 VCC.n8146 VCC.n7862 0.00317857
R58180 VCC.n8152 VCC.n8151 0.00317857
R58181 VCC.n8204 VCC.n7836 0.00317857
R58182 VCC.n8204 VCC.n8203 0.00317857
R58183 VCC.n8209 VCC.n7831 0.00317857
R58184 VCC.n8094 VCC.n8082 0.00317857
R58185 VCC.n8107 VCC.n7878 0.00317857
R58186 VCC.n8145 VCC.n8144 0.00317857
R58187 VCC.n8205 VCC.n7835 0.00317857
R58188 VCC.n8208 VCC.n7832 0.00317857
R58189 VCC.n7984 VCC.n7949 0.00317857
R58190 VCC.n8026 VCC.n7921 0.00317857
R58191 VCC.n8069 VCC.n8068 0.00317857
R58192 VCC.n8074 VCC.n7893 0.00317857
R58193 VCC.n7980 VCC.n7954 0.00317857
R58194 VCC.n7983 VCC.n7950 0.00317857
R58195 VCC.n8025 VCC.n7927 0.00317857
R58196 VCC.n8070 VCC.n7897 0.00317857
R58197 VCC.n8073 VCC.n7894 0.00317857
R58198 VCC.n8647 VCC.n8440 0.00317857
R58199 VCC.n8658 VCC.n8431 0.00317857
R58200 VCC.n8658 VCC.n8657 0.00317857
R58201 VCC.n8420 VCC.n8413 0.00317857
R58202 VCC.n8698 VCC.n8414 0.00317857
R58203 VCC.n8704 VCC.n8703 0.00317857
R58204 VCC.n8755 VCC.n8388 0.00317857
R58205 VCC.n8755 VCC.n8754 0.00317857
R58206 VCC.n8760 VCC.n8383 0.00317857
R58207 VCC.n8634 VCC.n8633 0.00317857
R58208 VCC.n8659 VCC.n8430 0.00317857
R58209 VCC.n8697 VCC.n8696 0.00317857
R58210 VCC.n8756 VCC.n8387 0.00317857
R58211 VCC.n8759 VCC.n8384 0.00317857
R58212 VCC.n8773 VCC.n8772 0.00317857
R58213 VCC.n8778 VCC.n8374 0.00317857
R58214 VCC.n8823 VCC.n8347 0.00317857
R58215 VCC.n8832 VCC.n8831 0.00317857
R58216 VCC.n8849 VCC.n8848 0.00317857
R58217 VCC.n8855 VCC.n8854 0.00317857
R58218 VCC.n8855 VCC.n8319 0.00317857
R58219 VCC.n8774 VCC.n8379 0.00317857
R58220 VCC.n8780 VCC.n8779 0.00317857
R58221 VCC.n8822 VCC.n8348 0.00317857
R58222 VCC.n8850 VCC.n8330 0.00317857
R58223 VCC.n8856 VCC.n8853 0.00317857
R58224 VCC.n8535 VCC.n8500 0.00317857
R58225 VCC.n8577 VCC.n8472 0.00317857
R58226 VCC.n8620 VCC.n8619 0.00317857
R58227 VCC.n8625 VCC.n8444 0.00317857
R58228 VCC.n8531 VCC.n8505 0.00317857
R58229 VCC.n8534 VCC.n8501 0.00317857
R58230 VCC.n8576 VCC.n8478 0.00317857
R58231 VCC.n8621 VCC.n8448 0.00317857
R58232 VCC.n8624 VCC.n8445 0.00317857
R58233 VCC.n9332 VCC.n9331 0.00317857
R58234 VCC.n9338 VCC.n8932 0.00317857
R58235 VCC.n9377 VCC.n8911 0.00317857
R58236 VCC.n8902 VCC.n8891 0.00317857
R58237 VCC.n9396 VCC.n8881 0.00317857
R58238 VCC.n9403 VCC.n9402 0.00317857
R58239 VCC.n9402 VCC.n8873 0.00317857
R58240 VCC.n9333 VCC.n8936 0.00317857
R58241 VCC.n9337 VCC.n9336 0.00317857
R58242 VCC.n9376 VCC.n8912 0.00317857
R58243 VCC.n9397 VCC.n8883 0.00317857
R58244 VCC.n9401 VCC.n9400 0.00317857
R58245 VCC.n9204 VCC.n8997 0.00317857
R58246 VCC.n9215 VCC.n8988 0.00317857
R58247 VCC.n9215 VCC.n9214 0.00317857
R58248 VCC.n8977 VCC.n8970 0.00317857
R58249 VCC.n9255 VCC.n8971 0.00317857
R58250 VCC.n9261 VCC.n9260 0.00317857
R58251 VCC.n9313 VCC.n8945 0.00317857
R58252 VCC.n9313 VCC.n9312 0.00317857
R58253 VCC.n9318 VCC.n8940 0.00317857
R58254 VCC.n9203 VCC.n9191 0.00317857
R58255 VCC.n9216 VCC.n8987 0.00317857
R58256 VCC.n9254 VCC.n9253 0.00317857
R58257 VCC.n9314 VCC.n8944 0.00317857
R58258 VCC.n9317 VCC.n8941 0.00317857
R58259 VCC.n9093 VCC.n9058 0.00317857
R58260 VCC.n9135 VCC.n9030 0.00317857
R58261 VCC.n9178 VCC.n9177 0.00317857
R58262 VCC.n9183 VCC.n9002 0.00317857
R58263 VCC.n9089 VCC.n9063 0.00317857
R58264 VCC.n9092 VCC.n9059 0.00317857
R58265 VCC.n9134 VCC.n9036 0.00317857
R58266 VCC.n9179 VCC.n9006 0.00317857
R58267 VCC.n9182 VCC.n9003 0.00317857
R58268 VCC.n9644 VCC.n9609 0.00317857
R58269 VCC.n9686 VCC.n9581 0.00317857
R58270 VCC.n9729 VCC.n9728 0.00317857
R58271 VCC.n9734 VCC.n9553 0.00317857
R58272 VCC.n9640 VCC.n9614 0.00317857
R58273 VCC.n9643 VCC.n9610 0.00317857
R58274 VCC.n9685 VCC.n9587 0.00317857
R58275 VCC.n9730 VCC.n9557 0.00317857
R58276 VCC.n9733 VCC.n9554 0.00317857
R58277 VCC.n9756 VCC.n9549 0.00317857
R58278 VCC.n9767 VCC.n9540 0.00317857
R58279 VCC.n9767 VCC.n9766 0.00317857
R58280 VCC.n9529 VCC.n9522 0.00317857
R58281 VCC.n9807 VCC.n9523 0.00317857
R58282 VCC.n9813 VCC.n9812 0.00317857
R58283 VCC.n9864 VCC.n9497 0.00317857
R58284 VCC.n9864 VCC.n9863 0.00317857
R58285 VCC.n9869 VCC.n9492 0.00317857
R58286 VCC.n9743 VCC.n9742 0.00317857
R58287 VCC.n9768 VCC.n9539 0.00317857
R58288 VCC.n9806 VCC.n9805 0.00317857
R58289 VCC.n9865 VCC.n9496 0.00317857
R58290 VCC.n9868 VCC.n9493 0.00317857
R58291 VCC.n9882 VCC.n9881 0.00317857
R58292 VCC.n9887 VCC.n9483 0.00317857
R58293 VCC.n9932 VCC.n9456 0.00317857
R58294 VCC.n9941 VCC.n9940 0.00317857
R58295 VCC.n9958 VCC.n9957 0.00317857
R58296 VCC.n9964 VCC.n9963 0.00317857
R58297 VCC.n9964 VCC.n9428 0.00317857
R58298 VCC.n9883 VCC.n9488 0.00317857
R58299 VCC.n9889 VCC.n9888 0.00317857
R58300 VCC.n9931 VCC.n9457 0.00317857
R58301 VCC.n9959 VCC.n9439 0.00317857
R58302 VCC.n9965 VCC.n9962 0.00317857
R58303 VCC.n10440 VCC.n10439 0.00317857
R58304 VCC.n10446 VCC.n10040 0.00317857
R58305 VCC.n10485 VCC.n10019 0.00317857
R58306 VCC.n10010 VCC.n9999 0.00317857
R58307 VCC.n10504 VCC.n9989 0.00317857
R58308 VCC.n10511 VCC.n10510 0.00317857
R58309 VCC.n10510 VCC.n9981 0.00317857
R58310 VCC.n10441 VCC.n10044 0.00317857
R58311 VCC.n10445 VCC.n10444 0.00317857
R58312 VCC.n10484 VCC.n10020 0.00317857
R58313 VCC.n10505 VCC.n9991 0.00317857
R58314 VCC.n10509 VCC.n10508 0.00317857
R58315 VCC.n10312 VCC.n10105 0.00317857
R58316 VCC.n10323 VCC.n10096 0.00317857
R58317 VCC.n10323 VCC.n10322 0.00317857
R58318 VCC.n10085 VCC.n10078 0.00317857
R58319 VCC.n10363 VCC.n10079 0.00317857
R58320 VCC.n10369 VCC.n10368 0.00317857
R58321 VCC.n10421 VCC.n10053 0.00317857
R58322 VCC.n10421 VCC.n10420 0.00317857
R58323 VCC.n10426 VCC.n10048 0.00317857
R58324 VCC.n10311 VCC.n10299 0.00317857
R58325 VCC.n10324 VCC.n10095 0.00317857
R58326 VCC.n10362 VCC.n10361 0.00317857
R58327 VCC.n10422 VCC.n10052 0.00317857
R58328 VCC.n10425 VCC.n10049 0.00317857
R58329 VCC.n10201 VCC.n10166 0.00317857
R58330 VCC.n10243 VCC.n10138 0.00317857
R58331 VCC.n10286 VCC.n10285 0.00317857
R58332 VCC.n10291 VCC.n10110 0.00317857
R58333 VCC.n10197 VCC.n10171 0.00317857
R58334 VCC.n10200 VCC.n10167 0.00317857
R58335 VCC.n10242 VCC.n10144 0.00317857
R58336 VCC.n10287 VCC.n10114 0.00317857
R58337 VCC.n10290 VCC.n10111 0.00317857
R58338 VCC.n10751 VCC.n10716 0.00317857
R58339 VCC.n10793 VCC.n10688 0.00317857
R58340 VCC.n10836 VCC.n10835 0.00317857
R58341 VCC.n10841 VCC.n10660 0.00317857
R58342 VCC.n10747 VCC.n10721 0.00317857
R58343 VCC.n10750 VCC.n10717 0.00317857
R58344 VCC.n10792 VCC.n10694 0.00317857
R58345 VCC.n10837 VCC.n10664 0.00317857
R58346 VCC.n10840 VCC.n10661 0.00317857
R58347 VCC.n10863 VCC.n10656 0.00317857
R58348 VCC.n10874 VCC.n10647 0.00317857
R58349 VCC.n10874 VCC.n10873 0.00317857
R58350 VCC.n10636 VCC.n10629 0.00317857
R58351 VCC.n10914 VCC.n10630 0.00317857
R58352 VCC.n10920 VCC.n10919 0.00317857
R58353 VCC.n10971 VCC.n10604 0.00317857
R58354 VCC.n10971 VCC.n10970 0.00317857
R58355 VCC.n10976 VCC.n10599 0.00317857
R58356 VCC.n10850 VCC.n10849 0.00317857
R58357 VCC.n10875 VCC.n10646 0.00317857
R58358 VCC.n10913 VCC.n10912 0.00317857
R58359 VCC.n10972 VCC.n10603 0.00317857
R58360 VCC.n10975 VCC.n10600 0.00317857
R58361 VCC.n10989 VCC.n10988 0.00317857
R58362 VCC.n10994 VCC.n10590 0.00317857
R58363 VCC.n11039 VCC.n10563 0.00317857
R58364 VCC.n11048 VCC.n11047 0.00317857
R58365 VCC.n11065 VCC.n11064 0.00317857
R58366 VCC.n11071 VCC.n11070 0.00317857
R58367 VCC.n11071 VCC.n10535 0.00317857
R58368 VCC.n10990 VCC.n10595 0.00317857
R58369 VCC.n10996 VCC.n10995 0.00317857
R58370 VCC.n11038 VCC.n10564 0.00317857
R58371 VCC.n11066 VCC.n10546 0.00317857
R58372 VCC.n11072 VCC.n11069 0.00317857
R58373 VCC.n11547 VCC.n11546 0.00317857
R58374 VCC.n11553 VCC.n11147 0.00317857
R58375 VCC.n11592 VCC.n11126 0.00317857
R58376 VCC.n11117 VCC.n11106 0.00317857
R58377 VCC.n11611 VCC.n11096 0.00317857
R58378 VCC.n11618 VCC.n11617 0.00317857
R58379 VCC.n11617 VCC.n11088 0.00317857
R58380 VCC.n11548 VCC.n11151 0.00317857
R58381 VCC.n11552 VCC.n11551 0.00317857
R58382 VCC.n11591 VCC.n11127 0.00317857
R58383 VCC.n11612 VCC.n11098 0.00317857
R58384 VCC.n11616 VCC.n11615 0.00317857
R58385 VCC.n11419 VCC.n11212 0.00317857
R58386 VCC.n11430 VCC.n11203 0.00317857
R58387 VCC.n11430 VCC.n11429 0.00317857
R58388 VCC.n11192 VCC.n11185 0.00317857
R58389 VCC.n11470 VCC.n11186 0.00317857
R58390 VCC.n11476 VCC.n11475 0.00317857
R58391 VCC.n11528 VCC.n11160 0.00317857
R58392 VCC.n11528 VCC.n11527 0.00317857
R58393 VCC.n11533 VCC.n11155 0.00317857
R58394 VCC.n11418 VCC.n11406 0.00317857
R58395 VCC.n11431 VCC.n11202 0.00317857
R58396 VCC.n11469 VCC.n11468 0.00317857
R58397 VCC.n11529 VCC.n11159 0.00317857
R58398 VCC.n11532 VCC.n11156 0.00317857
R58399 VCC.n11308 VCC.n11273 0.00317857
R58400 VCC.n11350 VCC.n11245 0.00317857
R58401 VCC.n11393 VCC.n11392 0.00317857
R58402 VCC.n11398 VCC.n11217 0.00317857
R58403 VCC.n11304 VCC.n11278 0.00317857
R58404 VCC.n11307 VCC.n11274 0.00317857
R58405 VCC.n11349 VCC.n11251 0.00317857
R58406 VCC.n11394 VCC.n11221 0.00317857
R58407 VCC.n11397 VCC.n11218 0.00317857
R58408 VCC.n11858 VCC.n11823 0.00317857
R58409 VCC.n11900 VCC.n11795 0.00317857
R58410 VCC.n11943 VCC.n11942 0.00317857
R58411 VCC.n11948 VCC.n11767 0.00317857
R58412 VCC.n11854 VCC.n11828 0.00317857
R58413 VCC.n11857 VCC.n11824 0.00317857
R58414 VCC.n11899 VCC.n11801 0.00317857
R58415 VCC.n11944 VCC.n11771 0.00317857
R58416 VCC.n11947 VCC.n11768 0.00317857
R58417 VCC.n11970 VCC.n11763 0.00317857
R58418 VCC.n11981 VCC.n11754 0.00317857
R58419 VCC.n11981 VCC.n11980 0.00317857
R58420 VCC.n11743 VCC.n11736 0.00317857
R58421 VCC.n12021 VCC.n11737 0.00317857
R58422 VCC.n12027 VCC.n12026 0.00317857
R58423 VCC.n12078 VCC.n11711 0.00317857
R58424 VCC.n12078 VCC.n12077 0.00317857
R58425 VCC.n12083 VCC.n11706 0.00317857
R58426 VCC.n11957 VCC.n11956 0.00317857
R58427 VCC.n11982 VCC.n11753 0.00317857
R58428 VCC.n12020 VCC.n12019 0.00317857
R58429 VCC.n12079 VCC.n11710 0.00317857
R58430 VCC.n12082 VCC.n11707 0.00317857
R58431 VCC.n12096 VCC.n12095 0.00317857
R58432 VCC.n12101 VCC.n11697 0.00317857
R58433 VCC.n12146 VCC.n11670 0.00317857
R58434 VCC.n12155 VCC.n12154 0.00317857
R58435 VCC.n12172 VCC.n12171 0.00317857
R58436 VCC.n12178 VCC.n12177 0.00317857
R58437 VCC.n12178 VCC.n11642 0.00317857
R58438 VCC.n12097 VCC.n11702 0.00317857
R58439 VCC.n12103 VCC.n12102 0.00317857
R58440 VCC.n12145 VCC.n11671 0.00317857
R58441 VCC.n12173 VCC.n11653 0.00317857
R58442 VCC.n12179 VCC.n12176 0.00317857
R58443 VCC.n12654 VCC.n12653 0.00317857
R58444 VCC.n12660 VCC.n12254 0.00317857
R58445 VCC.n12699 VCC.n12233 0.00317857
R58446 VCC.n12224 VCC.n12213 0.00317857
R58447 VCC.n12718 VCC.n12203 0.00317857
R58448 VCC.n12725 VCC.n12724 0.00317857
R58449 VCC.n12724 VCC.n12195 0.00317857
R58450 VCC.n12655 VCC.n12258 0.00317857
R58451 VCC.n12659 VCC.n12658 0.00317857
R58452 VCC.n12698 VCC.n12234 0.00317857
R58453 VCC.n12719 VCC.n12205 0.00317857
R58454 VCC.n12723 VCC.n12722 0.00317857
R58455 VCC.n12526 VCC.n12319 0.00317857
R58456 VCC.n12537 VCC.n12310 0.00317857
R58457 VCC.n12537 VCC.n12536 0.00317857
R58458 VCC.n12299 VCC.n12292 0.00317857
R58459 VCC.n12577 VCC.n12293 0.00317857
R58460 VCC.n12583 VCC.n12582 0.00317857
R58461 VCC.n12635 VCC.n12267 0.00317857
R58462 VCC.n12635 VCC.n12634 0.00317857
R58463 VCC.n12640 VCC.n12262 0.00317857
R58464 VCC.n12525 VCC.n12513 0.00317857
R58465 VCC.n12538 VCC.n12309 0.00317857
R58466 VCC.n12576 VCC.n12575 0.00317857
R58467 VCC.n12636 VCC.n12266 0.00317857
R58468 VCC.n12639 VCC.n12263 0.00317857
R58469 VCC.n12415 VCC.n12380 0.00317857
R58470 VCC.n12457 VCC.n12352 0.00317857
R58471 VCC.n12500 VCC.n12499 0.00317857
R58472 VCC.n12505 VCC.n12324 0.00317857
R58473 VCC.n12411 VCC.n12385 0.00317857
R58474 VCC.n12414 VCC.n12381 0.00317857
R58475 VCC.n12456 VCC.n12358 0.00317857
R58476 VCC.n12501 VCC.n12328 0.00317857
R58477 VCC.n12504 VCC.n12325 0.00317857
R58478 VCC.n12965 VCC.n12930 0.00317857
R58479 VCC.n13007 VCC.n12902 0.00317857
R58480 VCC.n13050 VCC.n13049 0.00317857
R58481 VCC.n13055 VCC.n12874 0.00317857
R58482 VCC.n12961 VCC.n12935 0.00317857
R58483 VCC.n12964 VCC.n12931 0.00317857
R58484 VCC.n13006 VCC.n12908 0.00317857
R58485 VCC.n13051 VCC.n12878 0.00317857
R58486 VCC.n13054 VCC.n12875 0.00317857
R58487 VCC.n13077 VCC.n12870 0.00317857
R58488 VCC.n13088 VCC.n12861 0.00317857
R58489 VCC.n13088 VCC.n13087 0.00317857
R58490 VCC.n12850 VCC.n12843 0.00317857
R58491 VCC.n13128 VCC.n12844 0.00317857
R58492 VCC.n13134 VCC.n13133 0.00317857
R58493 VCC.n13185 VCC.n12818 0.00317857
R58494 VCC.n13185 VCC.n13184 0.00317857
R58495 VCC.n13190 VCC.n12813 0.00317857
R58496 VCC.n13064 VCC.n13063 0.00317857
R58497 VCC.n13089 VCC.n12860 0.00317857
R58498 VCC.n13127 VCC.n13126 0.00317857
R58499 VCC.n13186 VCC.n12817 0.00317857
R58500 VCC.n13189 VCC.n12814 0.00317857
R58501 VCC.n13203 VCC.n13202 0.00317857
R58502 VCC.n13208 VCC.n12804 0.00317857
R58503 VCC.n13253 VCC.n12777 0.00317857
R58504 VCC.n13262 VCC.n13261 0.00317857
R58505 VCC.n13279 VCC.n13278 0.00317857
R58506 VCC.n13285 VCC.n13284 0.00317857
R58507 VCC.n13285 VCC.n12749 0.00317857
R58508 VCC.n13204 VCC.n12809 0.00317857
R58509 VCC.n13210 VCC.n13209 0.00317857
R58510 VCC.n13252 VCC.n12778 0.00317857
R58511 VCC.n13280 VCC.n12760 0.00317857
R58512 VCC.n13286 VCC.n13283 0.00317857
R58513 VCC.n13761 VCC.n13760 0.00317857
R58514 VCC.n13767 VCC.n13361 0.00317857
R58515 VCC.n13806 VCC.n13340 0.00317857
R58516 VCC.n13331 VCC.n13320 0.00317857
R58517 VCC.n13825 VCC.n13310 0.00317857
R58518 VCC.n13832 VCC.n13831 0.00317857
R58519 VCC.n13831 VCC.n13302 0.00317857
R58520 VCC.n13762 VCC.n13365 0.00317857
R58521 VCC.n13766 VCC.n13765 0.00317857
R58522 VCC.n13805 VCC.n13341 0.00317857
R58523 VCC.n13826 VCC.n13312 0.00317857
R58524 VCC.n13830 VCC.n13829 0.00317857
R58525 VCC.n13633 VCC.n13426 0.00317857
R58526 VCC.n13644 VCC.n13417 0.00317857
R58527 VCC.n13644 VCC.n13643 0.00317857
R58528 VCC.n13406 VCC.n13399 0.00317857
R58529 VCC.n13684 VCC.n13400 0.00317857
R58530 VCC.n13690 VCC.n13689 0.00317857
R58531 VCC.n13742 VCC.n13374 0.00317857
R58532 VCC.n13742 VCC.n13741 0.00317857
R58533 VCC.n13747 VCC.n13369 0.00317857
R58534 VCC.n13632 VCC.n13620 0.00317857
R58535 VCC.n13645 VCC.n13416 0.00317857
R58536 VCC.n13683 VCC.n13682 0.00317857
R58537 VCC.n13743 VCC.n13373 0.00317857
R58538 VCC.n13746 VCC.n13370 0.00317857
R58539 VCC.n13522 VCC.n13487 0.00317857
R58540 VCC.n13564 VCC.n13459 0.00317857
R58541 VCC.n13607 VCC.n13606 0.00317857
R58542 VCC.n13612 VCC.n13431 0.00317857
R58543 VCC.n13518 VCC.n13492 0.00317857
R58544 VCC.n13521 VCC.n13488 0.00317857
R58545 VCC.n13563 VCC.n13465 0.00317857
R58546 VCC.n13608 VCC.n13435 0.00317857
R58547 VCC.n13611 VCC.n13432 0.00317857
R58548 VCC.n14072 VCC.n14037 0.00317857
R58549 VCC.n14114 VCC.n14009 0.00317857
R58550 VCC.n14157 VCC.n14156 0.00317857
R58551 VCC.n14162 VCC.n13981 0.00317857
R58552 VCC.n14068 VCC.n14042 0.00317857
R58553 VCC.n14071 VCC.n14038 0.00317857
R58554 VCC.n14113 VCC.n14015 0.00317857
R58555 VCC.n14158 VCC.n13985 0.00317857
R58556 VCC.n14161 VCC.n13982 0.00317857
R58557 VCC.n14184 VCC.n13977 0.00317857
R58558 VCC.n14195 VCC.n13968 0.00317857
R58559 VCC.n14195 VCC.n14194 0.00317857
R58560 VCC.n13957 VCC.n13950 0.00317857
R58561 VCC.n14235 VCC.n13951 0.00317857
R58562 VCC.n14241 VCC.n14240 0.00317857
R58563 VCC.n14292 VCC.n13925 0.00317857
R58564 VCC.n14292 VCC.n14291 0.00317857
R58565 VCC.n14297 VCC.n13920 0.00317857
R58566 VCC.n14171 VCC.n14170 0.00317857
R58567 VCC.n14196 VCC.n13967 0.00317857
R58568 VCC.n14234 VCC.n14233 0.00317857
R58569 VCC.n14293 VCC.n13924 0.00317857
R58570 VCC.n14296 VCC.n13921 0.00317857
R58571 VCC.n14310 VCC.n14309 0.00317857
R58572 VCC.n14315 VCC.n13911 0.00317857
R58573 VCC.n14360 VCC.n13884 0.00317857
R58574 VCC.n14369 VCC.n14368 0.00317857
R58575 VCC.n14386 VCC.n14385 0.00317857
R58576 VCC.n14392 VCC.n14391 0.00317857
R58577 VCC.n14392 VCC.n13856 0.00317857
R58578 VCC.n14311 VCC.n13916 0.00317857
R58579 VCC.n14317 VCC.n14316 0.00317857
R58580 VCC.n14359 VCC.n13885 0.00317857
R58581 VCC.n14387 VCC.n13867 0.00317857
R58582 VCC.n14393 VCC.n14390 0.00317857
R58583 VCC.n14868 VCC.n14867 0.00317857
R58584 VCC.n14874 VCC.n14468 0.00317857
R58585 VCC.n14913 VCC.n14447 0.00317857
R58586 VCC.n14438 VCC.n14427 0.00317857
R58587 VCC.n14932 VCC.n14417 0.00317857
R58588 VCC.n14939 VCC.n14938 0.00317857
R58589 VCC.n14938 VCC.n14409 0.00317857
R58590 VCC.n14869 VCC.n14472 0.00317857
R58591 VCC.n14873 VCC.n14872 0.00317857
R58592 VCC.n14912 VCC.n14448 0.00317857
R58593 VCC.n14933 VCC.n14419 0.00317857
R58594 VCC.n14937 VCC.n14936 0.00317857
R58595 VCC.n14740 VCC.n14533 0.00317857
R58596 VCC.n14751 VCC.n14524 0.00317857
R58597 VCC.n14751 VCC.n14750 0.00317857
R58598 VCC.n14513 VCC.n14506 0.00317857
R58599 VCC.n14791 VCC.n14507 0.00317857
R58600 VCC.n14797 VCC.n14796 0.00317857
R58601 VCC.n14849 VCC.n14481 0.00317857
R58602 VCC.n14849 VCC.n14848 0.00317857
R58603 VCC.n14854 VCC.n14476 0.00317857
R58604 VCC.n14739 VCC.n14727 0.00317857
R58605 VCC.n14752 VCC.n14523 0.00317857
R58606 VCC.n14790 VCC.n14789 0.00317857
R58607 VCC.n14850 VCC.n14480 0.00317857
R58608 VCC.n14853 VCC.n14477 0.00317857
R58609 VCC.n14629 VCC.n14594 0.00317857
R58610 VCC.n14671 VCC.n14566 0.00317857
R58611 VCC.n14714 VCC.n14713 0.00317857
R58612 VCC.n14719 VCC.n14538 0.00317857
R58613 VCC.n14625 VCC.n14599 0.00317857
R58614 VCC.n14628 VCC.n14595 0.00317857
R58615 VCC.n14670 VCC.n14572 0.00317857
R58616 VCC.n14715 VCC.n14542 0.00317857
R58617 VCC.n14718 VCC.n14539 0.00317857
R58618 VCC.n15179 VCC.n15144 0.00317857
R58619 VCC.n15221 VCC.n15116 0.00317857
R58620 VCC.n15264 VCC.n15263 0.00317857
R58621 VCC.n15269 VCC.n15088 0.00317857
R58622 VCC.n15175 VCC.n15149 0.00317857
R58623 VCC.n15178 VCC.n15145 0.00317857
R58624 VCC.n15220 VCC.n15122 0.00317857
R58625 VCC.n15265 VCC.n15092 0.00317857
R58626 VCC.n15268 VCC.n15089 0.00317857
R58627 VCC.n15291 VCC.n15084 0.00317857
R58628 VCC.n15302 VCC.n15075 0.00317857
R58629 VCC.n15302 VCC.n15301 0.00317857
R58630 VCC.n15064 VCC.n15057 0.00317857
R58631 VCC.n15342 VCC.n15058 0.00317857
R58632 VCC.n15348 VCC.n15347 0.00317857
R58633 VCC.n15399 VCC.n15032 0.00317857
R58634 VCC.n15399 VCC.n15398 0.00317857
R58635 VCC.n15404 VCC.n15027 0.00317857
R58636 VCC.n15278 VCC.n15277 0.00317857
R58637 VCC.n15303 VCC.n15074 0.00317857
R58638 VCC.n15341 VCC.n15340 0.00317857
R58639 VCC.n15400 VCC.n15031 0.00317857
R58640 VCC.n15403 VCC.n15028 0.00317857
R58641 VCC.n15417 VCC.n15416 0.00317857
R58642 VCC.n15422 VCC.n15018 0.00317857
R58643 VCC.n15467 VCC.n14991 0.00317857
R58644 VCC.n15476 VCC.n15475 0.00317857
R58645 VCC.n15493 VCC.n15492 0.00317857
R58646 VCC.n15499 VCC.n15498 0.00317857
R58647 VCC.n15499 VCC.n14963 0.00317857
R58648 VCC.n15418 VCC.n15023 0.00317857
R58649 VCC.n15424 VCC.n15423 0.00317857
R58650 VCC.n15466 VCC.n14992 0.00317857
R58651 VCC.n15494 VCC.n14974 0.00317857
R58652 VCC.n15500 VCC.n15497 0.00317857
R58653 VCC.n15975 VCC.n15974 0.00317857
R58654 VCC.n15981 VCC.n15575 0.00317857
R58655 VCC.n16020 VCC.n15554 0.00317857
R58656 VCC.n15545 VCC.n15534 0.00317857
R58657 VCC.n16039 VCC.n15524 0.00317857
R58658 VCC.n16046 VCC.n16045 0.00317857
R58659 VCC.n16045 VCC.n15516 0.00317857
R58660 VCC.n15976 VCC.n15579 0.00317857
R58661 VCC.n15980 VCC.n15979 0.00317857
R58662 VCC.n16019 VCC.n15555 0.00317857
R58663 VCC.n16040 VCC.n15526 0.00317857
R58664 VCC.n16044 VCC.n16043 0.00317857
R58665 VCC.n15847 VCC.n15640 0.00317857
R58666 VCC.n15858 VCC.n15631 0.00317857
R58667 VCC.n15858 VCC.n15857 0.00317857
R58668 VCC.n15620 VCC.n15613 0.00317857
R58669 VCC.n15898 VCC.n15614 0.00317857
R58670 VCC.n15904 VCC.n15903 0.00317857
R58671 VCC.n15956 VCC.n15588 0.00317857
R58672 VCC.n15956 VCC.n15955 0.00317857
R58673 VCC.n15961 VCC.n15583 0.00317857
R58674 VCC.n15846 VCC.n15834 0.00317857
R58675 VCC.n15859 VCC.n15630 0.00317857
R58676 VCC.n15897 VCC.n15896 0.00317857
R58677 VCC.n15957 VCC.n15587 0.00317857
R58678 VCC.n15960 VCC.n15584 0.00317857
R58679 VCC.n15736 VCC.n15701 0.00317857
R58680 VCC.n15778 VCC.n15673 0.00317857
R58681 VCC.n15821 VCC.n15820 0.00317857
R58682 VCC.n15826 VCC.n15645 0.00317857
R58683 VCC.n15732 VCC.n15706 0.00317857
R58684 VCC.n15735 VCC.n15702 0.00317857
R58685 VCC.n15777 VCC.n15679 0.00317857
R58686 VCC.n15822 VCC.n15649 0.00317857
R58687 VCC.n15825 VCC.n15646 0.00317857
R58688 VCC.n16286 VCC.n16251 0.00317857
R58689 VCC.n16328 VCC.n16223 0.00317857
R58690 VCC.n16371 VCC.n16370 0.00317857
R58691 VCC.n16376 VCC.n16195 0.00317857
R58692 VCC.n16282 VCC.n16256 0.00317857
R58693 VCC.n16285 VCC.n16252 0.00317857
R58694 VCC.n16327 VCC.n16229 0.00317857
R58695 VCC.n16372 VCC.n16199 0.00317857
R58696 VCC.n16375 VCC.n16196 0.00317857
R58697 VCC.n16398 VCC.n16191 0.00317857
R58698 VCC.n16409 VCC.n16182 0.00317857
R58699 VCC.n16409 VCC.n16408 0.00317857
R58700 VCC.n16171 VCC.n16164 0.00317857
R58701 VCC.n16449 VCC.n16165 0.00317857
R58702 VCC.n16455 VCC.n16454 0.00317857
R58703 VCC.n16506 VCC.n16139 0.00317857
R58704 VCC.n16506 VCC.n16505 0.00317857
R58705 VCC.n16511 VCC.n16134 0.00317857
R58706 VCC.n16385 VCC.n16384 0.00317857
R58707 VCC.n16410 VCC.n16181 0.00317857
R58708 VCC.n16448 VCC.n16447 0.00317857
R58709 VCC.n16507 VCC.n16138 0.00317857
R58710 VCC.n16510 VCC.n16135 0.00317857
R58711 VCC.n16524 VCC.n16523 0.00317857
R58712 VCC.n16529 VCC.n16125 0.00317857
R58713 VCC.n16574 VCC.n16098 0.00317857
R58714 VCC.n16583 VCC.n16582 0.00317857
R58715 VCC.n16600 VCC.n16599 0.00317857
R58716 VCC.n16606 VCC.n16605 0.00317857
R58717 VCC.n16606 VCC.n16070 0.00317857
R58718 VCC.n16525 VCC.n16130 0.00317857
R58719 VCC.n16531 VCC.n16530 0.00317857
R58720 VCC.n16573 VCC.n16099 0.00317857
R58721 VCC.n16601 VCC.n16081 0.00317857
R58722 VCC.n16607 VCC.n16604 0.00317857
R58723 VCC.n17082 VCC.n17081 0.00317857
R58724 VCC.n17088 VCC.n16682 0.00317857
R58725 VCC.n17127 VCC.n16661 0.00317857
R58726 VCC.n16652 VCC.n16641 0.00317857
R58727 VCC.n17146 VCC.n16631 0.00317857
R58728 VCC.n17153 VCC.n17152 0.00317857
R58729 VCC.n17152 VCC.n16623 0.00317857
R58730 VCC.n17083 VCC.n16686 0.00317857
R58731 VCC.n17087 VCC.n17086 0.00317857
R58732 VCC.n17126 VCC.n16662 0.00317857
R58733 VCC.n17147 VCC.n16633 0.00317857
R58734 VCC.n17151 VCC.n17150 0.00317857
R58735 VCC.n16954 VCC.n16747 0.00317857
R58736 VCC.n16965 VCC.n16738 0.00317857
R58737 VCC.n16965 VCC.n16964 0.00317857
R58738 VCC.n16727 VCC.n16720 0.00317857
R58739 VCC.n17005 VCC.n16721 0.00317857
R58740 VCC.n17011 VCC.n17010 0.00317857
R58741 VCC.n17063 VCC.n16695 0.00317857
R58742 VCC.n17063 VCC.n17062 0.00317857
R58743 VCC.n17068 VCC.n16690 0.00317857
R58744 VCC.n16953 VCC.n16941 0.00317857
R58745 VCC.n16966 VCC.n16737 0.00317857
R58746 VCC.n17004 VCC.n17003 0.00317857
R58747 VCC.n17064 VCC.n16694 0.00317857
R58748 VCC.n17067 VCC.n16691 0.00317857
R58749 VCC.n16843 VCC.n16808 0.00317857
R58750 VCC.n16885 VCC.n16780 0.00317857
R58751 VCC.n16928 VCC.n16927 0.00317857
R58752 VCC.n16933 VCC.n16752 0.00317857
R58753 VCC.n16839 VCC.n16813 0.00317857
R58754 VCC.n16842 VCC.n16809 0.00317857
R58755 VCC.n16884 VCC.n16786 0.00317857
R58756 VCC.n16929 VCC.n16756 0.00317857
R58757 VCC.n16932 VCC.n16753 0.00317857
R58758 VCC.n17318 VCC.n17298 0.00317857
R58759 VCC.n17329 VCC.n17289 0.00317857
R58760 VCC.n17329 VCC.n17328 0.00317857
R58761 VCC.n17278 VCC.n17271 0.00317857
R58762 VCC.n17369 VCC.n17272 0.00317857
R58763 VCC.n17375 VCC.n17374 0.00317857
R58764 VCC.n17426 VCC.n17246 0.00317857
R58765 VCC.n17426 VCC.n17425 0.00317857
R58766 VCC.n17431 VCC.n17241 0.00317857
R58767 VCC.n17305 VCC.n17304 0.00317857
R58768 VCC.n17330 VCC.n17288 0.00317857
R58769 VCC.n17368 VCC.n17367 0.00317857
R58770 VCC.n17427 VCC.n17245 0.00317857
R58771 VCC.n17430 VCC.n17242 0.00317857
R58772 VCC.n17444 VCC.n17443 0.00317857
R58773 VCC.n17449 VCC.n17232 0.00317857
R58774 VCC.n17494 VCC.n17205 0.00317857
R58775 VCC.n17503 VCC.n17502 0.00317857
R58776 VCC.n17520 VCC.n17519 0.00317857
R58777 VCC.n17526 VCC.n17525 0.00317857
R58778 VCC.n17526 VCC.n17177 0.00317857
R58779 VCC.n17445 VCC.n17237 0.00317857
R58780 VCC.n17451 VCC.n17450 0.00317857
R58781 VCC.n17493 VCC.n17206 0.00317857
R58782 VCC.n17521 VCC.n17188 0.00317857
R58783 VCC.n17527 VCC.n17524 0.00317857
R58784 VCC.n8558 VCC.n8480 0.00316667
R58785 VCC.n8574 VCC.n8462 0.00316667
R58786 VCC.n215 VCC.n214 0.00228571
R58787 VCC.n222 VCC.n220 0.00228571
R58788 VCC.n162 VCC.n161 0.00228571
R58789 VCC.n278 VCC.n150 0.00228571
R58790 VCC.n352 VCC.n112 0.00228571
R58791 VCC.n478 VCC.n477 0.00228571
R58792 VCC.n489 VCC.n44 0.00228571
R58793 VCC.n501 VCC.n38 0.00228571
R58794 VCC.n522 VCC.n521 0.00228571
R58795 VCC.n502 VCC.n36 0.00228571
R58796 VCC.n767 VCC.n766 0.00228571
R58797 VCC.n774 VCC.n772 0.00228571
R58798 VCC.n714 VCC.n713 0.00228571
R58799 VCC.n830 VCC.n702 0.00228571
R58800 VCC.n904 VCC.n664 0.00228571
R58801 VCC.n1030 VCC.n1029 0.00228571
R58802 VCC.n1041 VCC.n596 0.00228571
R58803 VCC.n1053 VCC.n590 0.00228571
R58804 VCC.n1074 VCC.n1073 0.00228571
R58805 VCC.n1054 VCC.n588 0.00228571
R58806 VCC.n1596 VCC.n1595 0.00228571
R58807 VCC.n1592 VCC.n1588 0.00228571
R58808 VCC.n1605 VCC.n1146 0.00228571
R58809 VCC.n1624 VCC.n1134 0.00228571
R58810 VCC.n1607 VCC.n1606 0.00228571
R58811 VCC.n1461 VCC.n1221 0.00228571
R58812 VCC.n1325 VCC.n1324 0.00228571
R58813 VCC.n1332 VCC.n1330 0.00228571
R58814 VCC.n1272 VCC.n1271 0.00228571
R58815 VCC.n1388 VCC.n1260 0.00228571
R58816 VCC.n1876 VCC.n1875 0.00228571
R58817 VCC.n1883 VCC.n1881 0.00228571
R58818 VCC.n1823 VCC.n1822 0.00228571
R58819 VCC.n1939 VCC.n1811 0.00228571
R58820 VCC.n2013 VCC.n1773 0.00228571
R58821 VCC.n2139 VCC.n2138 0.00228571
R58822 VCC.n2150 VCC.n1705 0.00228571
R58823 VCC.n2162 VCC.n1699 0.00228571
R58824 VCC.n2183 VCC.n2182 0.00228571
R58825 VCC.n2163 VCC.n1697 0.00228571
R58826 VCC.n2705 VCC.n2704 0.00228571
R58827 VCC.n2701 VCC.n2697 0.00228571
R58828 VCC.n2714 VCC.n2255 0.00228571
R58829 VCC.n2733 VCC.n2243 0.00228571
R58830 VCC.n2716 VCC.n2715 0.00228571
R58831 VCC.n2570 VCC.n2330 0.00228571
R58832 VCC.n2434 VCC.n2433 0.00228571
R58833 VCC.n2441 VCC.n2439 0.00228571
R58834 VCC.n2381 VCC.n2380 0.00228571
R58835 VCC.n2497 VCC.n2369 0.00228571
R58836 VCC.n2985 VCC.n2984 0.00228571
R58837 VCC.n2992 VCC.n2990 0.00228571
R58838 VCC.n2932 VCC.n2931 0.00228571
R58839 VCC.n3048 VCC.n2920 0.00228571
R58840 VCC.n3122 VCC.n2882 0.00228571
R58841 VCC.n3248 VCC.n3247 0.00228571
R58842 VCC.n3259 VCC.n2814 0.00228571
R58843 VCC.n3271 VCC.n2808 0.00228571
R58844 VCC.n3292 VCC.n3291 0.00228571
R58845 VCC.n3272 VCC.n2806 0.00228571
R58846 VCC.n3814 VCC.n3813 0.00228571
R58847 VCC.n3810 VCC.n3806 0.00228571
R58848 VCC.n3823 VCC.n3364 0.00228571
R58849 VCC.n3842 VCC.n3352 0.00228571
R58850 VCC.n3825 VCC.n3824 0.00228571
R58851 VCC.n3679 VCC.n3439 0.00228571
R58852 VCC.n3543 VCC.n3542 0.00228571
R58853 VCC.n3550 VCC.n3548 0.00228571
R58854 VCC.n3490 VCC.n3489 0.00228571
R58855 VCC.n3606 VCC.n3478 0.00228571
R58856 VCC.n4094 VCC.n4093 0.00228571
R58857 VCC.n4101 VCC.n4099 0.00228571
R58858 VCC.n4041 VCC.n4040 0.00228571
R58859 VCC.n4157 VCC.n4029 0.00228571
R58860 VCC.n4231 VCC.n3991 0.00228571
R58861 VCC.n4357 VCC.n4356 0.00228571
R58862 VCC.n4368 VCC.n3923 0.00228571
R58863 VCC.n4380 VCC.n3917 0.00228571
R58864 VCC.n4401 VCC.n4400 0.00228571
R58865 VCC.n4381 VCC.n3915 0.00228571
R58866 VCC.n4923 VCC.n4922 0.00228571
R58867 VCC.n4919 VCC.n4915 0.00228571
R58868 VCC.n4932 VCC.n4473 0.00228571
R58869 VCC.n4951 VCC.n4461 0.00228571
R58870 VCC.n4934 VCC.n4933 0.00228571
R58871 VCC.n4788 VCC.n4548 0.00228571
R58872 VCC.n4652 VCC.n4651 0.00228571
R58873 VCC.n4659 VCC.n4657 0.00228571
R58874 VCC.n4599 VCC.n4598 0.00228571
R58875 VCC.n4715 VCC.n4587 0.00228571
R58876 VCC.n5203 VCC.n5202 0.00228571
R58877 VCC.n5210 VCC.n5208 0.00228571
R58878 VCC.n5150 VCC.n5149 0.00228571
R58879 VCC.n5266 VCC.n5138 0.00228571
R58880 VCC.n5340 VCC.n5100 0.00228571
R58881 VCC.n5466 VCC.n5465 0.00228571
R58882 VCC.n5477 VCC.n5032 0.00228571
R58883 VCC.n5489 VCC.n5026 0.00228571
R58884 VCC.n5510 VCC.n5509 0.00228571
R58885 VCC.n5490 VCC.n5024 0.00228571
R58886 VCC.n6032 VCC.n6031 0.00228571
R58887 VCC.n6028 VCC.n6024 0.00228571
R58888 VCC.n6041 VCC.n5582 0.00228571
R58889 VCC.n6060 VCC.n5570 0.00228571
R58890 VCC.n6043 VCC.n6042 0.00228571
R58891 VCC.n5897 VCC.n5657 0.00228571
R58892 VCC.n5761 VCC.n5760 0.00228571
R58893 VCC.n5768 VCC.n5766 0.00228571
R58894 VCC.n5708 VCC.n5707 0.00228571
R58895 VCC.n5824 VCC.n5696 0.00228571
R58896 VCC.n6312 VCC.n6311 0.00228571
R58897 VCC.n6319 VCC.n6317 0.00228571
R58898 VCC.n6259 VCC.n6258 0.00228571
R58899 VCC.n6375 VCC.n6247 0.00228571
R58900 VCC.n6449 VCC.n6209 0.00228571
R58901 VCC.n6575 VCC.n6574 0.00228571
R58902 VCC.n6586 VCC.n6141 0.00228571
R58903 VCC.n6598 VCC.n6135 0.00228571
R58904 VCC.n6619 VCC.n6618 0.00228571
R58905 VCC.n6599 VCC.n6133 0.00228571
R58906 VCC.n7141 VCC.n7140 0.00228571
R58907 VCC.n7137 VCC.n7133 0.00228571
R58908 VCC.n7150 VCC.n6691 0.00228571
R58909 VCC.n7169 VCC.n6679 0.00228571
R58910 VCC.n7152 VCC.n7151 0.00228571
R58911 VCC.n7006 VCC.n6766 0.00228571
R58912 VCC.n6870 VCC.n6869 0.00228571
R58913 VCC.n6877 VCC.n6875 0.00228571
R58914 VCC.n6817 VCC.n6816 0.00228571
R58915 VCC.n6933 VCC.n6805 0.00228571
R58916 VCC.n7421 VCC.n7420 0.00228571
R58917 VCC.n7428 VCC.n7426 0.00228571
R58918 VCC.n7368 VCC.n7367 0.00228571
R58919 VCC.n7484 VCC.n7356 0.00228571
R58920 VCC.n7558 VCC.n7318 0.00228571
R58921 VCC.n7684 VCC.n7683 0.00228571
R58922 VCC.n7695 VCC.n7250 0.00228571
R58923 VCC.n7707 VCC.n7244 0.00228571
R58924 VCC.n7728 VCC.n7727 0.00228571
R58925 VCC.n7708 VCC.n7242 0.00228571
R58926 VCC.n8250 VCC.n8249 0.00228571
R58927 VCC.n8246 VCC.n8242 0.00228571
R58928 VCC.n8259 VCC.n7800 0.00228571
R58929 VCC.n8278 VCC.n7788 0.00228571
R58930 VCC.n8261 VCC.n8260 0.00228571
R58931 VCC.n8115 VCC.n7875 0.00228571
R58932 VCC.n7979 VCC.n7978 0.00228571
R58933 VCC.n7986 VCC.n7984 0.00228571
R58934 VCC.n7926 VCC.n7925 0.00228571
R58935 VCC.n8042 VCC.n7914 0.00228571
R58936 VCC.n8667 VCC.n8427 0.00228571
R58937 VCC.n8793 VCC.n8792 0.00228571
R58938 VCC.n8804 VCC.n8359 0.00228571
R58939 VCC.n8816 VCC.n8353 0.00228571
R58940 VCC.n8837 VCC.n8836 0.00228571
R58941 VCC.n8817 VCC.n8351 0.00228571
R58942 VCC.n8530 VCC.n8529 0.00228571
R58943 VCC.n8537 VCC.n8535 0.00228571
R58944 VCC.n8477 VCC.n8476 0.00228571
R58945 VCC.n8593 VCC.n8465 0.00228571
R58946 VCC.n9359 VCC.n9358 0.00228571
R58947 VCC.n9355 VCC.n9351 0.00228571
R58948 VCC.n9368 VCC.n8909 0.00228571
R58949 VCC.n9387 VCC.n8897 0.00228571
R58950 VCC.n9370 VCC.n9369 0.00228571
R58951 VCC.n9224 VCC.n8984 0.00228571
R58952 VCC.n9088 VCC.n9087 0.00228571
R58953 VCC.n9095 VCC.n9093 0.00228571
R58954 VCC.n9035 VCC.n9034 0.00228571
R58955 VCC.n9151 VCC.n9023 0.00228571
R58956 VCC.n9639 VCC.n9638 0.00228571
R58957 VCC.n9646 VCC.n9644 0.00228571
R58958 VCC.n9586 VCC.n9585 0.00228571
R58959 VCC.n9702 VCC.n9574 0.00228571
R58960 VCC.n9776 VCC.n9536 0.00228571
R58961 VCC.n9902 VCC.n9901 0.00228571
R58962 VCC.n9913 VCC.n9468 0.00228571
R58963 VCC.n9925 VCC.n9462 0.00228571
R58964 VCC.n9946 VCC.n9945 0.00228571
R58965 VCC.n9926 VCC.n9460 0.00228571
R58966 VCC.n10467 VCC.n10466 0.00228571
R58967 VCC.n10463 VCC.n10459 0.00228571
R58968 VCC.n10476 VCC.n10017 0.00228571
R58969 VCC.n10495 VCC.n10005 0.00228571
R58970 VCC.n10478 VCC.n10477 0.00228571
R58971 VCC.n10332 VCC.n10092 0.00228571
R58972 VCC.n10196 VCC.n10195 0.00228571
R58973 VCC.n10203 VCC.n10201 0.00228571
R58974 VCC.n10143 VCC.n10142 0.00228571
R58975 VCC.n10259 VCC.n10131 0.00228571
R58976 VCC.n10746 VCC.n10745 0.00228571
R58977 VCC.n10753 VCC.n10751 0.00228571
R58978 VCC.n10693 VCC.n10692 0.00228571
R58979 VCC.n10809 VCC.n10681 0.00228571
R58980 VCC.n10883 VCC.n10643 0.00228571
R58981 VCC.n11009 VCC.n11008 0.00228571
R58982 VCC.n11020 VCC.n10575 0.00228571
R58983 VCC.n11032 VCC.n10569 0.00228571
R58984 VCC.n11053 VCC.n11052 0.00228571
R58985 VCC.n11033 VCC.n10567 0.00228571
R58986 VCC.n11574 VCC.n11573 0.00228571
R58987 VCC.n11570 VCC.n11566 0.00228571
R58988 VCC.n11583 VCC.n11124 0.00228571
R58989 VCC.n11602 VCC.n11112 0.00228571
R58990 VCC.n11585 VCC.n11584 0.00228571
R58991 VCC.n11439 VCC.n11199 0.00228571
R58992 VCC.n11303 VCC.n11302 0.00228571
R58993 VCC.n11310 VCC.n11308 0.00228571
R58994 VCC.n11250 VCC.n11249 0.00228571
R58995 VCC.n11366 VCC.n11238 0.00228571
R58996 VCC.n11853 VCC.n11852 0.00228571
R58997 VCC.n11860 VCC.n11858 0.00228571
R58998 VCC.n11800 VCC.n11799 0.00228571
R58999 VCC.n11916 VCC.n11788 0.00228571
R59000 VCC.n11990 VCC.n11750 0.00228571
R59001 VCC.n12116 VCC.n12115 0.00228571
R59002 VCC.n12127 VCC.n11682 0.00228571
R59003 VCC.n12139 VCC.n11676 0.00228571
R59004 VCC.n12160 VCC.n12159 0.00228571
R59005 VCC.n12140 VCC.n11674 0.00228571
R59006 VCC.n12681 VCC.n12680 0.00228571
R59007 VCC.n12677 VCC.n12673 0.00228571
R59008 VCC.n12690 VCC.n12231 0.00228571
R59009 VCC.n12709 VCC.n12219 0.00228571
R59010 VCC.n12692 VCC.n12691 0.00228571
R59011 VCC.n12546 VCC.n12306 0.00228571
R59012 VCC.n12410 VCC.n12409 0.00228571
R59013 VCC.n12417 VCC.n12415 0.00228571
R59014 VCC.n12357 VCC.n12356 0.00228571
R59015 VCC.n12473 VCC.n12345 0.00228571
R59016 VCC.n12960 VCC.n12959 0.00228571
R59017 VCC.n12967 VCC.n12965 0.00228571
R59018 VCC.n12907 VCC.n12906 0.00228571
R59019 VCC.n13023 VCC.n12895 0.00228571
R59020 VCC.n13097 VCC.n12857 0.00228571
R59021 VCC.n13223 VCC.n13222 0.00228571
R59022 VCC.n13234 VCC.n12789 0.00228571
R59023 VCC.n13246 VCC.n12783 0.00228571
R59024 VCC.n13267 VCC.n13266 0.00228571
R59025 VCC.n13247 VCC.n12781 0.00228571
R59026 VCC.n13788 VCC.n13787 0.00228571
R59027 VCC.n13784 VCC.n13780 0.00228571
R59028 VCC.n13797 VCC.n13338 0.00228571
R59029 VCC.n13816 VCC.n13326 0.00228571
R59030 VCC.n13799 VCC.n13798 0.00228571
R59031 VCC.n13653 VCC.n13413 0.00228571
R59032 VCC.n13517 VCC.n13516 0.00228571
R59033 VCC.n13524 VCC.n13522 0.00228571
R59034 VCC.n13464 VCC.n13463 0.00228571
R59035 VCC.n13580 VCC.n13452 0.00228571
R59036 VCC.n14067 VCC.n14066 0.00228571
R59037 VCC.n14074 VCC.n14072 0.00228571
R59038 VCC.n14014 VCC.n14013 0.00228571
R59039 VCC.n14130 VCC.n14002 0.00228571
R59040 VCC.n14204 VCC.n13964 0.00228571
R59041 VCC.n14330 VCC.n14329 0.00228571
R59042 VCC.n14341 VCC.n13896 0.00228571
R59043 VCC.n14353 VCC.n13890 0.00228571
R59044 VCC.n14374 VCC.n14373 0.00228571
R59045 VCC.n14354 VCC.n13888 0.00228571
R59046 VCC.n14895 VCC.n14894 0.00228571
R59047 VCC.n14891 VCC.n14887 0.00228571
R59048 VCC.n14904 VCC.n14445 0.00228571
R59049 VCC.n14923 VCC.n14433 0.00228571
R59050 VCC.n14906 VCC.n14905 0.00228571
R59051 VCC.n14760 VCC.n14520 0.00228571
R59052 VCC.n14624 VCC.n14623 0.00228571
R59053 VCC.n14631 VCC.n14629 0.00228571
R59054 VCC.n14571 VCC.n14570 0.00228571
R59055 VCC.n14687 VCC.n14559 0.00228571
R59056 VCC.n15174 VCC.n15173 0.00228571
R59057 VCC.n15181 VCC.n15179 0.00228571
R59058 VCC.n15121 VCC.n15120 0.00228571
R59059 VCC.n15237 VCC.n15109 0.00228571
R59060 VCC.n15311 VCC.n15071 0.00228571
R59061 VCC.n15437 VCC.n15436 0.00228571
R59062 VCC.n15448 VCC.n15003 0.00228571
R59063 VCC.n15460 VCC.n14997 0.00228571
R59064 VCC.n15481 VCC.n15480 0.00228571
R59065 VCC.n15461 VCC.n14995 0.00228571
R59066 VCC.n16002 VCC.n16001 0.00228571
R59067 VCC.n15998 VCC.n15994 0.00228571
R59068 VCC.n16011 VCC.n15552 0.00228571
R59069 VCC.n16030 VCC.n15540 0.00228571
R59070 VCC.n16013 VCC.n16012 0.00228571
R59071 VCC.n15867 VCC.n15627 0.00228571
R59072 VCC.n15731 VCC.n15730 0.00228571
R59073 VCC.n15738 VCC.n15736 0.00228571
R59074 VCC.n15678 VCC.n15677 0.00228571
R59075 VCC.n15794 VCC.n15666 0.00228571
R59076 VCC.n16281 VCC.n16280 0.00228571
R59077 VCC.n16288 VCC.n16286 0.00228571
R59078 VCC.n16228 VCC.n16227 0.00228571
R59079 VCC.n16344 VCC.n16216 0.00228571
R59080 VCC.n16418 VCC.n16178 0.00228571
R59081 VCC.n16544 VCC.n16543 0.00228571
R59082 VCC.n16555 VCC.n16110 0.00228571
R59083 VCC.n16567 VCC.n16104 0.00228571
R59084 VCC.n16588 VCC.n16587 0.00228571
R59085 VCC.n16568 VCC.n16102 0.00228571
R59086 VCC.n17109 VCC.n17108 0.00228571
R59087 VCC.n17105 VCC.n17101 0.00228571
R59088 VCC.n17118 VCC.n16659 0.00228571
R59089 VCC.n17137 VCC.n16647 0.00228571
R59090 VCC.n17120 VCC.n17119 0.00228571
R59091 VCC.n16974 VCC.n16734 0.00228571
R59092 VCC.n16838 VCC.n16837 0.00228571
R59093 VCC.n16845 VCC.n16843 0.00228571
R59094 VCC.n16785 VCC.n16784 0.00228571
R59095 VCC.n16901 VCC.n16773 0.00228571
R59096 VCC.n17338 VCC.n17285 0.00228571
R59097 VCC.n17464 VCC.n17463 0.00228571
R59098 VCC.n17475 VCC.n17217 0.00228571
R59099 VCC.n17487 VCC.n17211 0.00228571
R59100 VCC.n17508 VCC.n17507 0.00228571
R59101 VCC.n17488 VCC.n17209 0.00228571
R59102 VCC.n217 VCC.n188 0.00217857
R59103 VCC.n218 VCC.n173 0.00217857
R59104 VCC.n307 VCC.n131 0.00217857
R59105 VCC.n308 VCC.n127 0.00217857
R59106 VCC.n317 VCC.n316 0.00217857
R59107 VCC.n346 VCC.n114 0.00217857
R59108 VCC.n442 VCC.n70 0.00217857
R59109 VCC.n443 VCC.n66 0.00217857
R59110 VCC.n460 VCC.n62 0.00217857
R59111 VCC.n461 VCC.n49 0.00217857
R59112 VCC.n536 VCC.n13 0.00217857
R59113 VCC.n537 VCC.n0 0.00217857
R59114 VCC.n769 VCC.n740 0.00217857
R59115 VCC.n770 VCC.n725 0.00217857
R59116 VCC.n859 VCC.n683 0.00217857
R59117 VCC.n860 VCC.n679 0.00217857
R59118 VCC.n869 VCC.n868 0.00217857
R59119 VCC.n898 VCC.n666 0.00217857
R59120 VCC.n994 VCC.n622 0.00217857
R59121 VCC.n995 VCC.n618 0.00217857
R59122 VCC.n1012 VCC.n614 0.00217857
R59123 VCC.n1013 VCC.n601 0.00217857
R59124 VCC.n1088 VCC.n565 0.00217857
R59125 VCC.n1089 VCC.n554 0.00217857
R59126 VCC.n1327 VCC.n1298 0.00217857
R59127 VCC.n1328 VCC.n1283 0.00217857
R59128 VCC.n1417 VCC.n1241 0.00217857
R59129 VCC.n1418 VCC.n1237 0.00217857
R59130 VCC.n1427 VCC.n1426 0.00217857
R59131 VCC.n1455 VCC.n1223 0.00217857
R59132 VCC.n1552 VCC.n1179 0.00217857
R59133 VCC.n1553 VCC.n1175 0.00217857
R59134 VCC.n1571 VCC.n1171 0.00217857
R59135 VCC.n1572 VCC.n1154 0.00217857
R59136 VCC.n1635 VCC.n1126 0.00217857
R59137 VCC.n1636 VCC.n1108 0.00217857
R59138 VCC.n1878 VCC.n1849 0.00217857
R59139 VCC.n1879 VCC.n1834 0.00217857
R59140 VCC.n1968 VCC.n1792 0.00217857
R59141 VCC.n1969 VCC.n1788 0.00217857
R59142 VCC.n1978 VCC.n1977 0.00217857
R59143 VCC.n2007 VCC.n1775 0.00217857
R59144 VCC.n2103 VCC.n1731 0.00217857
R59145 VCC.n2104 VCC.n1727 0.00217857
R59146 VCC.n2121 VCC.n1723 0.00217857
R59147 VCC.n2122 VCC.n1710 0.00217857
R59148 VCC.n2197 VCC.n1674 0.00217857
R59149 VCC.n2198 VCC.n1663 0.00217857
R59150 VCC.n2436 VCC.n2407 0.00217857
R59151 VCC.n2437 VCC.n2392 0.00217857
R59152 VCC.n2526 VCC.n2350 0.00217857
R59153 VCC.n2527 VCC.n2346 0.00217857
R59154 VCC.n2536 VCC.n2535 0.00217857
R59155 VCC.n2564 VCC.n2332 0.00217857
R59156 VCC.n2661 VCC.n2288 0.00217857
R59157 VCC.n2662 VCC.n2284 0.00217857
R59158 VCC.n2680 VCC.n2280 0.00217857
R59159 VCC.n2681 VCC.n2263 0.00217857
R59160 VCC.n2744 VCC.n2235 0.00217857
R59161 VCC.n2745 VCC.n2217 0.00217857
R59162 VCC.n2987 VCC.n2958 0.00217857
R59163 VCC.n2988 VCC.n2943 0.00217857
R59164 VCC.n3077 VCC.n2901 0.00217857
R59165 VCC.n3078 VCC.n2897 0.00217857
R59166 VCC.n3087 VCC.n3086 0.00217857
R59167 VCC.n3116 VCC.n2884 0.00217857
R59168 VCC.n3212 VCC.n2840 0.00217857
R59169 VCC.n3213 VCC.n2836 0.00217857
R59170 VCC.n3230 VCC.n2832 0.00217857
R59171 VCC.n3231 VCC.n2819 0.00217857
R59172 VCC.n3306 VCC.n2783 0.00217857
R59173 VCC.n3307 VCC.n2772 0.00217857
R59174 VCC.n3545 VCC.n3516 0.00217857
R59175 VCC.n3546 VCC.n3501 0.00217857
R59176 VCC.n3635 VCC.n3459 0.00217857
R59177 VCC.n3636 VCC.n3455 0.00217857
R59178 VCC.n3645 VCC.n3644 0.00217857
R59179 VCC.n3673 VCC.n3441 0.00217857
R59180 VCC.n3770 VCC.n3397 0.00217857
R59181 VCC.n3771 VCC.n3393 0.00217857
R59182 VCC.n3789 VCC.n3389 0.00217857
R59183 VCC.n3790 VCC.n3372 0.00217857
R59184 VCC.n3853 VCC.n3344 0.00217857
R59185 VCC.n3854 VCC.n3326 0.00217857
R59186 VCC.n4096 VCC.n4067 0.00217857
R59187 VCC.n4097 VCC.n4052 0.00217857
R59188 VCC.n4186 VCC.n4010 0.00217857
R59189 VCC.n4187 VCC.n4006 0.00217857
R59190 VCC.n4196 VCC.n4195 0.00217857
R59191 VCC.n4225 VCC.n3993 0.00217857
R59192 VCC.n4321 VCC.n3949 0.00217857
R59193 VCC.n4322 VCC.n3945 0.00217857
R59194 VCC.n4339 VCC.n3941 0.00217857
R59195 VCC.n4340 VCC.n3928 0.00217857
R59196 VCC.n4415 VCC.n3892 0.00217857
R59197 VCC.n4416 VCC.n3881 0.00217857
R59198 VCC.n4654 VCC.n4625 0.00217857
R59199 VCC.n4655 VCC.n4610 0.00217857
R59200 VCC.n4744 VCC.n4568 0.00217857
R59201 VCC.n4745 VCC.n4564 0.00217857
R59202 VCC.n4754 VCC.n4753 0.00217857
R59203 VCC.n4782 VCC.n4550 0.00217857
R59204 VCC.n4879 VCC.n4506 0.00217857
R59205 VCC.n4880 VCC.n4502 0.00217857
R59206 VCC.n4898 VCC.n4498 0.00217857
R59207 VCC.n4899 VCC.n4481 0.00217857
R59208 VCC.n4962 VCC.n4453 0.00217857
R59209 VCC.n4963 VCC.n4435 0.00217857
R59210 VCC.n5205 VCC.n5176 0.00217857
R59211 VCC.n5206 VCC.n5161 0.00217857
R59212 VCC.n5295 VCC.n5119 0.00217857
R59213 VCC.n5296 VCC.n5115 0.00217857
R59214 VCC.n5305 VCC.n5304 0.00217857
R59215 VCC.n5334 VCC.n5102 0.00217857
R59216 VCC.n5430 VCC.n5058 0.00217857
R59217 VCC.n5431 VCC.n5054 0.00217857
R59218 VCC.n5448 VCC.n5050 0.00217857
R59219 VCC.n5449 VCC.n5037 0.00217857
R59220 VCC.n5524 VCC.n5001 0.00217857
R59221 VCC.n5525 VCC.n4990 0.00217857
R59222 VCC.n5763 VCC.n5734 0.00217857
R59223 VCC.n5764 VCC.n5719 0.00217857
R59224 VCC.n5853 VCC.n5677 0.00217857
R59225 VCC.n5854 VCC.n5673 0.00217857
R59226 VCC.n5863 VCC.n5862 0.00217857
R59227 VCC.n5891 VCC.n5659 0.00217857
R59228 VCC.n5988 VCC.n5615 0.00217857
R59229 VCC.n5989 VCC.n5611 0.00217857
R59230 VCC.n6007 VCC.n5607 0.00217857
R59231 VCC.n6008 VCC.n5590 0.00217857
R59232 VCC.n6071 VCC.n5562 0.00217857
R59233 VCC.n6072 VCC.n5544 0.00217857
R59234 VCC.n6314 VCC.n6285 0.00217857
R59235 VCC.n6315 VCC.n6270 0.00217857
R59236 VCC.n6404 VCC.n6228 0.00217857
R59237 VCC.n6405 VCC.n6224 0.00217857
R59238 VCC.n6414 VCC.n6413 0.00217857
R59239 VCC.n6443 VCC.n6211 0.00217857
R59240 VCC.n6539 VCC.n6167 0.00217857
R59241 VCC.n6540 VCC.n6163 0.00217857
R59242 VCC.n6557 VCC.n6159 0.00217857
R59243 VCC.n6558 VCC.n6146 0.00217857
R59244 VCC.n6633 VCC.n6110 0.00217857
R59245 VCC.n6634 VCC.n6099 0.00217857
R59246 VCC.n6872 VCC.n6843 0.00217857
R59247 VCC.n6873 VCC.n6828 0.00217857
R59248 VCC.n6962 VCC.n6786 0.00217857
R59249 VCC.n6963 VCC.n6782 0.00217857
R59250 VCC.n6972 VCC.n6971 0.00217857
R59251 VCC.n7000 VCC.n6768 0.00217857
R59252 VCC.n7097 VCC.n6724 0.00217857
R59253 VCC.n7098 VCC.n6720 0.00217857
R59254 VCC.n7116 VCC.n6716 0.00217857
R59255 VCC.n7117 VCC.n6699 0.00217857
R59256 VCC.n7180 VCC.n6671 0.00217857
R59257 VCC.n7181 VCC.n6653 0.00217857
R59258 VCC.n7423 VCC.n7394 0.00217857
R59259 VCC.n7424 VCC.n7379 0.00217857
R59260 VCC.n7513 VCC.n7337 0.00217857
R59261 VCC.n7514 VCC.n7333 0.00217857
R59262 VCC.n7523 VCC.n7522 0.00217857
R59263 VCC.n7552 VCC.n7320 0.00217857
R59264 VCC.n7648 VCC.n7276 0.00217857
R59265 VCC.n7649 VCC.n7272 0.00217857
R59266 VCC.n7666 VCC.n7268 0.00217857
R59267 VCC.n7667 VCC.n7255 0.00217857
R59268 VCC.n7742 VCC.n7219 0.00217857
R59269 VCC.n7743 VCC.n7208 0.00217857
R59270 VCC.n7981 VCC.n7952 0.00217857
R59271 VCC.n7982 VCC.n7937 0.00217857
R59272 VCC.n8071 VCC.n7895 0.00217857
R59273 VCC.n8072 VCC.n7891 0.00217857
R59274 VCC.n8081 VCC.n8080 0.00217857
R59275 VCC.n8109 VCC.n7877 0.00217857
R59276 VCC.n8206 VCC.n7833 0.00217857
R59277 VCC.n8207 VCC.n7829 0.00217857
R59278 VCC.n8225 VCC.n7825 0.00217857
R59279 VCC.n8226 VCC.n7808 0.00217857
R59280 VCC.n8289 VCC.n7780 0.00217857
R59281 VCC.n8290 VCC.n7762 0.00217857
R59282 VCC.n8632 VCC.n8631 0.00217857
R59283 VCC.n8661 VCC.n8429 0.00217857
R59284 VCC.n8757 VCC.n8385 0.00217857
R59285 VCC.n8758 VCC.n8381 0.00217857
R59286 VCC.n8775 VCC.n8377 0.00217857
R59287 VCC.n8776 VCC.n8364 0.00217857
R59288 VCC.n8851 VCC.n8328 0.00217857
R59289 VCC.n8852 VCC.n8317 0.00217857
R59290 VCC.n9090 VCC.n9061 0.00217857
R59291 VCC.n9091 VCC.n9046 0.00217857
R59292 VCC.n9180 VCC.n9004 0.00217857
R59293 VCC.n9181 VCC.n9000 0.00217857
R59294 VCC.n9190 VCC.n9189 0.00217857
R59295 VCC.n9218 VCC.n8986 0.00217857
R59296 VCC.n9315 VCC.n8942 0.00217857
R59297 VCC.n9316 VCC.n8938 0.00217857
R59298 VCC.n9334 VCC.n8934 0.00217857
R59299 VCC.n9335 VCC.n8917 0.00217857
R59300 VCC.n9398 VCC.n8889 0.00217857
R59301 VCC.n9399 VCC.n8871 0.00217857
R59302 VCC.n9641 VCC.n9612 0.00217857
R59303 VCC.n9642 VCC.n9597 0.00217857
R59304 VCC.n9731 VCC.n9555 0.00217857
R59305 VCC.n9732 VCC.n9551 0.00217857
R59306 VCC.n9741 VCC.n9740 0.00217857
R59307 VCC.n9770 VCC.n9538 0.00217857
R59308 VCC.n9866 VCC.n9494 0.00217857
R59309 VCC.n9867 VCC.n9490 0.00217857
R59310 VCC.n9884 VCC.n9486 0.00217857
R59311 VCC.n9885 VCC.n9473 0.00217857
R59312 VCC.n9960 VCC.n9437 0.00217857
R59313 VCC.n9961 VCC.n9426 0.00217857
R59314 VCC.n10198 VCC.n10169 0.00217857
R59315 VCC.n10199 VCC.n10154 0.00217857
R59316 VCC.n10288 VCC.n10112 0.00217857
R59317 VCC.n10289 VCC.n10108 0.00217857
R59318 VCC.n10298 VCC.n10297 0.00217857
R59319 VCC.n10326 VCC.n10094 0.00217857
R59320 VCC.n10423 VCC.n10050 0.00217857
R59321 VCC.n10424 VCC.n10046 0.00217857
R59322 VCC.n10442 VCC.n10042 0.00217857
R59323 VCC.n10443 VCC.n10025 0.00217857
R59324 VCC.n10506 VCC.n9997 0.00217857
R59325 VCC.n10507 VCC.n9979 0.00217857
R59326 VCC.n10748 VCC.n10719 0.00217857
R59327 VCC.n10749 VCC.n10704 0.00217857
R59328 VCC.n10838 VCC.n10662 0.00217857
R59329 VCC.n10839 VCC.n10658 0.00217857
R59330 VCC.n10848 VCC.n10847 0.00217857
R59331 VCC.n10877 VCC.n10645 0.00217857
R59332 VCC.n10973 VCC.n10601 0.00217857
R59333 VCC.n10974 VCC.n10597 0.00217857
R59334 VCC.n10991 VCC.n10593 0.00217857
R59335 VCC.n10992 VCC.n10580 0.00217857
R59336 VCC.n11067 VCC.n10544 0.00217857
R59337 VCC.n11068 VCC.n10533 0.00217857
R59338 VCC.n11305 VCC.n11276 0.00217857
R59339 VCC.n11306 VCC.n11261 0.00217857
R59340 VCC.n11395 VCC.n11219 0.00217857
R59341 VCC.n11396 VCC.n11215 0.00217857
R59342 VCC.n11405 VCC.n11404 0.00217857
R59343 VCC.n11433 VCC.n11201 0.00217857
R59344 VCC.n11530 VCC.n11157 0.00217857
R59345 VCC.n11531 VCC.n11153 0.00217857
R59346 VCC.n11549 VCC.n11149 0.00217857
R59347 VCC.n11550 VCC.n11132 0.00217857
R59348 VCC.n11613 VCC.n11104 0.00217857
R59349 VCC.n11614 VCC.n11086 0.00217857
R59350 VCC.n11855 VCC.n11826 0.00217857
R59351 VCC.n11856 VCC.n11811 0.00217857
R59352 VCC.n11945 VCC.n11769 0.00217857
R59353 VCC.n11946 VCC.n11765 0.00217857
R59354 VCC.n11955 VCC.n11954 0.00217857
R59355 VCC.n11984 VCC.n11752 0.00217857
R59356 VCC.n12080 VCC.n11708 0.00217857
R59357 VCC.n12081 VCC.n11704 0.00217857
R59358 VCC.n12098 VCC.n11700 0.00217857
R59359 VCC.n12099 VCC.n11687 0.00217857
R59360 VCC.n12174 VCC.n11651 0.00217857
R59361 VCC.n12175 VCC.n11640 0.00217857
R59362 VCC.n12412 VCC.n12383 0.00217857
R59363 VCC.n12413 VCC.n12368 0.00217857
R59364 VCC.n12502 VCC.n12326 0.00217857
R59365 VCC.n12503 VCC.n12322 0.00217857
R59366 VCC.n12512 VCC.n12511 0.00217857
R59367 VCC.n12540 VCC.n12308 0.00217857
R59368 VCC.n12637 VCC.n12264 0.00217857
R59369 VCC.n12638 VCC.n12260 0.00217857
R59370 VCC.n12656 VCC.n12256 0.00217857
R59371 VCC.n12657 VCC.n12239 0.00217857
R59372 VCC.n12720 VCC.n12211 0.00217857
R59373 VCC.n12721 VCC.n12193 0.00217857
R59374 VCC.n12962 VCC.n12933 0.00217857
R59375 VCC.n12963 VCC.n12918 0.00217857
R59376 VCC.n13052 VCC.n12876 0.00217857
R59377 VCC.n13053 VCC.n12872 0.00217857
R59378 VCC.n13062 VCC.n13061 0.00217857
R59379 VCC.n13091 VCC.n12859 0.00217857
R59380 VCC.n13187 VCC.n12815 0.00217857
R59381 VCC.n13188 VCC.n12811 0.00217857
R59382 VCC.n13205 VCC.n12807 0.00217857
R59383 VCC.n13206 VCC.n12794 0.00217857
R59384 VCC.n13281 VCC.n12758 0.00217857
R59385 VCC.n13282 VCC.n12747 0.00217857
R59386 VCC.n13519 VCC.n13490 0.00217857
R59387 VCC.n13520 VCC.n13475 0.00217857
R59388 VCC.n13609 VCC.n13433 0.00217857
R59389 VCC.n13610 VCC.n13429 0.00217857
R59390 VCC.n13619 VCC.n13618 0.00217857
R59391 VCC.n13647 VCC.n13415 0.00217857
R59392 VCC.n13744 VCC.n13371 0.00217857
R59393 VCC.n13745 VCC.n13367 0.00217857
R59394 VCC.n13763 VCC.n13363 0.00217857
R59395 VCC.n13764 VCC.n13346 0.00217857
R59396 VCC.n13827 VCC.n13318 0.00217857
R59397 VCC.n13828 VCC.n13300 0.00217857
R59398 VCC.n14069 VCC.n14040 0.00217857
R59399 VCC.n14070 VCC.n14025 0.00217857
R59400 VCC.n14159 VCC.n13983 0.00217857
R59401 VCC.n14160 VCC.n13979 0.00217857
R59402 VCC.n14169 VCC.n14168 0.00217857
R59403 VCC.n14198 VCC.n13966 0.00217857
R59404 VCC.n14294 VCC.n13922 0.00217857
R59405 VCC.n14295 VCC.n13918 0.00217857
R59406 VCC.n14312 VCC.n13914 0.00217857
R59407 VCC.n14313 VCC.n13901 0.00217857
R59408 VCC.n14388 VCC.n13865 0.00217857
R59409 VCC.n14389 VCC.n13854 0.00217857
R59410 VCC.n14626 VCC.n14597 0.00217857
R59411 VCC.n14627 VCC.n14582 0.00217857
R59412 VCC.n14716 VCC.n14540 0.00217857
R59413 VCC.n14717 VCC.n14536 0.00217857
R59414 VCC.n14726 VCC.n14725 0.00217857
R59415 VCC.n14754 VCC.n14522 0.00217857
R59416 VCC.n14851 VCC.n14478 0.00217857
R59417 VCC.n14852 VCC.n14474 0.00217857
R59418 VCC.n14870 VCC.n14470 0.00217857
R59419 VCC.n14871 VCC.n14453 0.00217857
R59420 VCC.n14934 VCC.n14425 0.00217857
R59421 VCC.n14935 VCC.n14407 0.00217857
R59422 VCC.n15176 VCC.n15147 0.00217857
R59423 VCC.n15177 VCC.n15132 0.00217857
R59424 VCC.n15266 VCC.n15090 0.00217857
R59425 VCC.n15267 VCC.n15086 0.00217857
R59426 VCC.n15276 VCC.n15275 0.00217857
R59427 VCC.n15305 VCC.n15073 0.00217857
R59428 VCC.n15401 VCC.n15029 0.00217857
R59429 VCC.n15402 VCC.n15025 0.00217857
R59430 VCC.n15419 VCC.n15021 0.00217857
R59431 VCC.n15420 VCC.n15008 0.00217857
R59432 VCC.n15495 VCC.n14972 0.00217857
R59433 VCC.n15496 VCC.n14961 0.00217857
R59434 VCC.n15733 VCC.n15704 0.00217857
R59435 VCC.n15734 VCC.n15689 0.00217857
R59436 VCC.n15823 VCC.n15647 0.00217857
R59437 VCC.n15824 VCC.n15643 0.00217857
R59438 VCC.n15833 VCC.n15832 0.00217857
R59439 VCC.n15861 VCC.n15629 0.00217857
R59440 VCC.n15958 VCC.n15585 0.00217857
R59441 VCC.n15959 VCC.n15581 0.00217857
R59442 VCC.n15977 VCC.n15577 0.00217857
R59443 VCC.n15978 VCC.n15560 0.00217857
R59444 VCC.n16041 VCC.n15532 0.00217857
R59445 VCC.n16042 VCC.n15514 0.00217857
R59446 VCC.n16283 VCC.n16254 0.00217857
R59447 VCC.n16284 VCC.n16239 0.00217857
R59448 VCC.n16373 VCC.n16197 0.00217857
R59449 VCC.n16374 VCC.n16193 0.00217857
R59450 VCC.n16383 VCC.n16382 0.00217857
R59451 VCC.n16412 VCC.n16180 0.00217857
R59452 VCC.n16508 VCC.n16136 0.00217857
R59453 VCC.n16509 VCC.n16132 0.00217857
R59454 VCC.n16526 VCC.n16128 0.00217857
R59455 VCC.n16527 VCC.n16115 0.00217857
R59456 VCC.n16602 VCC.n16079 0.00217857
R59457 VCC.n16603 VCC.n16068 0.00217857
R59458 VCC.n16840 VCC.n16811 0.00217857
R59459 VCC.n16841 VCC.n16796 0.00217857
R59460 VCC.n16930 VCC.n16754 0.00217857
R59461 VCC.n16931 VCC.n16750 0.00217857
R59462 VCC.n16940 VCC.n16939 0.00217857
R59463 VCC.n16968 VCC.n16736 0.00217857
R59464 VCC.n17065 VCC.n16692 0.00217857
R59465 VCC.n17066 VCC.n16688 0.00217857
R59466 VCC.n17084 VCC.n16684 0.00217857
R59467 VCC.n17085 VCC.n16667 0.00217857
R59468 VCC.n17148 VCC.n16639 0.00217857
R59469 VCC.n17149 VCC.n16621 0.00217857
R59470 VCC.n17303 VCC.n17302 0.00217857
R59471 VCC.n17332 VCC.n17287 0.00217857
R59472 VCC.n17428 VCC.n17243 0.00217857
R59473 VCC.n17429 VCC.n17239 0.00217857
R59474 VCC.n17446 VCC.n17235 0.00217857
R59475 VCC.n17447 VCC.n17222 0.00217857
R59476 VCC.n17522 VCC.n17186 0.00217857
R59477 VCC.n17523 VCC.n17175 0.00217857
R59478 VCC.n8532 VCC.n8503 0.00216667
R59479 VCC.n8533 VCC.n8488 0.00216667
R59480 VCC.n8622 VCC.n8446 0.00216667
R59481 VCC.n8623 VCC.n8442 0.00216667
R59482 VCC.n214 VCC.n193 0.00139286
R59483 VCC.n237 VCC.n236 0.00139286
R59484 VCC.n254 VCC.n253 0.00139286
R59485 VCC.n294 VCC.n129 0.00139286
R59486 VCC.n252 VCC.n167 0.00139286
R59487 VCC.n350 VCC.n104 0.00139286
R59488 VCC.n405 VCC.n90 0.00139286
R59489 VCC.n532 VCC.n19 0.00139286
R59490 VCC.n543 VCC.n8 0.00139286
R59491 VCC.n766 VCC.n745 0.00139286
R59492 VCC.n789 VCC.n788 0.00139286
R59493 VCC.n806 VCC.n805 0.00139286
R59494 VCC.n846 VCC.n681 0.00139286
R59495 VCC.n804 VCC.n719 0.00139286
R59496 VCC.n902 VCC.n656 0.00139286
R59497 VCC.n957 VCC.n642 0.00139286
R59498 VCC.n1084 VCC.n571 0.00139286
R59499 VCC.n1097 VCC.n562 0.00139286
R59500 VCC.n1647 VCC.n1646 0.00139286
R59501 VCC.n1125 VCC.n1122 0.00139286
R59502 VCC.n1459 VCC.n1213 0.00139286
R59503 VCC.n1514 VCC.n1199 0.00139286
R59504 VCC.n1324 VCC.n1303 0.00139286
R59505 VCC.n1347 VCC.n1346 0.00139286
R59506 VCC.n1364 VCC.n1363 0.00139286
R59507 VCC.n1404 VCC.n1239 0.00139286
R59508 VCC.n1362 VCC.n1277 0.00139286
R59509 VCC.n1875 VCC.n1854 0.00139286
R59510 VCC.n1898 VCC.n1897 0.00139286
R59511 VCC.n1915 VCC.n1914 0.00139286
R59512 VCC.n1955 VCC.n1790 0.00139286
R59513 VCC.n1913 VCC.n1828 0.00139286
R59514 VCC.n2011 VCC.n1765 0.00139286
R59515 VCC.n2066 VCC.n1751 0.00139286
R59516 VCC.n2193 VCC.n1680 0.00139286
R59517 VCC.n2206 VCC.n1671 0.00139286
R59518 VCC.n2756 VCC.n2755 0.00139286
R59519 VCC.n2234 VCC.n2231 0.00139286
R59520 VCC.n2568 VCC.n2322 0.00139286
R59521 VCC.n2623 VCC.n2308 0.00139286
R59522 VCC.n2433 VCC.n2412 0.00139286
R59523 VCC.n2456 VCC.n2455 0.00139286
R59524 VCC.n2473 VCC.n2472 0.00139286
R59525 VCC.n2513 VCC.n2348 0.00139286
R59526 VCC.n2471 VCC.n2386 0.00139286
R59527 VCC.n2984 VCC.n2963 0.00139286
R59528 VCC.n3007 VCC.n3006 0.00139286
R59529 VCC.n3024 VCC.n3023 0.00139286
R59530 VCC.n3064 VCC.n2899 0.00139286
R59531 VCC.n3022 VCC.n2937 0.00139286
R59532 VCC.n3120 VCC.n2874 0.00139286
R59533 VCC.n3175 VCC.n2860 0.00139286
R59534 VCC.n3302 VCC.n2789 0.00139286
R59535 VCC.n3315 VCC.n2780 0.00139286
R59536 VCC.n3865 VCC.n3864 0.00139286
R59537 VCC.n3343 VCC.n3340 0.00139286
R59538 VCC.n3677 VCC.n3431 0.00139286
R59539 VCC.n3732 VCC.n3417 0.00139286
R59540 VCC.n3542 VCC.n3521 0.00139286
R59541 VCC.n3565 VCC.n3564 0.00139286
R59542 VCC.n3582 VCC.n3581 0.00139286
R59543 VCC.n3622 VCC.n3457 0.00139286
R59544 VCC.n3580 VCC.n3495 0.00139286
R59545 VCC.n4093 VCC.n4072 0.00139286
R59546 VCC.n4116 VCC.n4115 0.00139286
R59547 VCC.n4133 VCC.n4132 0.00139286
R59548 VCC.n4173 VCC.n4008 0.00139286
R59549 VCC.n4131 VCC.n4046 0.00139286
R59550 VCC.n4229 VCC.n3983 0.00139286
R59551 VCC.n4284 VCC.n3969 0.00139286
R59552 VCC.n4411 VCC.n3898 0.00139286
R59553 VCC.n4424 VCC.n3889 0.00139286
R59554 VCC.n4974 VCC.n4973 0.00139286
R59555 VCC.n4452 VCC.n4449 0.00139286
R59556 VCC.n4786 VCC.n4540 0.00139286
R59557 VCC.n4841 VCC.n4526 0.00139286
R59558 VCC.n4651 VCC.n4630 0.00139286
R59559 VCC.n4674 VCC.n4673 0.00139286
R59560 VCC.n4691 VCC.n4690 0.00139286
R59561 VCC.n4731 VCC.n4566 0.00139286
R59562 VCC.n4689 VCC.n4604 0.00139286
R59563 VCC.n5202 VCC.n5181 0.00139286
R59564 VCC.n5225 VCC.n5224 0.00139286
R59565 VCC.n5242 VCC.n5241 0.00139286
R59566 VCC.n5282 VCC.n5117 0.00139286
R59567 VCC.n5240 VCC.n5155 0.00139286
R59568 VCC.n5338 VCC.n5092 0.00139286
R59569 VCC.n5393 VCC.n5078 0.00139286
R59570 VCC.n5520 VCC.n5007 0.00139286
R59571 VCC.n5533 VCC.n4998 0.00139286
R59572 VCC.n6083 VCC.n6082 0.00139286
R59573 VCC.n5561 VCC.n5558 0.00139286
R59574 VCC.n5895 VCC.n5649 0.00139286
R59575 VCC.n5950 VCC.n5635 0.00139286
R59576 VCC.n5760 VCC.n5739 0.00139286
R59577 VCC.n5783 VCC.n5782 0.00139286
R59578 VCC.n5800 VCC.n5799 0.00139286
R59579 VCC.n5840 VCC.n5675 0.00139286
R59580 VCC.n5798 VCC.n5713 0.00139286
R59581 VCC.n6311 VCC.n6290 0.00139286
R59582 VCC.n6334 VCC.n6333 0.00139286
R59583 VCC.n6351 VCC.n6350 0.00139286
R59584 VCC.n6391 VCC.n6226 0.00139286
R59585 VCC.n6349 VCC.n6264 0.00139286
R59586 VCC.n6447 VCC.n6201 0.00139286
R59587 VCC.n6502 VCC.n6187 0.00139286
R59588 VCC.n6629 VCC.n6116 0.00139286
R59589 VCC.n6642 VCC.n6107 0.00139286
R59590 VCC.n7192 VCC.n7191 0.00139286
R59591 VCC.n6670 VCC.n6667 0.00139286
R59592 VCC.n7004 VCC.n6758 0.00139286
R59593 VCC.n7059 VCC.n6744 0.00139286
R59594 VCC.n6869 VCC.n6848 0.00139286
R59595 VCC.n6892 VCC.n6891 0.00139286
R59596 VCC.n6909 VCC.n6908 0.00139286
R59597 VCC.n6949 VCC.n6784 0.00139286
R59598 VCC.n6907 VCC.n6822 0.00139286
R59599 VCC.n7420 VCC.n7399 0.00139286
R59600 VCC.n7443 VCC.n7442 0.00139286
R59601 VCC.n7460 VCC.n7459 0.00139286
R59602 VCC.n7500 VCC.n7335 0.00139286
R59603 VCC.n7458 VCC.n7373 0.00139286
R59604 VCC.n7556 VCC.n7310 0.00139286
R59605 VCC.n7611 VCC.n7296 0.00139286
R59606 VCC.n7738 VCC.n7225 0.00139286
R59607 VCC.n7751 VCC.n7216 0.00139286
R59608 VCC.n8301 VCC.n8300 0.00139286
R59609 VCC.n7779 VCC.n7776 0.00139286
R59610 VCC.n8113 VCC.n7867 0.00139286
R59611 VCC.n8168 VCC.n7853 0.00139286
R59612 VCC.n7978 VCC.n7957 0.00139286
R59613 VCC.n8001 VCC.n8000 0.00139286
R59614 VCC.n8018 VCC.n8017 0.00139286
R59615 VCC.n8058 VCC.n7893 0.00139286
R59616 VCC.n8016 VCC.n7931 0.00139286
R59617 VCC.n8665 VCC.n8419 0.00139286
R59618 VCC.n8720 VCC.n8405 0.00139286
R59619 VCC.n8847 VCC.n8334 0.00139286
R59620 VCC.n8860 VCC.n8325 0.00139286
R59621 VCC.n8529 VCC.n8508 0.00139286
R59622 VCC.n8552 VCC.n8551 0.00139286
R59623 VCC.n8569 VCC.n8568 0.00139286
R59624 VCC.n8609 VCC.n8444 0.00139286
R59625 VCC.n8567 VCC.n8482 0.00139286
R59626 VCC.n9410 VCC.n9409 0.00139286
R59627 VCC.n8888 VCC.n8885 0.00139286
R59628 VCC.n9222 VCC.n8976 0.00139286
R59629 VCC.n9277 VCC.n8962 0.00139286
R59630 VCC.n9087 VCC.n9066 0.00139286
R59631 VCC.n9110 VCC.n9109 0.00139286
R59632 VCC.n9127 VCC.n9126 0.00139286
R59633 VCC.n9167 VCC.n9002 0.00139286
R59634 VCC.n9125 VCC.n9040 0.00139286
R59635 VCC.n9638 VCC.n9617 0.00139286
R59636 VCC.n9661 VCC.n9660 0.00139286
R59637 VCC.n9678 VCC.n9677 0.00139286
R59638 VCC.n9718 VCC.n9553 0.00139286
R59639 VCC.n9676 VCC.n9591 0.00139286
R59640 VCC.n9774 VCC.n9528 0.00139286
R59641 VCC.n9829 VCC.n9514 0.00139286
R59642 VCC.n9956 VCC.n9443 0.00139286
R59643 VCC.n9969 VCC.n9434 0.00139286
R59644 VCC.n10518 VCC.n10517 0.00139286
R59645 VCC.n9996 VCC.n9993 0.00139286
R59646 VCC.n10330 VCC.n10084 0.00139286
R59647 VCC.n10385 VCC.n10070 0.00139286
R59648 VCC.n10195 VCC.n10174 0.00139286
R59649 VCC.n10218 VCC.n10217 0.00139286
R59650 VCC.n10235 VCC.n10234 0.00139286
R59651 VCC.n10275 VCC.n10110 0.00139286
R59652 VCC.n10233 VCC.n10148 0.00139286
R59653 VCC.n10745 VCC.n10724 0.00139286
R59654 VCC.n10768 VCC.n10767 0.00139286
R59655 VCC.n10785 VCC.n10784 0.00139286
R59656 VCC.n10825 VCC.n10660 0.00139286
R59657 VCC.n10783 VCC.n10698 0.00139286
R59658 VCC.n10881 VCC.n10635 0.00139286
R59659 VCC.n10936 VCC.n10621 0.00139286
R59660 VCC.n11063 VCC.n10550 0.00139286
R59661 VCC.n11076 VCC.n10541 0.00139286
R59662 VCC.n11625 VCC.n11624 0.00139286
R59663 VCC.n11103 VCC.n11100 0.00139286
R59664 VCC.n11437 VCC.n11191 0.00139286
R59665 VCC.n11492 VCC.n11177 0.00139286
R59666 VCC.n11302 VCC.n11281 0.00139286
R59667 VCC.n11325 VCC.n11324 0.00139286
R59668 VCC.n11342 VCC.n11341 0.00139286
R59669 VCC.n11382 VCC.n11217 0.00139286
R59670 VCC.n11340 VCC.n11255 0.00139286
R59671 VCC.n11852 VCC.n11831 0.00139286
R59672 VCC.n11875 VCC.n11874 0.00139286
R59673 VCC.n11892 VCC.n11891 0.00139286
R59674 VCC.n11932 VCC.n11767 0.00139286
R59675 VCC.n11890 VCC.n11805 0.00139286
R59676 VCC.n11988 VCC.n11742 0.00139286
R59677 VCC.n12043 VCC.n11728 0.00139286
R59678 VCC.n12170 VCC.n11657 0.00139286
R59679 VCC.n12183 VCC.n11648 0.00139286
R59680 VCC.n12732 VCC.n12731 0.00139286
R59681 VCC.n12210 VCC.n12207 0.00139286
R59682 VCC.n12544 VCC.n12298 0.00139286
R59683 VCC.n12599 VCC.n12284 0.00139286
R59684 VCC.n12409 VCC.n12388 0.00139286
R59685 VCC.n12432 VCC.n12431 0.00139286
R59686 VCC.n12449 VCC.n12448 0.00139286
R59687 VCC.n12489 VCC.n12324 0.00139286
R59688 VCC.n12447 VCC.n12362 0.00139286
R59689 VCC.n12959 VCC.n12938 0.00139286
R59690 VCC.n12982 VCC.n12981 0.00139286
R59691 VCC.n12999 VCC.n12998 0.00139286
R59692 VCC.n13039 VCC.n12874 0.00139286
R59693 VCC.n12997 VCC.n12912 0.00139286
R59694 VCC.n13095 VCC.n12849 0.00139286
R59695 VCC.n13150 VCC.n12835 0.00139286
R59696 VCC.n13277 VCC.n12764 0.00139286
R59697 VCC.n13290 VCC.n12755 0.00139286
R59698 VCC.n13839 VCC.n13838 0.00139286
R59699 VCC.n13317 VCC.n13314 0.00139286
R59700 VCC.n13651 VCC.n13405 0.00139286
R59701 VCC.n13706 VCC.n13391 0.00139286
R59702 VCC.n13516 VCC.n13495 0.00139286
R59703 VCC.n13539 VCC.n13538 0.00139286
R59704 VCC.n13556 VCC.n13555 0.00139286
R59705 VCC.n13596 VCC.n13431 0.00139286
R59706 VCC.n13554 VCC.n13469 0.00139286
R59707 VCC.n14066 VCC.n14045 0.00139286
R59708 VCC.n14089 VCC.n14088 0.00139286
R59709 VCC.n14106 VCC.n14105 0.00139286
R59710 VCC.n14146 VCC.n13981 0.00139286
R59711 VCC.n14104 VCC.n14019 0.00139286
R59712 VCC.n14202 VCC.n13956 0.00139286
R59713 VCC.n14257 VCC.n13942 0.00139286
R59714 VCC.n14384 VCC.n13871 0.00139286
R59715 VCC.n14397 VCC.n13862 0.00139286
R59716 VCC.n14946 VCC.n14945 0.00139286
R59717 VCC.n14424 VCC.n14421 0.00139286
R59718 VCC.n14758 VCC.n14512 0.00139286
R59719 VCC.n14813 VCC.n14498 0.00139286
R59720 VCC.n14623 VCC.n14602 0.00139286
R59721 VCC.n14646 VCC.n14645 0.00139286
R59722 VCC.n14663 VCC.n14662 0.00139286
R59723 VCC.n14703 VCC.n14538 0.00139286
R59724 VCC.n14661 VCC.n14576 0.00139286
R59725 VCC.n15173 VCC.n15152 0.00139286
R59726 VCC.n15196 VCC.n15195 0.00139286
R59727 VCC.n15213 VCC.n15212 0.00139286
R59728 VCC.n15253 VCC.n15088 0.00139286
R59729 VCC.n15211 VCC.n15126 0.00139286
R59730 VCC.n15309 VCC.n15063 0.00139286
R59731 VCC.n15364 VCC.n15049 0.00139286
R59732 VCC.n15491 VCC.n14978 0.00139286
R59733 VCC.n15504 VCC.n14969 0.00139286
R59734 VCC.n16053 VCC.n16052 0.00139286
R59735 VCC.n15531 VCC.n15528 0.00139286
R59736 VCC.n15865 VCC.n15619 0.00139286
R59737 VCC.n15920 VCC.n15605 0.00139286
R59738 VCC.n15730 VCC.n15709 0.00139286
R59739 VCC.n15753 VCC.n15752 0.00139286
R59740 VCC.n15770 VCC.n15769 0.00139286
R59741 VCC.n15810 VCC.n15645 0.00139286
R59742 VCC.n15768 VCC.n15683 0.00139286
R59743 VCC.n16280 VCC.n16259 0.00139286
R59744 VCC.n16303 VCC.n16302 0.00139286
R59745 VCC.n16320 VCC.n16319 0.00139286
R59746 VCC.n16360 VCC.n16195 0.00139286
R59747 VCC.n16318 VCC.n16233 0.00139286
R59748 VCC.n16416 VCC.n16170 0.00139286
R59749 VCC.n16471 VCC.n16156 0.00139286
R59750 VCC.n16598 VCC.n16085 0.00139286
R59751 VCC.n16611 VCC.n16076 0.00139286
R59752 VCC.n17160 VCC.n17159 0.00139286
R59753 VCC.n16638 VCC.n16635 0.00139286
R59754 VCC.n16972 VCC.n16726 0.00139286
R59755 VCC.n17027 VCC.n16712 0.00139286
R59756 VCC.n16837 VCC.n16816 0.00139286
R59757 VCC.n16860 VCC.n16859 0.00139286
R59758 VCC.n16877 VCC.n16876 0.00139286
R59759 VCC.n16917 VCC.n16752 0.00139286
R59760 VCC.n16875 VCC.n16790 0.00139286
R59761 VCC.n17336 VCC.n17277 0.00139286
R59762 VCC.n17391 VCC.n17263 0.00139286
R59763 VCC.n17518 VCC.n17192 0.00139286
R59764 VCC.n17531 VCC.n17183 0.00139286
R59765 VCC.n17541 VCC.n17174 0.00054824
R59766 VCC.n17543 VCC.n16067 0.00054824
R59767 VCC.n17545 VCC.n14960 0.00054824
R59768 VCC.n17547 VCC.n13853 0.00054824
R59769 VCC.n17549 VCC.n12746 0.00054824
R59770 VCC.n17551 VCC.n11639 0.00054824
R59771 VCC.n17553 VCC.n10532 0.00054824
R59772 VCC.n9425 VCC.n9424 0.00054824
R59773 VCC.n8316 VCC.n8315 0.00054824
R59774 VCC.n7207 VCC.n7206 0.00054824
R59775 VCC.n6098 VCC.n6097 0.00054824
R59776 VCC.n4989 VCC.n4988 0.00054824
R59777 VCC.n3880 VCC.n3879 0.00054824
R59778 VCC.n2771 VCC.n2770 0.00054824
R59779 VCC.n1662 VCC.n1661 0.00054824
R59780 6_bit_dac_0[1].5_bit_dac_1.D3.n0 6_bit_dac_0[1].5_bit_dac_1.D3.n1 173.293
R59781 6_bit_dac_0[1].5_bit_dac_1.D3 6_bit_dac_0[1].5_bit_dac_1.D3.n2 125.046
R59782 6_bit_dac_0[1].5_bit_dac_1.D3.n1 6_bit_dac_0[1].5_bit_dac_1.D3.t4 84.3505
R59783 6_bit_dac_0[1].5_bit_dac_1.D3.n2 6_bit_dac_0[1].5_bit_dac_1.D3.t3 77.1205
R59784 6_bit_dac_0[1].5_bit_dac_1.D3.n2 6_bit_dac_0[1].5_bit_dac_1.D3.t2 61.6965
R59785 6_bit_dac_0[1].5_bit_dac_1.D3.n1 6_bit_dac_0[1].5_bit_dac_1.D3.t5 53.5025
R59786 6_bit_dac_0[1].5_bit_dac_1.D3.n0 6_bit_dac_0[1].5_bit_dac_1.D3.t0 46.9077
R59787 6_bit_dac_0[1].5_bit_dac_1.D3.n0 6_bit_dac_0[1].5_bit_dac_1.D3.t1 35.0239
R59788 6_bit_dac_0[1].5_bit_dac_1.D3 6_bit_dac_0[1].5_bit_dac_1.D3.n0 3.95473
R59789 6_bit_dac_0[1].5_bit_dac_1.D4.n0 6_bit_dac_0[1].5_bit_dac_1.D4.n1 173.293
R59790 6_bit_dac_0[1].5_bit_dac_1.D4 6_bit_dac_0[1].5_bit_dac_1.D4.n2 125.046
R59791 6_bit_dac_0[1].5_bit_dac_1.D4.n1 6_bit_dac_0[1].5_bit_dac_1.D4.t5 84.3505
R59792 6_bit_dac_0[1].5_bit_dac_1.D4.n2 6_bit_dac_0[1].5_bit_dac_1.D4.t2 77.1205
R59793 6_bit_dac_0[1].5_bit_dac_1.D4.n2 6_bit_dac_0[1].5_bit_dac_1.D4.t4 61.6965
R59794 6_bit_dac_0[1].5_bit_dac_1.D4.n1 6_bit_dac_0[1].5_bit_dac_1.D4.t3 53.5025
R59795 6_bit_dac_0[1].5_bit_dac_1.D4.n0 6_bit_dac_0[1].5_bit_dac_1.D4.t0 46.9077
R59796 6_bit_dac_0[1].5_bit_dac_1.D4.n0 6_bit_dac_0[1].5_bit_dac_1.D4.t1 35.0239
R59797 6_bit_dac_0[1].5_bit_dac_1.D4 6_bit_dac_0[1].5_bit_dac_1.D4.n0 3.95498
R59798 6_bit_dac_0[0].5_bit_dac_0.VOUT.n1 6_bit_dac_0[0].5_bit_dac_0.VOUT.t5 49.5021
R59799 6_bit_dac_0[0].5_bit_dac_0.VOUT.n2 6_bit_dac_0[0].5_bit_dac_0.VOUT.t1 46.8495
R59800 6_bit_dac_0[0].5_bit_dac_0.VOUT.n2 6_bit_dac_0[0].5_bit_dac_0.VOUT.t4 46.5654
R59801 6_bit_dac_0[0].5_bit_dac_0.VOUT.n1 6_bit_dac_0[0].5_bit_dac_0.VOUT.t3 40.9453
R59802 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 6_bit_dac_0[0].5_bit_dac_0.VOUT.t0 34.8869
R59803 6_bit_dac_0[0].5_bit_dac_0.VOUT.n8 6_bit_dac_0[0].5_bit_dac_0.VOUT.t2 27.6955
R59804 6_bit_dac_0[0].5_bit_dac_0.VOUT.n5 6_bit_dac_0[0].5_bit_dac_0.VOUT.n4 13.362
R59805 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 6_bit_dac_0[0].5_bit_dac_0.VOUT.n6 9.3005
R59806 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 6_bit_dac_0[0].5_bit_dac_0.VOUT.n3 9.3005
R59807 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 6_bit_dac_0[0].5_bit_dac_0.VOUT.n7 9.3005
R59808 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 6_bit_dac_0[0].5_bit_dac_0.VOUT.n9 9.3005
R59809 6_bit_dac_0[0].5_bit_dac_0.VOUT.n9 6_bit_dac_0[0].5_bit_dac_0.VOUT.n8 9.02061
R59810 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 6_bit_dac_0[0].5_bit_dac_0.VOUT.n5 4.55875
R59811 6_bit_dac_0[0].5_bit_dac_0.VOUT.n2 6_bit_dac_0[0].5_bit_dac_0.VOUT 2.96822
R59812 6_bit_dac_0[0].5_bit_dac_0.VOUT 6_bit_dac_0[0].5_bit_dac_0.VOUT.n1 1.26728
R59813 6_bit_dac_0[0].5_bit_dac_0.VOUT 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 0.815717
R59814 6_bit_dac_0[0].5_bit_dac_0.VOUT.n0 6_bit_dac_0[0].5_bit_dac_0.VOUT.n2 0.716261
R59815 switch_n_3v3_1.D5.n0 switch_n_3v3_1.D5.n1 173.293
R59816 switch_n_3v3_1.D5 switch_n_3v3_1.D5.n2 125.046
R59817 switch_n_3v3_1.D5.n1 switch_n_3v3_1.D5.t2 84.3505
R59818 switch_n_3v3_1.D5.n2 switch_n_3v3_1.D5.t5 77.1205
R59819 switch_n_3v3_1.D5.n2 switch_n_3v3_1.D5.t4 61.6965
R59820 switch_n_3v3_1.D5.n1 switch_n_3v3_1.D5.t3 53.5025
R59821 switch_n_3v3_1.D5.n0 switch_n_3v3_1.D5.t0 46.9077
R59822 switch_n_3v3_1.D5.n0 switch_n_3v3_1.D5.t1 35.0239
R59823 switch_n_3v3_1.D5 switch_n_3v3_1.D5.n0 3.95338
R59824 D1.n1 D1.n0 127.099
R59825 D1.n0 D1.t0 77.6025
R59826 D1.n0 D1.t1 61.2145
R59827 D1.n1 D1 0.0485769
R59828 D1 D1.n1 0.0365577
R59829 D3 D3.n0 125.046
R59830 D3.n0 D3.t0 77.1205
R59831 D3.n0 D3.t1 61.6965
R59832 D5 D5.n0 125.046
R59833 D5.n0 D5.t0 77.1205
R59834 D5.n0 D5.t1 61.6965
R59835 VREFL.n1 VREFL.t2 99.7169
R59836 VREFL.n0 VREFL.t1 44.9543
R59837 VREFL.n0 VREFL.t0 37.5373
R59838 VREFL.n1 VREFL.n0 2.88557
R59839 VREFL VREFL.n1 1.84958
R59840 D6_BUF.n2 D6_BUF.n1 173.293
R59841 D6_BUF.n1 D6_BUF.t2 84.3505
R59842 D6_BUF.n1 D6_BUF.t3 53.5025
R59843 D6_BUF.n0 D6_BUF.t0 46.9077
R59844 D6_BUF.n0 D6_BUF.t1 35.0239
R59845 D6_BUF D6_BUF.n2 3.75226
R59846 D6_BUF.n2 D6_BUF.n0 0.204238
R59847 6_bit_dac_0[1].VOUT.n1 6_bit_dac_0[1].VOUT.n0 0.0523282
R59848 6_bit_dac_0[1].VOUT.n3 6_bit_dac_0[1].VOUT.t0 49.5021
R59849 6_bit_dac_0[1].VOUT.n2 6_bit_dac_0[1].VOUT.t2 46.8495
R59850 6_bit_dac_0[1].VOUT.n2 6_bit_dac_0[1].VOUT.t5 46.5654
R59851 6_bit_dac_0[1].VOUT.n3 6_bit_dac_0[1].VOUT.t1 40.9445
R59852 6_bit_dac_0[1].VOUT.n1 6_bit_dac_0[1].VOUT.t3 34.887
R59853 6_bit_dac_0[1].VOUT.n0 6_bit_dac_0[1].VOUT.t4 34.5611
R59854 6_bit_dac_0[1].VOUT.n2 6_bit_dac_0[1].VOUT 3.09322
R59855 6_bit_dac_0[1].VOUT 6_bit_dac_0[1].VOUT.n3 1.26445
R59856 6_bit_dac_0[1].VOUT 6_bit_dac_0[1].VOUT.n0 0.867541
R59857 6_bit_dac_0[1].VOUT.n1 6_bit_dac_0[1].VOUT.n2 0.613
R59858 VOUT.n0 VOUT.t0 46.8495
R59859 VOUT.n0 VOUT.t3 46.5654
R59860 VOUT.n5 VOUT.t1 34.887
R59861 VOUT.n10 VOUT.t2 27.6955
R59862 VOUT.n4 VOUT.n3 13.362
R59863 VOUT.n2 VOUT.n1 9.3005
R59864 VOUT.n7 VOUT.n6 9.3005
R59865 VOUT.n9 VOUT.n8 9.3005
R59866 VOUT.n12 VOUT.n11 9.3005
R59867 VOUT.n11 VOUT.n10 9.02061
R59868 VOUT.n5 VOUT.n4 4.55875
R59869 VOUT.n0 VOUT 3.09322
R59870 VOUT VOUT.n12 0.815717
R59871 VOUT.n2 VOUT.n0 0.613
R59872 VOUT.n12 VOUT.n9 0.0439783
R59873 VOUT.n7 VOUT.n5 0.0439783
R59874 VOUT.n5 VOUT.n2 0.014087
R59875 VOUT.n9 VOUT.n7 0.00321739
R59876 D2_BUF.n2 D2_BUF.n1 173.293
R59877 D2_BUF.n1 D2_BUF.t3 84.3505
R59878 D2_BUF.n1 D2_BUF.t2 53.5025
R59879 D2_BUF.n0 D2_BUF.t0 46.9077
R59880 D2_BUF.n0 D2_BUF.t1 35.0239
R59881 D2_BUF D2_BUF.n2 3.75226
R59882 D2_BUF.n2 D2_BUF.n0 0.204238
R59883 6_bit_dac_0[0].5_bit_dac_1.D4.n0 6_bit_dac_0[0].5_bit_dac_1.D4.n1 173.293
R59884 6_bit_dac_0[0].5_bit_dac_1.D4 6_bit_dac_0[0].5_bit_dac_1.D4.n2 125.046
R59885 6_bit_dac_0[0].5_bit_dac_1.D4.n1 6_bit_dac_0[0].5_bit_dac_1.D4.t5 84.3505
R59886 6_bit_dac_0[0].5_bit_dac_1.D4.n2 6_bit_dac_0[0].5_bit_dac_1.D4.t4 77.1205
R59887 6_bit_dac_0[0].5_bit_dac_1.D4.n2 6_bit_dac_0[0].5_bit_dac_1.D4.t3 61.6965
R59888 6_bit_dac_0[0].5_bit_dac_1.D4.n1 6_bit_dac_0[0].5_bit_dac_1.D4.t2 53.5025
R59889 6_bit_dac_0[0].5_bit_dac_1.D4.n0 6_bit_dac_0[0].5_bit_dac_1.D4.t0 46.9077
R59890 6_bit_dac_0[0].5_bit_dac_1.D4.n0 6_bit_dac_0[0].5_bit_dac_1.D4.t1 35.0239
R59891 6_bit_dac_0[0].5_bit_dac_1.D4 6_bit_dac_0[0].5_bit_dac_1.D4.n0 3.95498
R59892 D5_BUF.n2 D5_BUF.n1 173.293
R59893 D5_BUF.n1 D5_BUF.t2 84.3505
R59894 D5_BUF.n1 D5_BUF.t3 53.5025
R59895 D5_BUF.n0 D5_BUF.t0 46.9077
R59896 D5_BUF.n0 D5_BUF.t1 35.0239
R59897 D5_BUF D5_BUF.n2 3.74964
R59898 D5_BUF.n2 D5_BUF.n0 0.204238
R59899 6_bit_dac_0[0].VOUT.n0 6_bit_dac_0[0].VOUT.n1 0.0523299
R59900 6_bit_dac_0[0].VOUT 6_bit_dac_0[0].VOUT.t3 49.82
R59901 6_bit_dac_0[0].VOUT.n2 6_bit_dac_0[0].VOUT.t4 46.8495
R59902 6_bit_dac_0[0].VOUT.n2 6_bit_dac_0[0].VOUT.t2 46.5654
R59903 6_bit_dac_0[0].VOUT 6_bit_dac_0[0].VOUT.t0 36.7243
R59904 6_bit_dac_0[0].VOUT.n1 6_bit_dac_0[0].VOUT.t5 34.887
R59905 6_bit_dac_0[0].VOUT.t1 6_bit_dac_0[0].VOUT.n0 34.5609
R59906 6_bit_dac_0[0].VOUT.n2 6_bit_dac_0[0].VOUT 3.09322
R59907 6_bit_dac_0[0].VOUT 6_bit_dac_0[0].VOUT.n0 0.86754
R59908 6_bit_dac_0[0].VOUT.n1 6_bit_dac_0[0].VOUT.n2 0.613
R59909 6_bit_dac_0[0].5_bit_dac_1.D3.n0 6_bit_dac_0[0].5_bit_dac_1.D3.n1 173.293
R59910 6_bit_dac_0[0].5_bit_dac_1.D3 6_bit_dac_0[0].5_bit_dac_1.D3.n2 125.046
R59911 6_bit_dac_0[0].5_bit_dac_1.D3.n1 6_bit_dac_0[0].5_bit_dac_1.D3.t3 84.3505
R59912 6_bit_dac_0[0].5_bit_dac_1.D3.n2 6_bit_dac_0[0].5_bit_dac_1.D3.t2 77.1205
R59913 6_bit_dac_0[0].5_bit_dac_1.D3.n2 6_bit_dac_0[0].5_bit_dac_1.D3.t5 61.6965
R59914 6_bit_dac_0[0].5_bit_dac_1.D3.n1 6_bit_dac_0[0].5_bit_dac_1.D3.t4 53.5025
R59915 6_bit_dac_0[0].5_bit_dac_1.D3.n0 6_bit_dac_0[0].5_bit_dac_1.D3.t0 46.9077
R59916 6_bit_dac_0[0].5_bit_dac_1.D3.n0 6_bit_dac_0[0].5_bit_dac_1.D3.t1 35.0239
R59917 6_bit_dac_0[0].5_bit_dac_1.D3 6_bit_dac_0[0].5_bit_dac_1.D3.n0 3.95473
R59918 D4_BUF.n2 D4_BUF.n1 173.293
R59919 D4_BUF.n1 D4_BUF.t3 84.3505
R59920 D4_BUF.n1 D4_BUF.t2 53.5025
R59921 D4_BUF.n0 D4_BUF.t0 46.9077
R59922 D4_BUF.n0 D4_BUF.t1 35.0239
R59923 D4_BUF D4_BUF.n2 3.75124
R59924 D4_BUF.n2 D4_BUF.n0 0.204238
R59925 D3_BUF.n2 D3_BUF.n1 173.293
R59926 D3_BUF.n1 D3_BUF.t2 84.3505
R59927 D3_BUF.n1 D3_BUF.t3 53.5025
R59928 D3_BUF.n0 D3_BUF.t0 46.9077
R59929 D3_BUF.n0 D3_BUF.t1 35.0239
R59930 D3_BUF D3_BUF.n2 3.75099
R59931 D3_BUF.n2 D3_BUF.n0 0.204238
R59932 switch_n_3v3_1.D3.n0 switch_n_3v3_1.D3.n1 173.293
R59933 switch_n_3v3_1.D3 switch_n_3v3_1.D3.n2 125.046
R59934 switch_n_3v3_1.D3.n1 switch_n_3v3_1.D3.t5 84.3505
R59935 switch_n_3v3_1.D3.n2 switch_n_3v3_1.D3.t4 77.1205
R59936 switch_n_3v3_1.D3.n2 switch_n_3v3_1.D3.t2 61.6965
R59937 switch_n_3v3_1.D3.n1 switch_n_3v3_1.D3.t3 53.5025
R59938 switch_n_3v3_1.D3.n0 switch_n_3v3_1.D3.t0 46.9077
R59939 switch_n_3v3_1.D3.n0 switch_n_3v3_1.D3.t1 35.0239
R59940 switch_n_3v3_1.D3 switch_n_3v3_1.D3.n0 3.95473
R59941 switch_n_3v3_1.D4.n0 switch_n_3v3_1.D4.n1 173.293
R59942 switch_n_3v3_1.D4 switch_n_3v3_1.D4.n2 125.046
R59943 switch_n_3v3_1.D4.n1 switch_n_3v3_1.D4.t3 84.3505
R59944 switch_n_3v3_1.D4.n2 switch_n_3v3_1.D4.t5 77.1205
R59945 switch_n_3v3_1.D4.n2 switch_n_3v3_1.D4.t2 61.6965
R59946 switch_n_3v3_1.D4.n1 switch_n_3v3_1.D4.t4 53.5025
R59947 switch_n_3v3_1.D4.n0 switch_n_3v3_1.D4.t0 46.9077
R59948 switch_n_3v3_1.D4.n0 switch_n_3v3_1.D4.t1 35.0239
R59949 switch_n_3v3_1.D4 switch_n_3v3_1.D4.n0 3.95498
R59950 6_bit_dac_0[1].5_bit_dac_1.VOUT 6_bit_dac_0[1].5_bit_dac_1.VOUT.t5 49.82
R59951 6_bit_dac_0[1].5_bit_dac_1.VOUT.n8 6_bit_dac_0[1].5_bit_dac_1.VOUT.t3 46.8495
R59952 6_bit_dac_0[1].5_bit_dac_1.VOUT.n8 6_bit_dac_0[1].5_bit_dac_1.VOUT.t0 46.5654
R59953 6_bit_dac_0[1].5_bit_dac_1.VOUT 6_bit_dac_0[1].5_bit_dac_1.VOUT.t4 36.7243
R59954 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 6_bit_dac_0[1].5_bit_dac_1.VOUT.t2 34.887
R59955 6_bit_dac_0[1].5_bit_dac_1.VOUT.n6 6_bit_dac_0[1].5_bit_dac_1.VOUT.t1 27.6955
R59956 6_bit_dac_0[1].5_bit_dac_1.VOUT.n5 6_bit_dac_0[1].5_bit_dac_1.VOUT.n4 13.362
R59957 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 6_bit_dac_0[1].5_bit_dac_1.VOUT.n3 9.3005
R59958 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 6_bit_dac_0[1].5_bit_dac_1.VOUT.n2 9.3005
R59959 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 6_bit_dac_0[1].5_bit_dac_1.VOUT.n1 9.3005
R59960 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 6_bit_dac_0[1].5_bit_dac_1.VOUT.n7 9.3005
R59961 6_bit_dac_0[1].5_bit_dac_1.VOUT.n7 6_bit_dac_0[1].5_bit_dac_1.VOUT.n6 9.0206
R59962 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 6_bit_dac_0[1].5_bit_dac_1.VOUT.n5 4.55875
R59963 6_bit_dac_0[1].5_bit_dac_1.VOUT 6_bit_dac_0[1].5_bit_dac_1.VOUT.n8 2.96822
R59964 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 6_bit_dac_0[1].5_bit_dac_1.VOUT 0.815717
R59965 6_bit_dac_0[1].5_bit_dac_1.VOUT.n8 6_bit_dac_0[1].5_bit_dac_1.VOUT.n0 0.716261
R59966 D2 D2.n0 125.046
R59967 D2.n0 D2.t1 77.1205
R59968 D2.n0 D2.t0 61.6965
R59969 D4 D4.n0 125.046
R59970 D4.n0 D4.t1 77.1205
R59971 D4.n0 D4.t0 61.6965
R59972 D1_BUF.n2 D1_BUF.n1 169.566
R59973 D1_BUF.n1 D1_BUF.t2 84.8325
R59974 D1_BUF.n1 D1_BUF.t3 53.0205
R59975 D1_BUF.n0 D1_BUF.t0 46.9158
R59976 D1_BUF.n0 D1_BUF.t1 35.0302
R59977 D1_BUF.n3 D1_BUF.n2 3.65455
R59978 D1_BUF D1_BUF.n3 2.56683
R59979 D1_BUF.n2 D1_BUF.n0 0.199588
R59980 D1_BUF.n3 D1_BUF 0.0389615
R59981 VREFH.n0 VREFH.t0 96.9442
R59982 VREFH VREFH.n0 1.07866
R59983 VREFH.n0 VREFH 0.00100409
R59984 D6 D6.n0 125.046
R59985 D6.n0 D6.t1 77.1205
R59986 D6.n0 D6.t0 61.6965
R59987 D0 D0.n0 115.853
R59988 D0.n0 D0.t1 81.9405
R59989 D0.n0 D0.t0 56.8765
C0 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C1 a_544_22941# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C2 VCC 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C3 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C4 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 D4 1.25f
C5 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 1.29f
C6 VCC 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.18f
C7 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C8 VCC 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.18f
C9 VCC 6_bit_dac_0[1].5_bit_dac_1.D0 1.18f
C10 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.06f
C11 VCC 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 1.18f
C12 a_544_31537# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C13 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C14 VCC 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 1.18f
C15 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C16 a_544_19257# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C17 a_544_30309# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C18 a_544_13117# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C19 switch_n_3v3_1.D3 switch_n_3v3_1.D2 1.29f
C20 6_bit_dac_0[0].5_bit_dac_1.VREFL 6_bit_dac_0[0].5_bit_dac_1.D0 1.06f
C21 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.06f
C22 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C23 a_544_15573# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C24 VCC D6_BUF 1.16f
C25 switch_n_3v3_1.D5 D6 5.01f
C26 a_544_16801# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C27 switch_n_3v3_1.D5 switch_n_3v3_1.D4 5.04f
C28 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C29 VCC 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.18f
C30 D5_BUF D4_BUF 2.18f
C31 switch_n_3v3_1.D4 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 1.25f
C32 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C33 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C34 VCC 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C35 VCC 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 1.18f
C36 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C37 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 1.06f
C38 D6_BUF switch_n_3v3_1.D7 9.7f
C39 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 1.06f
C40 VCC 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C41 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C42 D3 D4 1.02f
C43 VCC switch_n_3v3_1.D7 4.34f
C44 a_544_37677# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C45 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.06f
C46 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C47 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C48 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 1.29f
C49 a_544_11889# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C50 VCC 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C51 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.06f
C52 VCC 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.18f
C53 a_544_10661# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C54 VCC 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.17f
C55 6_bit_dac_0[0].VOUT 6_bit_dac_0[0].5_bit_dac_0.VOUT 2.26f
C56 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 switch_n_3v3_1.D4 1.25f
C57 VCC 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.18f
C58 a_544_33993# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C59 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C60 VCC 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C61 a_544_5749# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C62 VCC 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C63 a_544_29081# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C64 VCC 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C65 VCC 6_bit_dac_0[1].VOUT 1.26f
C66 a_544_24169# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C67 a_544_21713# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C68 a_544_38905# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C69 VCC 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C70 6_bit_dac_0[1].5_bit_dac_1.VOUT 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT 1.52f
C71 VCC 6_bit_dac_0[0].D0 1.18f
C72 a_544_25397# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C73 VCC 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C74 VCC 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C75 a_544_35221# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C76 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 D4_BUF 1.25f
C77 VCC 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.18f
C78 a_544_837# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C79 a_544_26625# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C80 a_544_36449# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C81 switch_n_3v3_1.D5 D6_BUF 5.01f
C82 a_544_18029# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C83 VCC switch_n_3v3_1.D5 1.41f
C84 a_544_2065# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C85 6_bit_dac_0[0].5_bit_dac_1.VOUT 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT 1.52f
C86 VCC 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C87 VCC 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.18f
C88 a_544_14345# 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C89 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.06f
C90 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 1.29f
C91 a_544_9433# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C92 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 1.29f
C93 6_bit_dac_0[1].VREFH 6_bit_dac_0[0].D0 1.06f
C94 VCC 6_bit_dac_0[0].5_bit_dac_1.D0 1.18f
C95 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.06f
C96 VCC 6_bit_dac_0[0].VOUT 1.07f
C97 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.06f
C98 a_544_8205# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C99 VCC 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C100 D6_BUF D5_BUF 4.69f
C101 VCC 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 1.18f
C102 D5 D6 4.78f
C103 6_bit_dac_0[1].VOUT 6_bit_dac_0[1].5_bit_dac_1.VOUT 2.21f
C104 VCC D6 1.1f
C105 VCC 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 1.18f
C106 a_544_4521# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C107 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 1.06f
C108 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C109 D4 D5 2.27f
C110 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C111 a_544_3293# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C112 a_544_6977# 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C113 VCC 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C114 a_544_32765# 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C115 6_bit_dac_0[1].5_bit_dac_1.VREFL 6_bit_dac_0[1].5_bit_dac_1.D0 1.06f
C116 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 1.06f
C117 switch_n_3v3_1.D4 switch_n_3v3_1.D3 2.53f
C118 D6 switch_n_3v3_1.D7 9.8f
C119 VCC 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C120 a_544_20485# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C121 VCC 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C122 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VREFH 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 1.06f
C123 a_544_27853# 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C124 switch_n_3v3_1.D7 VSS 7f
C125 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.53f
C126 D1_BUF VSS 1.17f
C127 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.13f
C128 D0_BUF VSS 2.53f
C129 a_1556_406# VSS 1.22f
C130 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.32f
C131 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.08f
C132 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C133 D2_BUF VSS 1.14f
C134 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.14f
C135 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.63f
C136 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C137 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.26f
C138 a_1556_1634# VSS 1.16f
C139 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.5f
C140 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C141 D3_BUF VSS 1.17f
C142 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.09f
C143 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS 1.61f
C144 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C145 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS 3.25f
C146 a_1556_2862# VSS 1.16f
C147 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS 1.42f
C148 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C149 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS 1.87f
C150 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f
C151 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C152 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C153 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f
C154 a_1556_4090# VSS 1.16f
C155 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C156 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].VOUT VSS 1.46f
C157 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f
C158 D4_BUF VSS 2.68f
C159 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.DX_ VSS 1.08f
C160 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D1 VSS 1.61f
C161 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C162 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[0].D0 VSS 3.25f
C163 a_1556_5318# VSS 1.16f
C164 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS 1.42f
C165 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f
C166 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f
C167 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C168 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D2 VSS 1.86f
C169 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f
C170 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f
C171 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C172 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f
C173 a_1556_6546# VSS 1.16f
C174 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f
C175 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].VOUT VSS 1.24f
C176 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C177 6_bit_dac_0[0].5_bit_dac_1.switch_n_3v3_0.D3 VSS 1.89f
C178 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.08f
C179 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS 1.61f
C180 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C181 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS 3.25f
C182 a_1556_7774# VSS 1.16f
C183 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS 1.42f
C184 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 1.04f
C185 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C186 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS 1.86f
C187 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f
C188 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C189 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C190 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f
C191 a_1556_9002# VSS 1.16f
C192 6_bit_dac_0[0].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C193 6_bit_dac_0[0].5_bit_dac_1.VOUT VSS 2.63f
C194 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f
C195 D5_BUF VSS 8.89f
C196 6_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.09f
C197 6_bit_dac_0[0].5_bit_dac_1.D1 VSS 1.61f
C198 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C199 6_bit_dac_0[0].5_bit_dac_1.D0 VSS 3.25f
C200 a_1556_10230# VSS 1.16f
C201 6_bit_dac_0[0].5_bit_dac_1.VREFL VSS 1.42f
C202 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f
C203 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f
C204 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C205 6_bit_dac_0[0].5_bit_dac_1.D2 VSS 1.86f
C206 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f
C207 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f
C208 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C209 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f
C210 a_1556_11458# VSS 1.16f
C211 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f
C212 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C213 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.08f
C214 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS 1.61f
C215 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C216 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS 3.25f
C217 a_1556_12686# VSS 1.16f
C218 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS 1.42f
C219 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C220 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS 1.86f
C221 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f
C222 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C223 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C224 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f
C225 a_1556_13914# VSS 1.16f
C226 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C227 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].VOUT VSS 1.22f
C228 6_bit_dac_0[0].5_bit_dac_0.VOUT VSS 2.75f
C229 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f
C230 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.DX_ VSS 1.08f
C231 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D1 VSS 1.61f
C232 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C233 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[0].D0 VSS 3.25f
C234 a_1556_15142# VSS 1.16f
C235 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS 1.42f
C236 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f
C237 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f
C238 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C239 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D2 VSS 1.86f
C240 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f
C241 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f
C242 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C243 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f
C244 a_1556_16370# VSS 1.16f
C245 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f
C246 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].VOUT VSS 1.32f
C247 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C248 6_bit_dac_0[0].5_bit_dac_0.switch_n_3v3_0.D3 VSS 1.89f
C249 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.08f
C250 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS 1.61f
C251 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C252 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS 3.25f
C253 a_1556_17598# VSS 1.16f
C254 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS 1.42f
C255 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 1.05f
C256 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C257 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS 1.86f
C258 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f
C259 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C260 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C261 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f
C262 a_1556_18826# VSS 1.16f
C263 6_bit_dac_0[0].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C264 6_bit_dac_0[0].VOUT VSS 5.69f
C265 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f
C266 D6_BUF VSS 19.3f
C267 switch_n_3v3_1.DX_ VSS 1.09f
C268 D6 VSS 20.5f
C269 6_bit_dac_0[0].D1 VSS 1.61f
C270 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C271 6_bit_dac_0[0].D0 VSS 3.25f
C272 a_1556_20054# VSS 1.16f
C273 6_bit_dac_0[1].VREFH VSS 1.42f
C274 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f
C275 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f
C276 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C277 switch_n_3v3_1.D2 VSS 1.86f
C278 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f
C279 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f
C280 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C281 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f
C282 a_1556_21282# VSS 1.16f
C283 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f
C284 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C285 switch_n_3v3_1.D3 VSS 3.39f
C286 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.08f
C287 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS 1.61f
C288 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C289 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS 3.25f
C290 a_1556_22510# VSS 1.16f
C291 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS 1.42f
C292 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C293 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS 1.86f
C294 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f
C295 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C296 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C297 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f
C298 a_1556_23738# VSS 1.16f
C299 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C300 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].VOUT VSS 1.25f
C301 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f
C302 switch_n_3v3_1.D4 VSS 7.7f
C303 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.DX_ VSS 1.08f
C304 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D1 VSS 1.61f
C305 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C306 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[0].D0 VSS 3.25f
C307 a_1556_24966# VSS 1.16f
C308 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VREFH VSS 1.42f
C309 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f
C310 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f
C311 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C312 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D2 VSS 1.86f
C313 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f
C314 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f
C315 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C316 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f
C317 a_1556_26194# VSS 1.16f
C318 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f
C319 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].VOUT VSS 1.24f
C320 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C321 6_bit_dac_0[1].5_bit_dac_1.switch_n_3v3_0.D3 VSS 1.89f
C322 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.08f
C323 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS 1.61f
C324 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C325 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS 3.25f
C326 a_1556_27422# VSS 1.16f
C327 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS 1.42f
C328 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 1.04f
C329 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C330 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS 1.86f
C331 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f
C332 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C333 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C334 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f
C335 a_1556_28650# VSS 1.16f
C336 6_bit_dac_0[1].5_bit_dac_1.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C337 6_bit_dac_0[1].5_bit_dac_1.VOUT VSS 3.31f
C338 6_bit_dac_0[1].VOUT VSS 5.53f
C339 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f
C340 switch_n_3v3_1.D5 VSS 19.7f
C341 6_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.08f
C342 D5 VSS 9.87f
C343 6_bit_dac_0[1].5_bit_dac_1.D1 VSS 1.61f
C344 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C345 6_bit_dac_0[1].5_bit_dac_1.D0 VSS 3.25f
C346 a_1556_29878# VSS 1.16f
C347 6_bit_dac_0[1].5_bit_dac_1.VREFL VSS 1.42f
C348 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f
C349 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f
C350 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C351 6_bit_dac_0[1].5_bit_dac_1.D2 VSS 1.86f
C352 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f
C353 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f
C354 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C355 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f
C356 a_1556_31106# VSS 1.16f
C357 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f
C358 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C359 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.08f
C360 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS 1.61f
C361 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C362 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS 3.25f
C363 a_1556_32334# VSS 1.16f
C364 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS 1.42f
C365 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C366 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].switch_n_3v3_0.D2 VSS 1.86f
C367 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f
C368 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C369 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C370 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f
C371 a_1556_33562# VSS 1.16f
C372 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C373 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].VOUT VSS 1.22f
C374 6_bit_dac_0[1].5_bit_dac_0.VOUT VSS 2.37f
C375 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f
C376 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.DX_ VSS 1.09f
C377 D4 VSS 2.71f
C378 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D1 VSS 1.61f
C379 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C380 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[0].D0 VSS 3.25f
C381 a_1556_34790# VSS 1.16f
C382 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VREFH VSS 1.42f
C383 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f
C384 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f
C385 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f
C386 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D2 VSS 1.86f
C387 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f
C388 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f
C389 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f
C390 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f
C391 a_1556_36018# VSS 1.16f
C392 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f
C393 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].VOUT VSS 1.73f
C394 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f
C395 6_bit_dac_0[1].5_bit_dac_0.switch_n_3v3_0.D3 VSS 1.89f
C396 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.08f
C397 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS 1.61f
C398 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f
C399 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS 3.25f
C400 a_1556_37246# VSS 1.16f
C401 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS 1.42f
C402 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 1.36f
C403 VREFL VSS 1.15f
C404 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.11f
C405 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].switch_n_3v3_0.D2 VSS 1.86f
C406 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.1f
C407 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f
C408 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.08f
C409 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.35f
C410 a_1556_38474# VSS 1.18f
C411 6_bit_dac_0[1].5_bit_dac_0.4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f
C412 VCC VSS 0.374p
C413 switch_n_3v3_1.D5.n0 VSS 1.4f
.ends

X1 D0 VREFL D1 D2 D3 D5 D6 D0_BUF VREFH D1_BUF D2_BUF D3_BUF
+ D5_BUF D6_BUF VOUT D4_BUF D4 VSS VCC 7_bit_dac


.param mc_mm_switch=0
.param mc_pr_switch=0
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red" tt

V1 VSS 0 dc 0
V2 VCC 0 dc 3.3

V3 VREFL 0 dc 0
V4 VREFH 0 dc 3.3

V5  D0 0 PULSE(0 1.8 4u 1p 1p 4u 8u)
V6  D1 0 PULSE(0 1.8 8u 1p 1p 8u 16u)
V7  D2 0 PULSE(0 1.8 16u 1p 1p 16u 32u)
V8  D3 0 PULSE(0 1.8 32u 1p 1p 32u 64u)
V9  D4 0 PULSE(0 1.8 64u 1p 1p 64u 128u)
V10 D5 0 PULSE(0 1.8 128u 1p 1p 128u 256u)
V11 D6 0 PULSE(0 1.8 256u 1p 1p 256u 512u)

.tran 50u 513u uic


.control
run
set filetype=ascii
set xbrushwidth=3
set hcopydevtype = svg

plot D3 D4 D5 D6 VOUT
write 7_bit_dac.raw D0 VOUT
*hardcopy 4_bit_dac_RCX.svg D0 D1 D2 D3 VOUT

.endc
.end
