magic
tech sky130A
magscale 1 2
timestamp 1687488057
<< nwell >>
rect 2852 916 3140 926
rect 2852 406 3192 916
rect 2852 398 2954 406
<< locali >>
rect 2116 -7 2170 448
<< viali >>
rect 2116 -61 2170 -7
<< metal1 >>
rect 2946 959 4381 998
rect 2946 762 2985 959
rect 4212 917 4218 924
rect 4032 878 4218 917
rect 4212 872 4218 878
rect 4270 872 4276 924
rect 4342 617 4381 959
rect -148 592 -93 598
rect -148 307 -93 537
rect -154 252 -148 307
rect -93 252 -87 307
rect -148 208 -92 214
rect -92 152 82 208
rect -148 146 -92 152
rect 2110 -7 2176 5
rect -254 -61 -248 -7
rect -194 -61 2116 -7
rect 2170 -61 2176 -7
rect 2110 -73 2176 -61
rect 2949 -102 2991 93
rect 4495 -102 4537 294
rect 2949 -144 4537 -102
<< via1 >>
rect 4218 872 4270 924
rect -148 537 -93 592
rect -148 252 -93 307
rect -148 152 -92 208
rect -248 -61 -194 -7
<< metal2 >>
rect -252 421 -197 1046
rect -148 592 -93 1046
rect 3038 910 3079 1046
rect 4218 924 4270 930
rect 4270 879 4549 918
rect 4218 866 4270 872
rect -154 537 -148 592
rect -93 537 -87 592
rect -252 366 137 421
rect -148 307 -93 313
rect -93 252 93 307
rect -148 246 -93 252
rect -252 -1 -197 188
rect -154 152 -148 208
rect -92 152 -86 208
rect -252 -7 -194 -1
rect -252 -61 -248 -7
rect -249 -182 -194 -61
rect -148 -20 -92 152
rect -148 -182 -93 -20
rect 3038 -182 3079 -67
<< metal3 >>
rect -528 728 7198 868
rect -528 38 7198 178
use /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_layout/switch2n_3v3  switch2n_3v3_0
timestamp 1687488057
transform 1 0 7554 0 1 722
box -7582 -710 -4563 214
use /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_layout/switch_n_3v3_v2  switch_n_3v3_v2_0
timestamp 1687027365
transform 1 0 9520 0 1 722
box -6614 -860 -4922 237
<< labels >>
rlabel metal3 -378 809 -378 809 7 VCC
rlabel metal3 -360 104 -360 104 7 VSS
rlabel metal2 -231 1004 -231 1004 7 D0
rlabel metal2 -120 1004 -120 1004 7 VREFL
rlabel metal2 -225 -146 -225 -146 7 D0_BUF
rlabel metal2 -117 -163 -117 -163 7 VREFH
rlabel metal2 4530 895 4530 895 7 VOUT
rlabel metal2 3060 -164 3060 -164 7 D1_BUF
rlabel metal2 3058 1022 3058 1022 7 D1
<< end >>
