magic
tech sky130A
magscale 1 2
timestamp 1692509756
<< error_p >>
rect -223 130 223 164
rect -253 -202 253 130
<< nwell >>
rect -223 -198 223 164
<< mvpmos >>
rect -129 -136 -29 64
rect 29 -136 129 64
<< mvpdiff >>
rect -187 52 -129 64
rect -187 -124 -175 52
rect -141 -124 -129 52
rect -187 -136 -129 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 129 52 187 64
rect 129 -124 141 52
rect 175 -124 187 52
rect 129 -136 187 -124
<< mvpdiffc >>
rect -175 -124 -141 52
rect -17 -124 17 52
rect 141 -124 175 52
<< poly >>
rect -129 145 -29 161
rect -129 111 -113 145
rect -45 111 -29 145
rect -129 64 -29 111
rect 29 145 129 161
rect 29 111 45 145
rect 113 111 129 145
rect 29 64 129 111
rect -129 -162 -29 -136
rect 29 -162 129 -136
<< polycont >>
rect -113 111 -45 145
rect 45 111 113 145
<< locali >>
rect -129 111 -113 145
rect -45 111 -29 145
rect 29 111 45 145
rect 113 111 129 145
rect -175 52 -141 68
rect -175 -140 -141 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 141 52 175 68
rect 141 -140 175 -124
<< viali >>
rect -113 111 -45 145
rect 45 111 113 145
rect -175 -124 -141 52
rect -17 -124 17 52
rect 141 -124 175 52
<< metal1 >>
rect -125 145 -33 151
rect -125 111 -113 145
rect -45 111 -33 145
rect -125 105 -33 111
rect 33 145 125 151
rect 33 111 45 145
rect 113 111 125 145
rect 33 105 125 111
rect -181 52 -135 64
rect -181 -124 -175 52
rect -141 -124 -135 52
rect -181 -136 -135 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 135 52 181 64
rect 135 -124 141 52
rect 175 -124 181 52
rect 135 -136 181 -124
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
