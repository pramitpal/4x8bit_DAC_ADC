** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/2bitdac/2_bit_dac.sch
.subckt 2_bit_dac D1 D0 D0_BUF D1_BUF VOUT VREFL VREFH VCC VSS
*.PININFO D1:I D0:I D0_BUF:O D1_BUF:O VOUT:O VREFL:I VREFH:I VCC:B VSS:B
x1 VCC D0_BUF D0 VREFH VSS VINL VINH VREFL switch2n_3v3
x2 VCC D1 D1_BUF VSS VINH VOUT VINL switch_n_3v3
.ends

* expanding   symbol:
*+  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch2n_3v3.sym # of pins=8
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch2n_3v3.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch2n_3v3.sch
.subckt switch2n_3v3 VCC DX_BUF DX VREFH VSS VOUTL VOUTH VREFL
*.PININFO VCC:B VSS:B VOUTL:O DX:I VOUTH:O DX_BUF:O VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUTL net1 VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUTL net1 net2 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 net2 DX_BUF VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM9 VOUTH net1 net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM10 VOUTH net1 net4 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM11 net3 DX_BUF VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM12 net4 DX_BUF VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XR1 net3 net4 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR2 net2 net3 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR3 VREFL net2 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR4 net4 VREFH VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch_n_3v3.sym # of pins=7
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch_n_3v3.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch_n_3v3.sch
.subckt switch_n_3v3 VCC DX DX_BUF VSS VREFH VOUT VREFL
*.PININFO VCC:B VSS:B DX_BUF:O VOUT:O DX:I VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUT net1 VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUT net1 VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 VREFH DX_BUF VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends

.end
