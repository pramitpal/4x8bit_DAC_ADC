* NGSPICE file created from 4x8_bit_dac.ext - technology: sky130A

.subckt switch_n_3v3_v2 VREFH DX_BUF DX VCC VSS VOUT VREFL
X0 VOUT DX_BUF VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 DX_ DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 DX_BUF DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT DX_BUF VREFL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 DX_ DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 VREFL DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 DX_BUF DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VREFH DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt switch2n_3v3 VOUTL DX_BUF VREFH VOUTH DX VCC VSS VREFL
X0 VOUTH a_n6524_n498# a_n7536_n67# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 a_n7536_n67# DX_BUF VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2 a_n7536_n67# R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3 DX_BUF a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4 VREFL DX_BUF VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X5 a_n7536_n67# VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6 a_n6524_n498# DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VOUTL a_n6524_n498# VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8 VOUTH a_n6524_n498# R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 R_H DX_BUF VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 R_H R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X11 R_L VREFL VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X12 R_L DX_BUF VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 DX_BUF a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 a_n6524_n498# DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X15 VOUTL a_n6524_n498# R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt x2_bit_dac VREFH D1_BUF D1 D0 VCC D0_BUF VOUT VREFL VSS
Xswitch_n_3v3_v2_0 switch2n_3v3_0/VOUTH D1_BUF D1 VCC VSS VOUT switch2n_3v3_0/VOUTL
+ switch_n_3v3_v2
Xswitch2n_3v3_0 switch2n_3v3_0/VOUTL D0_BUF VREFH switch2n_3v3_0/VOUTH D0 VCC VSS
+ VREFL switch2n_3v3
.ends

.subckt switch_n_3v3 VREFH DX_BUF m2_n6802_n990# m2_n6562_n990# D7 D6 D5 D4 DX m2_n6722_n990#
+ D3 D2 m2_n6482_n990# m2_n6882_n990# VCC VSS VOUT m2_n6642_n990# VREFL
X0 VOUT DX_BUF VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 DX_ DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 DX_BUF DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT DX_BUF VREFL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 DX_ DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 VREFL DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 DX_BUF DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VREFH DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt x3_bit_dac VREFH D1_BUF switch_n_3v3_1/D6 switch_n_3v3_1/D7 switch_n_3v3_1/D3
+ D2_BUF switch_n_3v3_1/D4 D2 D1 D0 D0_BUF VCC VOUT VREFL switch_n_3v3_1/D5 VSS
X2_bit_dac_0[0] VREFH D1_BUF 2_bit_dac_0[0]/D1 2_bit_dac_0[0]/D0 VCC D0_BUF 2_bit_dac_0[0]/VOUT
+ 2_bit_dac_0[1]/VREFH VSS x2_bit_dac
X2_bit_dac_0[1] 2_bit_dac_0[1]/VREFH 2_bit_dac_0[0]/D1 D1 D0 VCC 2_bit_dac_0[0]/D0
+ 2_bit_dac_0[1]/VOUT VREFL VSS x2_bit_dac
Xswitch_n_3v3_1 2_bit_dac_0[0]/VOUT D2_BUF switch_n_3v3_1/D3 switch_n_3v3_1/D6 switch_n_3v3_1/D7
+ switch_n_3v3_1/D6 switch_n_3v3_1/D5 switch_n_3v3_1/D4 D2 switch_n_3v3_1/D4 switch_n_3v3_1/D3
+ D2 switch_n_3v3_1/D7 D2_BUF VCC VSS VOUT switch_n_3v3_1/D5 2_bit_dac_0[1]/VOUT switch_n_3v3
.ends

.subckt x4_bit_dac VREFH D1_BUF D2_BUF D3 D2 switch_n_3v3_0/D7 D1 switch_n_3v3_0/D6
+ D0 switch_n_3v3_0/D5 switch_n_3v3_0/D4 D3_BUF D0_BUF VCC VOUT VREFL VSS
X3_bit_dac_0[0] VREFH D1_BUF switch_n_3v3_0/D6 switch_n_3v3_0/D7 D3_BUF D2_BUF switch_n_3v3_0/D4
+ switch_n_3v3_0/D2 3_bit_dac_0[0]/D1 3_bit_dac_0[0]/D0 D0_BUF VCC 3_bit_dac_0[0]/VOUT
+ 3_bit_dac_0[1]/VREFH switch_n_3v3_0/D5 VSS x3_bit_dac
X3_bit_dac_0[1] 3_bit_dac_0[1]/VREFH 3_bit_dac_0[0]/D1 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ D3 switch_n_3v3_0/D2 switch_n_3v3_0/D4 D2 D1 D0 3_bit_dac_0[0]/D0 VCC 3_bit_dac_0[1]/VOUT
+ VREFL switch_n_3v3_0/D5 VSS x3_bit_dac
Xswitch_n_3v3_0 3_bit_dac_0[0]/VOUT D3_BUF D3_BUF switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 switch_n_3v3_0/D5 switch_n_3v3_0/D4 D3 switch_n_3v3_0/D4 D3 switch_n_3v3_0/D2
+ switch_n_3v3_0/D7 switch_n_3v3_0/D2 VCC VSS VOUT switch_n_3v3_0/D5 3_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt x5_bit_dac D4_BUF VREFH D1_BUF D2_BUF D4 D3 D2 D1 switch_n_3v3_0/D6 D0 D3_BUF
+ switch_n_3v3_0/D7 D0_BUF VOUT VCC VREFL switch_n_3v3_0/D5 VSS
X4_bit_dac_0[0] VREFH D1_BUF D2_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D2 switch_n_3v3_0/D7
+ 4_bit_dac_0[0]/D1 switch_n_3v3_0/D6 4_bit_dac_0[0]/D0 switch_n_3v3_0/D5 D4_BUF D3_BUF
+ D0_BUF VCC 4_bit_dac_0[0]/VOUT 4_bit_dac_0[1]/VREFH VSS x4_bit_dac
X4_bit_dac_0[1] 4_bit_dac_0[1]/VREFH 4_bit_dac_0[0]/D1 switch_n_3v3_0/D2 D3 D2 switch_n_3v3_0/D7
+ D1 switch_n_3v3_0/D6 D0 switch_n_3v3_0/D5 D4 switch_n_3v3_0/D3 4_bit_dac_0[0]/D0
+ VCC 4_bit_dac_0[1]/VOUT VREFL VSS x4_bit_dac
Xswitch_n_3v3_0 4_bit_dac_0[0]/VOUT D4_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 switch_n_3v3_0/D5 D4 D4 D4_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D2
+ switch_n_3v3_0/D7 switch_n_3v3_0/D2 VCC VSS VOUT switch_n_3v3_0/D5 4_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt x6_bit_dac D0 D1 D2 D5 VREFH VREFL D0_BUF D1_BUF D2_BUF D5_BUF VOUT VCC D3
+ D3_BUF D4 D4_BUF switch_n_3v3_0/D7 switch_n_3v3_0/D6 VSS
X5_bit_dac_1 D4_BUF VREFH D1_BUF D2_BUF 5_bit_dac_1/D4 5_bit_dac_1/D3 5_bit_dac_1/D2
+ 5_bit_dac_1/D1 switch_n_3v3_0/D6 5_bit_dac_1/D0 D3_BUF switch_n_3v3_0/D7 D0_BUF
+ 5_bit_dac_1/VOUT VCC 5_bit_dac_1/VREFL D5_BUF VSS x5_bit_dac
Xswitch_n_3v3_0 5_bit_dac_1/VOUT D5_BUF 5_bit_dac_1/D3 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 D5 5_bit_dac_1/D4 D5 5_bit_dac_1/D4 5_bit_dac_1/D3 5_bit_dac_1/D2
+ switch_n_3v3_0/D7 5_bit_dac_1/D2 VCC VSS VOUT D5_BUF 5_bit_dac_0/VOUT switch_n_3v3
X5_bit_dac_0 5_bit_dac_1/D4 5_bit_dac_1/VREFL 5_bit_dac_1/D1 5_bit_dac_1/D2 D4 D3
+ D2 D1 switch_n_3v3_0/D6 D0 5_bit_dac_1/D3 switch_n_3v3_0/D7 5_bit_dac_1/D0 5_bit_dac_0/VOUT
+ VCC VREFL D5 VSS x5_bit_dac
.ends

.subckt x7_bit_dac VREFH D1_BUF D6 D5 D4 D3 D2 D1 D0 D4_BUF D3_BUF VCC D0_BUF VOUT
+ switch_n_3v3_1/D7 D6_BUF D5_BUF VREFL VSS D2_BUF
X6_bit_dac_0[0] 6_bit_dac_0[0]/D0 6_bit_dac_0[0]/D1 switch_n_3v3_1/D2 switch_n_3v3_1/D5
+ VREFH 6_bit_dac_0[1]/VREFH D0_BUF D1_BUF D2_BUF D5_BUF 6_bit_dac_0[0]/VOUT VCC switch_n_3v3_1/D3
+ D3_BUF switch_n_3v3_1/D4 D4_BUF switch_n_3v3_1/D7 D6_BUF VSS x6_bit_dac
X6_bit_dac_0[1] D0 D1 D2 D5 6_bit_dac_0[1]/VREFH VREFL 6_bit_dac_0[0]/D0 6_bit_dac_0[0]/D1
+ switch_n_3v3_1/D2 switch_n_3v3_1/D5 6_bit_dac_0[1]/VOUT VCC D3 switch_n_3v3_1/D3
+ D4 switch_n_3v3_1/D4 switch_n_3v3_1/D7 D6 VSS x6_bit_dac
Xswitch_n_3v3_1 6_bit_dac_0[0]/VOUT D6_BUF switch_n_3v3_1/D3 D6_BUF switch_n_3v3_1/D7
+ D6 switch_n_3v3_1/D5 switch_n_3v3_1/D4 D6 switch_n_3v3_1/D4 switch_n_3v3_1/D3 switch_n_3v3_1/D2
+ switch_n_3v3_1/D7 switch_n_3v3_1/D2 VCC VSS VOUT switch_n_3v3_1/D5 6_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt x8_bit_dac VREFH D7 D6 D5 D4 D3 D2 D0 D1 VOUT VREFL VCC VSS
X7_bit_dac_0 7_bit_dac_1/VREFL 7_bit_dac_1/D1 D6 D5 D4 D3 D2 D1 D0 7_bit_dac_1/D4
+ 7_bit_dac_1/D3 VCC 7_bit_dac_1/D0 7_bit_dac_0/VOUT D7 7_bit_dac_1/D6 7_bit_dac_1/D5
+ VREFL VSS 7_bit_dac_1/D2 x7_bit_dac
X7_bit_dac_1 VREFH D1_BUF 7_bit_dac_1/D6 7_bit_dac_1/D5 7_bit_dac_1/D4 7_bit_dac_1/D3
+ 7_bit_dac_1/D2 7_bit_dac_1/D1 7_bit_dac_1/D0 D4_BUF D3_BUF VCC D0_BUF 7_bit_dac_1/VOUT
+ D7_BUF D6_BUF D5_BUF 7_bit_dac_1/VREFL VSS D2_BUF x7_bit_dac
Xswitch_n_3v3_1 7_bit_dac_1/VOUT D7_BUF 7_bit_dac_1/D3 7_bit_dac_1/D6 D7 7_bit_dac_1/D6
+ 7_bit_dac_1/D5 7_bit_dac_1/D4 D7 7_bit_dac_1/D4 7_bit_dac_1/D3 7_bit_dac_1/D2 D7_BUF
+ 7_bit_dac_1/D2 VCC VSS VOUT 7_bit_dac_1/D5 7_bit_dac_0/VOUT switch_n_3v3
.ends

.subckt level_tx_1bit VCCD VSSD VIN VOUT VDDA
X0 a_n1423_1248# VOUT VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 VSSD VIN a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.2
X2 VSSD VIN a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4 a_n1353_675# VIN VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.2
X5 VOUT a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt level_tx_8bit VIN7 VIN6 VIN5 VIN4 VIN3 VIN2 VIN1 VIN0 VCCD VOUT7 VSSD VOUT6
+ VOUT5 VOUT4 VOUT3 VOUT2 VOUT1 VOUT0 VDDA
Xlevel_tx_1bit_0[0] VCCD VSSD VIN0 VOUT0 VDDA level_tx_1bit
Xlevel_tx_1bit_0[1] VCCD VSSD VIN1 VOUT1 VDDA level_tx_1bit
Xlevel_tx_1bit_0[2] VCCD VSSD VIN2 VOUT2 VDDA level_tx_1bit
Xlevel_tx_1bit_0[3] VCCD VSSD VIN3 VOUT3 VDDA level_tx_1bit
Xlevel_tx_1bit_0[4] VCCD VSSD VIN4 VOUT4 VDDA level_tx_1bit
Xlevel_tx_1bit_0[5] VCCD VSSD VIN5 VOUT5 VDDA level_tx_1bit
Xlevel_tx_1bit_0[6] VCCD VSSD VIN6 VOUT6 VDDA level_tx_1bit
Xlevel_tx_1bit_0[7] VCCD VSSD VIN7 VOUT7 VDDA level_tx_1bit
.ends

.subckt opamp VSSA VIN VOUT VDDA
X0 VSSA a_3246_n774# VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X1 VOUT a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 VDDA a_1618_n334# VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X3 VDDA a_394_n920# a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X4 a_1704_376# VOUT a_1446_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X5 VDDA a_1618_n334# VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X6 a_408_552# VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.48 l=4.46
X7 VSSA a_1022_n914# a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X8 a_2158_n774# VOUT a_1900_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X9 VSSA a_2894_292# a_2894_292# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X10 a_1022_n914# a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X11 a_1776_n834# a_408_552# a_1618_n334# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X12 VSSA a_1022_n914# a_1446_376# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X13 a_2894_292# a_408_552# a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X14 VDDA a_408_552# VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=8.32
X15 a_2416_n774# a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X16 VDDA a_394_n920# a_394_n920# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
X17 a_1446_376# a_408_552# a_1300_n354# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X18 VOUT a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X19 a_2416_n774# VIN a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X20 VOUT a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
X21 VOUT a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X22 a_1776_n834# VIN a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X23 a_1618_n334# a_1300_n354# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X24 VSSA a_3246_n774# VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X25 VSSA a_1022_n914# a_1022_n914# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X26 a_1776_n834# a_1022_n914# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X27 a_3246_n774# a_2894_292# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X28 VSSA a_394_n920# VSSA sky130_fd_pr__res_generic_nd__hv w=0.41 l=15.7
X29 VDDA a_394_n920# a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X30 a_3246_n774# a_408_552# a_2416_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X31 VDDA a_1300_n354# a_1300_n354# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
.ends

.subckt x8_bit_dac_tx_buffer VREFH VCCD D7 D6 D5 D4 D3 D2 D1 D0 VOUT_BUF VSSD VSSA
+ VDDA
X8_bit_dac_0 VREFH 8_bit_dac_0/D7 8_bit_dac_0/D6 8_bit_dac_0/D5 8_bit_dac_0/D4 8_bit_dac_0/D3
+ 8_bit_dac_0/D2 8_bit_dac_0/D0 8_bit_dac_0/D1 VOUT VSSA VDDA VSSA x8_bit_dac
Xlevel_tx_8bit_0 D7 D6 D5 D4 D3 D2 D1 D0 VCCD 8_bit_dac_0/D7 VSSD 8_bit_dac_0/D6 8_bit_dac_0/D5
+ 8_bit_dac_0/D4 8_bit_dac_0/D3 8_bit_dac_0/D2 8_bit_dac_0/D1 8_bit_dac_0/D0 VDDA
+ level_tx_8bit
Xopamp_0 VSSA VOUT VOUT_BUF VDDA opamp
.ends

.subckt x4x8_bit_dac Din0[0] Din0[1] Din0[2] Din0[3] Din0[4] Din0[5] Din0[6] Din0[7]
+ VOUT0 Din1[0] Din1[1] Din1[2] Din1[3] Din1[4] Din1[5] Din1[6] Din1[7] VOUT1 Din2[0]
+ Din2[1] Din2[2] Din2[3] Din2[4] Din2[5] Din2[6] Din2[7] VOUT2 Din3[0] Din3[1] Din3[2]
+ Din3[3] Din3[4] Din3[5] Din3[6] Din3[7] VOUT3 VDDA VSSA VSSD VCCD VREFH
X8_bit_dac_tx_buffer_0[0] VREFH VCCD Din0[7] Din0[6] Din0[5] Din0[4] Din0[3] Din0[2]
+ Din0[1] Din0[0] VOUT0 VSSD VSSA VDDA x8_bit_dac_tx_buffer
X8_bit_dac_tx_buffer_0[1] VREFH VCCD Din1[7] Din1[6] Din1[5] Din1[4] Din1[3] Din1[2]
+ Din1[1] Din1[0] VOUT1 VSSD VSSA VDDA x8_bit_dac_tx_buffer
X8_bit_dac_tx_buffer_0[2] VREFH VCCD Din2[7] Din2[6] Din2[5] Din2[4] Din2[3] Din2[2]
+ Din2[1] Din2[0] VOUT2 VSSD VSSA VDDA x8_bit_dac_tx_buffer
X8_bit_dac_tx_buffer_0[3] VREFH VCCD Din3[7] Din3[6] Din3[5] Din3[4] Din3[3] Din3[2]
+ Din3[1] Din3[0] VOUT3 VSSD VSSA VDDA x8_bit_dac_tx_buffer
.ends

