magic
tech sky130A
magscale 1 2
timestamp 1692514852
<< nwell >>
rect 670 638 2433 1085
rect 671 250 2433 638
rect 671 -22 2100 250
rect 671 -80 1910 -22
<< mvpsubdiff >>
rect 755 -479 2487 -458
rect 755 -546 784 -479
rect 2441 -546 2487 -479
rect 755 -564 2487 -546
<< mvnsubdiff >>
rect 884 901 2351 919
rect 884 833 912 901
rect 2327 833 2351 901
rect 884 813 2351 833
<< mvpsubdiffcont >>
rect 784 -546 2441 -479
<< mvnsubdiffcont >>
rect 912 833 2327 901
<< poly >>
rect 2156 316 2256 350
rect 2156 282 2172 316
rect 2240 282 2256 316
rect 2156 272 2256 282
rect 2557 238 2657 254
rect 2557 204 2573 238
rect 2641 204 2657 238
rect 2557 174 2657 204
rect 962 -31 1062 65
rect 804 -61 904 -45
rect 804 -95 814 -61
rect 894 -95 904 -61
rect 804 -134 904 -95
rect 962 -65 972 -31
rect 1052 -65 1062 -31
rect 1529 24 1629 40
rect 1529 -10 1539 24
rect 1619 -10 1629 24
rect 962 -157 1062 -65
rect 1250 -75 1350 -59
rect 1250 -109 1260 -75
rect 1340 -109 1350 -75
rect 1250 -133 1350 -109
rect 1529 -152 1629 -10
rect 1687 -40 1787 -24
rect 1687 -74 1697 -40
rect 1777 -74 1787 -40
rect 1687 -166 1787 -74
rect 1845 -30 1945 88
rect 1845 -64 1872 -30
rect 1906 -64 1945 -30
rect 1845 -159 1945 -64
<< polycont >>
rect 2172 282 2240 316
rect 2573 204 2641 238
rect 814 -95 894 -61
rect 972 -65 1052 -31
rect 1539 -10 1619 24
rect 1260 -109 1340 -75
rect 1697 -74 1777 -40
rect 1872 -64 1906 -30
<< locali >>
rect 860 901 2365 936
rect 860 833 912 901
rect 2327 833 2365 901
rect 860 796 2365 833
rect 2156 282 2172 316
rect 2240 282 2256 316
rect 789 33 823 110
rect 789 8 1067 33
rect 1440 8 1474 273
rect 2557 204 2573 238
rect 2641 204 2657 238
rect 1542 152 1597 186
rect 1542 118 1552 152
rect 1586 118 1597 152
rect 1542 63 1597 118
rect 1541 44 1597 63
rect 1529 38 1629 44
rect 789 -1 1474 8
rect 952 -26 1474 -1
rect 1522 24 1635 38
rect 1522 -10 1539 24
rect 1619 -10 1635 24
rect 1522 -20 1635 -10
rect 952 -31 1067 -26
rect 1529 -31 1629 -20
rect 1679 -26 1793 -17
rect 800 -47 910 -41
rect 798 -61 829 -47
rect 887 -61 910 -47
rect 798 -95 814 -61
rect 894 -95 910 -61
rect 952 -65 972 -31
rect 1052 -65 1067 -31
rect 1679 -40 1712 -26
rect 1770 -40 1793 -26
rect 952 -81 1067 -65
rect 1243 -74 1354 -61
rect 1679 -74 1697 -40
rect 1777 -74 1793 -40
rect 1856 -64 1872 -30
rect 1907 -64 1922 -30
rect 1243 -75 1517 -74
rect 798 -105 829 -95
rect 887 -105 910 -95
rect 800 -112 910 -105
rect 1243 -109 1260 -75
rect 1340 -109 1482 -75
rect 1243 -119 1354 -109
rect 1679 -84 1712 -74
rect 1770 -84 1793 -74
rect 1679 -92 1793 -84
rect 1482 -118 1517 -110
rect 687 -479 2544 -444
rect 687 -546 784 -479
rect 2441 -546 2544 -479
rect 687 -584 2544 -546
<< viali >>
rect 912 833 2327 901
rect 1440 273 1474 307
rect 2172 282 2240 316
rect 789 110 823 144
rect 2573 204 2641 238
rect 1552 118 1586 152
rect 829 -61 887 -47
rect 829 -95 887 -61
rect 1712 -40 1770 -26
rect 1872 -30 1907 -29
rect 1712 -74 1770 -40
rect 1872 -64 1906 -30
rect 1906 -64 1907 -30
rect 829 -105 887 -95
rect 1482 -110 1517 -75
rect 1712 -84 1770 -74
rect 784 -546 2441 -479
<< metal1 >>
rect 808 901 2365 936
rect 808 833 912 901
rect 2327 833 2365 901
rect 808 796 2365 833
rect 808 541 854 796
rect 976 668 1028 674
rect 960 619 976 665
rect 1467 624 1993 659
rect 976 610 1028 616
rect 1418 559 1453 576
rect 808 495 956 541
rect 1404 507 1410 559
rect 1462 507 1468 559
rect 910 248 956 495
rect 1059 437 1065 489
rect 1117 437 1123 489
rect 1068 402 1114 437
rect 1418 404 1453 507
rect 1578 466 1612 578
rect 1737 560 1772 576
rect 1722 508 1728 560
rect 1780 508 1786 560
rect 1563 414 1569 466
rect 1621 414 1627 466
rect 1068 289 1336 335
rect 1434 308 1480 319
rect 1629 308 1635 317
rect 1434 307 1635 308
rect 901 196 907 248
rect 959 196 965 248
rect 783 153 829 156
rect 774 101 780 153
rect 832 101 838 153
rect 783 98 829 101
rect 823 -41 893 -35
rect 817 -111 823 -41
rect 881 -47 893 -41
rect 887 -105 893 -47
rect 881 -111 893 -105
rect 823 -117 893 -111
rect 1068 -204 1114 289
rect 1434 273 1440 307
rect 1474 274 1635 307
rect 1474 273 1480 274
rect 1434 261 1480 273
rect 1629 265 1635 274
rect 1687 265 1693 317
rect 1210 163 1235 201
rect 1186 111 1192 163
rect 1248 111 1254 163
rect 1360 129 1395 196
rect 1958 179 1993 624
rect 2110 528 2144 796
rect 2259 490 2311 496
rect 2311 447 2318 481
rect 2259 432 2311 438
rect 2132 327 2226 328
rect 2131 321 2348 327
rect 2191 316 2348 321
rect 2240 282 2348 316
rect 2191 261 2348 282
rect 2131 255 2191 261
rect 2274 244 2348 261
rect 2274 238 2653 244
rect 2274 204 2573 238
rect 2641 204 2653 238
rect 2274 198 2653 204
rect 1546 164 1598 170
rect 1201 86 1240 111
rect 1360 94 1517 129
rect 1598 112 1835 158
rect 1546 106 1598 112
rect 1482 -69 1517 94
rect 1549 88 1595 106
rect 1706 -20 1776 -14
rect 1470 -75 1529 -69
rect 1470 -110 1482 -75
rect 1517 -110 1529 -75
rect 1700 -90 1706 -20
rect 1764 -26 1776 -20
rect 1864 -20 1916 -14
rect 1770 -84 1776 -26
rect 1860 -70 1864 -23
rect 1916 -70 1919 -23
rect 1864 -78 1916 -72
rect 1764 -90 1776 -84
rect 1706 -96 1776 -90
rect 1470 -116 1529 -110
rect 1068 -250 1241 -204
rect 1482 -235 1517 -116
rect 1951 -183 1997 138
rect 2392 90 2426 143
rect 2121 64 2181 70
rect 2181 4 2265 64
rect 2377 38 2383 90
rect 2435 38 2441 90
rect 2495 66 2501 118
rect 2553 66 2559 118
rect 2121 -2 2181 4
rect 2510 -11 2544 66
rect 2464 -74 2524 -68
rect 2099 -121 2464 -86
rect 2309 -122 2464 -121
rect 2464 -140 2524 -134
rect 2234 -192 2268 -169
rect 2669 -176 2703 -21
rect 900 -309 906 -257
rect 958 -309 964 -257
rect 1347 -309 1353 -257
rect 1405 -309 1411 -257
rect 1468 -287 1474 -235
rect 1526 -287 1532 -235
rect 2219 -244 2225 -192
rect 2277 -244 2283 -192
rect 2478 -210 2703 -176
rect 2061 -324 2067 -272
rect 2119 -324 2125 -272
rect 757 -444 792 -338
rect 1799 -444 1833 -348
rect 2076 -349 2110 -324
rect 2234 -363 2268 -251
rect 2392 -272 2426 -266
rect 2377 -324 2383 -272
rect 2435 -324 2441 -272
rect 2478 -444 2512 -210
rect 687 -479 2544 -444
rect 687 -546 784 -479
rect 2441 -546 2544 -479
rect 687 -584 2544 -546
<< via1 >>
rect 912 833 2327 901
rect 976 616 1028 668
rect 1410 507 1462 559
rect 1065 437 1117 489
rect 1728 508 1780 560
rect 1569 414 1621 466
rect 907 196 959 248
rect 780 144 832 153
rect 780 110 789 144
rect 789 110 823 144
rect 823 110 832 144
rect 780 101 832 110
rect 823 -47 881 -41
rect 823 -105 829 -47
rect 829 -105 881 -47
rect 823 -111 881 -105
rect 1635 265 1687 317
rect 1192 111 1248 163
rect 2259 438 2311 490
rect 2131 316 2191 321
rect 2131 282 2172 316
rect 2172 282 2191 316
rect 2131 261 2191 282
rect 1546 152 1598 164
rect 1546 118 1552 152
rect 1552 118 1586 152
rect 1586 118 1598 152
rect 1546 112 1598 118
rect 1706 -26 1764 -20
rect 1706 -84 1712 -26
rect 1712 -84 1764 -26
rect 1864 -29 1916 -20
rect 1864 -64 1872 -29
rect 1872 -64 1907 -29
rect 1907 -64 1916 -29
rect 1864 -72 1916 -64
rect 1706 -90 1764 -84
rect 2121 4 2181 64
rect 2383 38 2435 90
rect 2501 66 2553 118
rect 2464 -134 2524 -74
rect 906 -309 958 -257
rect 1353 -309 1405 -257
rect 1474 -287 1526 -235
rect 2225 -244 2277 -192
rect 2067 -324 2119 -272
rect 2383 -324 2435 -272
rect 784 -546 2441 -479
<< metal2 >>
rect 684 1046 693 1106
rect 753 1046 762 1106
rect 700 486 746 1046
rect 860 901 2365 936
rect 860 833 912 901
rect 2327 833 2365 901
rect 860 796 2365 833
rect 800 714 1456 753
rect 800 612 839 714
rect 972 672 1032 681
rect 970 616 972 668
rect 1032 616 1034 668
rect 790 603 850 612
rect 972 603 1032 612
rect 1417 565 1456 714
rect 790 534 850 543
rect 1410 559 1462 565
rect 1728 560 1780 566
rect 1462 516 1728 555
rect 1065 489 1117 495
rect 700 440 1065 486
rect 1190 493 1250 502
rect 1410 501 1462 507
rect 1780 521 2079 555
rect 1728 502 1780 508
rect 1117 440 1190 486
rect 1065 431 1117 437
rect 1190 424 1250 433
rect 1569 466 1621 472
rect 1621 423 2014 457
rect 1569 408 1621 414
rect 792 391 848 400
rect 603 342 792 385
rect 792 326 848 335
rect 1635 321 1687 323
rect 1622 261 1631 321
rect 1691 261 1700 321
rect 1635 259 1687 261
rect 907 248 959 254
rect 959 199 1489 245
rect 907 190 959 196
rect 1192 167 1248 169
rect 780 153 832 159
rect 626 110 780 144
rect 1183 111 1192 167
rect 1248 111 1257 167
rect 1443 161 1489 199
rect 1540 161 1546 164
rect 1443 115 1546 161
rect 1540 112 1546 115
rect 1598 112 1604 164
rect 1696 131 1705 191
rect 1765 131 1774 191
rect 1192 105 1248 111
rect 780 95 832 101
rect 1340 57 1349 64
rect 697 11 1349 57
rect 697 -260 743 11
rect 1340 4 1349 11
rect 1409 4 1418 64
rect 1706 -20 1764 131
rect 815 -41 899 -32
rect 815 -111 823 -41
rect 881 -111 899 -41
rect 1691 -90 1706 -24
rect 1764 -26 1778 -24
rect 1764 -84 1794 -26
rect 1858 -72 1864 -20
rect 1916 -72 1922 -20
rect 1764 -90 1778 -84
rect 1691 -97 1778 -90
rect 815 -133 899 -111
rect 1706 -133 1764 -97
rect 815 -191 1764 -133
rect 1471 -230 1531 -221
rect 906 -257 958 -251
rect 697 -306 906 -260
rect 1353 -257 1405 -251
rect 958 -306 1353 -260
rect 906 -315 958 -309
rect 1873 -243 1908 -72
rect 1531 -278 1908 -243
rect 1471 -299 1531 -290
rect 1980 -281 2014 423
rect 2045 -201 2079 521
rect 2253 438 2259 490
rect 2311 438 2317 490
rect 2133 321 2189 328
rect 2125 261 2131 321
rect 2191 261 2197 321
rect 2133 254 2189 261
rect 2115 191 2171 198
rect 2113 190 2179 191
rect 2268 190 2302 438
rect 2113 189 2544 190
rect 2113 133 2115 189
rect 2171 156 2544 189
rect 2171 133 2179 156
rect 2113 131 2179 133
rect 2115 124 2171 131
rect 2510 124 2544 156
rect 2501 118 2553 124
rect 2383 90 2435 96
rect 2123 64 2179 71
rect 2115 4 2121 64
rect 2181 4 2187 64
rect 2501 60 2553 66
rect 2383 32 2435 38
rect 2123 -3 2179 4
rect 2392 -76 2426 32
rect 2466 -74 2522 -67
rect 2235 -110 2426 -76
rect 2235 -186 2269 -110
rect 2458 -134 2464 -74
rect 2524 -134 2530 -74
rect 2466 -141 2522 -134
rect 2225 -192 2277 -186
rect 2045 -235 2225 -201
rect 2277 -235 2288 -201
rect 2225 -250 2277 -244
rect 2067 -272 2119 -266
rect 1353 -315 1405 -309
rect 1980 -315 2067 -281
rect 2383 -272 2435 -266
rect 2119 -315 2383 -281
rect 2067 -330 2119 -324
rect 2435 -315 2941 -281
rect 2383 -330 2435 -324
rect 687 -479 2544 -444
rect 687 -546 784 -479
rect 2441 -546 2544 -479
rect 687 -584 2544 -546
rect 2679 -676 2713 -315
rect 2666 -685 2726 -676
rect 2666 -754 2726 -745
<< via2 >>
rect 693 1046 753 1106
rect 912 833 2327 901
rect 972 668 1032 672
rect 972 616 976 668
rect 976 616 1028 668
rect 1028 616 1032 668
rect 972 612 1032 616
rect 790 543 850 603
rect 1190 433 1250 493
rect 792 335 848 391
rect 1631 317 1691 321
rect 1631 265 1635 317
rect 1635 265 1687 317
rect 1687 265 1691 317
rect 1631 261 1691 265
rect 1192 163 1248 167
rect 1192 111 1248 163
rect 1705 131 1765 191
rect 1349 4 1409 64
rect 1471 -235 1531 -230
rect 1471 -287 1474 -235
rect 1474 -287 1526 -235
rect 1526 -287 1531 -235
rect 1471 -290 1531 -287
rect 2133 263 2189 319
rect 2115 133 2171 189
rect 2123 6 2179 62
rect 2466 -132 2522 -76
rect 784 -546 2441 -479
rect 2666 -745 2726 -685
<< metal3 >>
rect 688 1106 758 1111
rect 1558 1108 1622 1114
rect 688 1046 693 1106
rect 753 1046 1558 1106
rect 688 1041 758 1046
rect 1558 1038 1622 1044
rect 460 901 3028 936
rect 460 833 912 901
rect 2327 833 3028 901
rect 460 796 3028 833
rect 960 672 1044 678
rect 960 612 972 672
rect 1032 612 1044 672
rect 2837 619 2901 625
rect 785 603 855 608
rect 960 604 1044 612
rect 785 543 790 603
rect 850 543 855 603
rect 785 538 855 543
rect 790 396 850 538
rect 787 391 853 396
rect 787 335 792 391
rect 848 335 853 391
rect 787 330 853 335
rect 980 -74 1040 604
rect 2428 557 2837 617
rect 1185 493 1255 498
rect 1185 433 1190 493
rect 1250 433 1255 493
rect 1185 428 1255 433
rect 1190 172 1250 428
rect 1626 321 1696 326
rect 2128 321 2194 324
rect 1626 261 1631 321
rect 1691 319 2194 321
rect 1691 263 2133 319
rect 2189 263 2194 319
rect 1691 261 2194 263
rect 1626 256 1696 261
rect 2128 258 2194 261
rect 1700 191 1770 196
rect 2110 191 2176 194
rect 1187 167 1253 172
rect 1187 111 1192 167
rect 1248 111 1253 167
rect 1700 131 1705 191
rect 1765 189 2176 191
rect 1765 133 2115 189
rect 2171 133 2176 189
rect 1765 131 2176 133
rect 1700 126 1770 131
rect 2110 128 2176 131
rect 1187 106 1253 111
rect 1344 64 1414 69
rect 2118 64 2184 67
rect 2428 64 2488 557
rect 2837 549 2901 555
rect 1344 4 1349 64
rect 1409 62 2488 64
rect 1409 6 2123 62
rect 2179 6 2488 62
rect 1409 4 2488 6
rect 1344 -1 1414 4
rect 2118 1 2184 4
rect 2461 -74 2527 -71
rect 980 -76 2527 -74
rect 980 -132 2466 -76
rect 2522 -132 2527 -76
rect 980 -134 2527 -132
rect 1471 -225 1531 -134
rect 2461 -137 2527 -134
rect 1466 -230 1536 -225
rect 1466 -290 1471 -230
rect 1531 -290 1536 -230
rect 1466 -295 1536 -290
rect 628 -479 2934 -444
rect 628 -546 784 -479
rect 2441 -546 2934 -479
rect 628 -584 2934 -546
rect 1567 -683 1631 -677
rect 2661 -685 2731 -680
rect 1631 -745 2666 -685
rect 2726 -745 2731 -685
rect 2830 -720 2934 -584
rect 1567 -753 1631 -747
rect 2661 -750 2731 -745
rect 2825 -822 2831 -720
rect 2933 -822 2939 -720
rect 2830 -823 2934 -822
rect 460 -1122 3028 -982
<< via3 >>
rect 1558 1044 1622 1108
rect 2837 555 2901 619
rect 1567 -747 1631 -683
rect 2831 -822 2933 -720
<< metal4 >>
rect 1560 1132 1620 1223
rect 1536 1108 1640 1132
rect 1536 1044 1558 1108
rect 1622 1044 1640 1108
rect 1536 1025 1640 1044
rect 2816 619 2920 1223
rect 2816 555 2837 619
rect 2901 555 2920 619
rect 2816 531 2920 555
rect 1550 -683 1654 -666
rect 1550 -747 1567 -683
rect 1631 -747 1654 -683
rect 1550 -982 1654 -747
rect 2830 -720 2934 -719
rect 2830 -822 2831 -720
rect 2933 -822 2934 -720
rect 2830 -953 2934 -822
use sky130_fd_pr__cap_mim_m3_1_3DGTNZ  sky130_fd_pr__cap_mim_m3_1_3DGTNZ_0
timestamp 1692509756
transform 1 0 1748 0 1 -3169
box -1186 -2320 1186 2320
use sky130_fd_pr__cap_mim_m3_1_3DGTNZ  sky130_fd_pr__cap_mim_m3_1_3DGTNZ_1
timestamp 1692509756
transform 1 0 1734 0 1 3421
box -1186 -2320 1186 2320
use sky130_fd_pr__cap_mim_m3_1_DMGF22  sky130_fd_pr__cap_mim_m3_1_DMGF22_0
timestamp 1692509756
transform 1 0 1888 0 1 2688
box 0 0 1 1
use sky130_fd_pr__nfet_g5v0d10v5_LWV9XU  sky130_fd_pr__nfet_g5v0d10v5_LWV9XU_0
timestamp 1692509756
transform 1 0 2251 0 1 -228
box -187 -157 187 157
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_0
timestamp 1692509756
transform 1 0 854 0 1 -259
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_1
timestamp 1692509756
transform 1 0 1895 0 1 -259
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_2
timestamp 1692509756
transform 1 0 1012 0 1 -259
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_3
timestamp 1692509756
transform 1 0 1737 0 1 -259
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_4
timestamp 1692509756
transform 1 0 1300 0 1 -259
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_5
timestamp 1692509756
transform 1 0 1579 0 1 -259
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_6
timestamp 1692509756
transform 1 0 2607 0 1 64
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_SACDK5  sky130_fd_pr__nfet_g5v0d10v5_SACDK5_7
timestamp 1692509756
transform 1 0 2330 0 1 55
box -108 -126 108 126
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_0
timestamp 1692509756
transform 1 0 1895 0 1 177
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_1
timestamp 1692509756
transform 1 0 1012 0 1 182
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7  sky130_fd_pr__pfet_g5v0d10v5_NQ4LZ7_2
timestamp 1692509756
transform 1 0 2206 0 1 463
box -174 -166 174 166
use sky130_fd_pr__pfet_g5v0d10v5_TUZSY8  sky130_fd_pr__pfet_g5v0d10v5_TUZSY8_0
timestamp 1692509756
transform 1 0 1595 0 1 514
box -253 -202 253 164
use sky130_fd_pr__pfet_g5v0d10v5_YM4LZ5  sky130_fd_pr__pfet_g5v0d10v5_YM4LZ5_0
timestamp 1692509756
transform -1 0 1012 0 -1 514
box -174 -164 174 202
use sky130_fd_pr__pfet_g5v0d10v5_YM4LZ5  sky130_fd_pr__pfet_g5v0d10v5_YM4LZ5_1
timestamp 1692509756
transform -1 0 1300 0 -1 184
box -174 -164 174 202
<< labels >>
flabel metal2 s 637 125 637 125 7 FreeSans 1600 0 0 0 CLK
flabel metal2 s 619 367 619 367 7 FreeSans 1600 0 0 0 VIN
flabel metal2 s 2924 -301 2924 -301 3 FreeSans 1600 0 0 0 VOUT
flabel metal3 s 520 874 520 874 7 FreeSans 1600 0 0 0 VCC
flabel metal3 s 649 -511 649 -511 7 FreeSans 1600 0 0 0 VSS
<< end >>
