magic
tech sky130A
magscale 1 2
timestamp 1687977505
<< nwell >>
rect 1280 19332 1946 19538
rect 3378 19520 4292 19528
rect 5622 19520 6250 19528
rect 3378 19332 4984 19520
rect 1280 19260 4984 19332
rect 1328 19008 4984 19260
rect 5622 19008 6942 19520
rect 1328 19000 3480 19008
rect 1328 18998 3408 19000
rect 2832 18994 3146 18998
rect 1280 18104 1946 18310
rect 3378 18292 4292 18300
rect 5622 18292 6250 18300
rect 3378 18104 4984 18292
rect 1280 18032 4984 18104
rect 1328 17780 4984 18032
rect 5622 17780 6942 18292
rect 1328 17772 3480 17780
rect 1328 17770 3408 17772
rect 2832 17766 3146 17770
rect 1280 16876 1946 17082
rect 3378 17064 4292 17072
rect 5622 17064 6250 17072
rect 3378 16876 4984 17064
rect 1280 16804 4984 16876
rect 1328 16552 4984 16804
rect 5622 16552 6942 17064
rect 1328 16544 3480 16552
rect 1328 16542 3408 16544
rect 2832 16538 3146 16542
rect 1280 15648 1946 15854
rect 3378 15836 4292 15844
rect 5622 15836 6250 15844
rect 3378 15648 4984 15836
rect 1280 15576 4984 15648
rect 1328 15324 4984 15576
rect 5622 15324 6942 15836
rect 1328 15316 3480 15324
rect 1328 15314 3408 15316
rect 2832 15310 3146 15314
rect 1280 14420 1946 14626
rect 3378 14608 4292 14616
rect 5622 14608 6250 14616
rect 3378 14420 4984 14608
rect 1280 14348 4984 14420
rect 1328 14096 4984 14348
rect 5622 14096 6942 14608
rect 1328 14088 3480 14096
rect 1328 14086 3408 14088
rect 2832 14082 3146 14086
rect 1280 13192 1946 13398
rect 3378 13380 4292 13388
rect 5622 13380 6250 13388
rect 3378 13192 4984 13380
rect 1280 13120 4984 13192
rect 1328 12868 4984 13120
rect 5622 12868 6942 13380
rect 1328 12860 3480 12868
rect 1328 12858 3408 12860
rect 2832 12854 3146 12858
rect 1280 11964 1946 12170
rect 3378 12152 4292 12160
rect 5622 12152 6250 12160
rect 3378 11964 4984 12152
rect 1280 11892 4984 11964
rect 1328 11640 4984 11892
rect 5622 11640 6942 12152
rect 1328 11632 3480 11640
rect 1328 11630 3408 11632
rect 2832 11626 3146 11630
rect 1280 10736 1946 10942
rect 3378 10924 4292 10932
rect 5622 10924 6250 10932
rect 3378 10736 4984 10924
rect 1280 10664 4984 10736
rect 1328 10412 4984 10664
rect 5622 10412 6942 10924
rect 1328 10404 3480 10412
rect 1328 10402 3408 10404
rect 2832 10398 3146 10402
rect 1280 9508 1946 9714
rect 3378 9696 4292 9704
rect 5622 9696 6250 9704
rect 3378 9508 4984 9696
rect 1280 9436 4984 9508
rect 1328 9184 4984 9436
rect 5622 9184 6942 9696
rect 1328 9176 3480 9184
rect 1328 9174 3408 9176
rect 2832 9170 3146 9174
rect 1280 8280 1946 8486
rect 3378 8468 4292 8476
rect 5622 8468 6250 8476
rect 3378 8280 4984 8468
rect 1280 8208 4984 8280
rect 1328 7956 4984 8208
rect 5622 7956 6942 8468
rect 1328 7948 3480 7956
rect 1328 7946 3408 7948
rect 2832 7942 3146 7946
rect 1280 7052 1946 7258
rect 3378 7240 4292 7248
rect 5622 7240 6250 7248
rect 3378 7052 4984 7240
rect 1280 6980 4984 7052
rect 1328 6728 4984 6980
rect 5622 6728 6942 7240
rect 1328 6720 3480 6728
rect 1328 6718 3408 6720
rect 2832 6714 3146 6718
rect 1280 5824 1946 6030
rect 3378 6012 4292 6020
rect 5622 6012 6250 6020
rect 3378 5824 4984 6012
rect 1280 5752 4984 5824
rect 1328 5500 4984 5752
rect 5622 5500 6942 6012
rect 1328 5492 3480 5500
rect 1328 5490 3408 5492
rect 2832 5486 3146 5490
rect 1280 4596 1946 4802
rect 3378 4784 4292 4792
rect 5622 4784 6250 4792
rect 3378 4596 4984 4784
rect 1280 4524 4984 4596
rect 1328 4272 4984 4524
rect 5622 4272 6942 4784
rect 1328 4264 3480 4272
rect 1328 4262 3408 4264
rect 2832 4258 3146 4262
rect 1280 3368 1946 3574
rect 3378 3556 4292 3564
rect 5622 3556 6250 3564
rect 3378 3368 4984 3556
rect 1280 3296 4984 3368
rect 1328 3044 4984 3296
rect 5622 3044 6942 3556
rect 1328 3036 3480 3044
rect 1328 3034 3408 3036
rect 2832 3030 3146 3034
rect 1280 2140 1946 2346
rect 3378 2328 4292 2336
rect 5622 2328 6250 2336
rect 3378 2140 4984 2328
rect 1280 2068 4984 2140
rect 1328 1816 4984 2068
rect 5622 1816 6942 2328
rect 1328 1808 3480 1816
rect 1328 1806 3408 1808
rect 2832 1802 3146 1806
rect 1280 912 1946 1118
rect 3378 1100 4292 1108
rect 3378 912 4984 1100
rect 1280 840 4984 912
rect 1328 588 4984 840
rect 1328 580 3480 588
rect 1328 578 3408 580
rect 2832 574 3146 578
<< pwell >>
rect 808 19386 1098 19392
rect 518 18714 1098 19386
rect 4364 18962 4940 18964
rect 6322 18962 6898 18964
rect 1372 18800 3350 18952
rect 3704 18812 4940 18962
rect 5662 18812 6898 18962
rect 3704 18810 4280 18812
rect 5662 18810 6238 18812
rect 3704 18806 4270 18810
rect 5662 18806 6228 18810
rect 1372 18794 1985 18800
rect 518 18708 800 18714
rect 1298 18614 1985 18794
rect 3678 18614 4270 18806
rect 5636 18614 6228 18806
rect 808 18158 1098 18164
rect 518 17486 1098 18158
rect 4364 17734 4940 17736
rect 6322 17734 6898 17736
rect 1372 17572 3350 17724
rect 3704 17584 4940 17734
rect 5662 17584 6898 17734
rect 3704 17582 4280 17584
rect 5662 17582 6238 17584
rect 3704 17578 4270 17582
rect 5662 17578 6228 17582
rect 1372 17566 1985 17572
rect 518 17480 800 17486
rect 1298 17386 1985 17566
rect 3678 17386 4270 17578
rect 5636 17386 6228 17578
rect 808 16930 1098 16936
rect 518 16258 1098 16930
rect 4364 16506 4940 16508
rect 6322 16506 6898 16508
rect 1372 16344 3350 16496
rect 3704 16356 4940 16506
rect 5662 16356 6898 16506
rect 3704 16354 4280 16356
rect 5662 16354 6238 16356
rect 3704 16350 4270 16354
rect 5662 16350 6228 16354
rect 1372 16338 1985 16344
rect 518 16252 800 16258
rect 1298 16158 1985 16338
rect 3678 16158 4270 16350
rect 5636 16158 6228 16350
rect 808 15702 1098 15708
rect 518 15030 1098 15702
rect 4364 15278 4940 15280
rect 6322 15278 6898 15280
rect 1372 15116 3350 15268
rect 3704 15128 4940 15278
rect 5662 15128 6898 15278
rect 3704 15126 4280 15128
rect 5662 15126 6238 15128
rect 3704 15122 4270 15126
rect 5662 15122 6228 15126
rect 1372 15110 1985 15116
rect 518 15024 800 15030
rect 1298 14930 1985 15110
rect 3678 14930 4270 15122
rect 5636 14930 6228 15122
rect 808 14474 1098 14480
rect 518 13802 1098 14474
rect 4364 14050 4940 14052
rect 6322 14050 6898 14052
rect 1372 13888 3350 14040
rect 3704 13900 4940 14050
rect 5662 13900 6898 14050
rect 3704 13898 4280 13900
rect 5662 13898 6238 13900
rect 3704 13894 4270 13898
rect 5662 13894 6228 13898
rect 1372 13882 1985 13888
rect 518 13796 800 13802
rect 1298 13702 1985 13882
rect 3678 13702 4270 13894
rect 5636 13702 6228 13894
rect 808 13246 1098 13252
rect 518 12574 1098 13246
rect 4364 12822 4940 12824
rect 6322 12822 6898 12824
rect 1372 12660 3350 12812
rect 3704 12672 4940 12822
rect 5662 12672 6898 12822
rect 3704 12670 4280 12672
rect 5662 12670 6238 12672
rect 3704 12666 4270 12670
rect 5662 12666 6228 12670
rect 1372 12654 1985 12660
rect 518 12568 800 12574
rect 1298 12474 1985 12654
rect 3678 12474 4270 12666
rect 5636 12474 6228 12666
rect 808 12018 1098 12024
rect 518 11346 1098 12018
rect 4364 11594 4940 11596
rect 6322 11594 6898 11596
rect 1372 11432 3350 11584
rect 3704 11444 4940 11594
rect 5662 11444 6898 11594
rect 3704 11442 4280 11444
rect 5662 11442 6238 11444
rect 3704 11438 4270 11442
rect 5662 11438 6228 11442
rect 1372 11426 1985 11432
rect 518 11340 800 11346
rect 1298 11246 1985 11426
rect 3678 11246 4270 11438
rect 5636 11246 6228 11438
rect 808 10790 1098 10796
rect 518 10118 1098 10790
rect 4364 10366 4940 10368
rect 6322 10366 6898 10368
rect 1372 10204 3350 10356
rect 3704 10216 4940 10366
rect 5662 10216 6898 10366
rect 3704 10214 4280 10216
rect 5662 10214 6238 10216
rect 3704 10210 4270 10214
rect 5662 10210 6228 10214
rect 1372 10198 1985 10204
rect 518 10112 800 10118
rect 1298 10018 1985 10198
rect 3678 10018 4270 10210
rect 5636 10018 6228 10210
rect 808 9562 1098 9568
rect 518 8890 1098 9562
rect 4364 9138 4940 9140
rect 6322 9138 6898 9140
rect 1372 8976 3350 9128
rect 3704 8988 4940 9138
rect 5662 8988 6898 9138
rect 3704 8986 4280 8988
rect 5662 8986 6238 8988
rect 3704 8982 4270 8986
rect 5662 8982 6228 8986
rect 1372 8970 1985 8976
rect 518 8884 800 8890
rect 1298 8790 1985 8970
rect 3678 8790 4270 8982
rect 5636 8790 6228 8982
rect 808 8334 1098 8340
rect 518 7662 1098 8334
rect 4364 7910 4940 7912
rect 6322 7910 6898 7912
rect 1372 7748 3350 7900
rect 3704 7760 4940 7910
rect 5662 7760 6898 7910
rect 3704 7758 4280 7760
rect 5662 7758 6238 7760
rect 3704 7754 4270 7758
rect 5662 7754 6228 7758
rect 1372 7742 1985 7748
rect 518 7656 800 7662
rect 1298 7562 1985 7742
rect 3678 7562 4270 7754
rect 5636 7562 6228 7754
rect 808 7106 1098 7112
rect 518 6434 1098 7106
rect 4364 6682 4940 6684
rect 6322 6682 6898 6684
rect 1372 6520 3350 6672
rect 3704 6532 4940 6682
rect 5662 6532 6898 6682
rect 3704 6530 4280 6532
rect 5662 6530 6238 6532
rect 3704 6526 4270 6530
rect 5662 6526 6228 6530
rect 1372 6514 1985 6520
rect 518 6428 800 6434
rect 1298 6334 1985 6514
rect 3678 6334 4270 6526
rect 5636 6334 6228 6526
rect 808 5878 1098 5884
rect 518 5206 1098 5878
rect 4364 5454 4940 5456
rect 6322 5454 6898 5456
rect 1372 5292 3350 5444
rect 3704 5304 4940 5454
rect 5662 5304 6898 5454
rect 3704 5302 4280 5304
rect 5662 5302 6238 5304
rect 3704 5298 4270 5302
rect 5662 5298 6228 5302
rect 1372 5286 1985 5292
rect 518 5200 800 5206
rect 1298 5106 1985 5286
rect 3678 5106 4270 5298
rect 5636 5106 6228 5298
rect 808 4650 1098 4656
rect 518 3978 1098 4650
rect 4364 4226 4940 4228
rect 6322 4226 6898 4228
rect 1372 4064 3350 4216
rect 3704 4076 4940 4226
rect 5662 4076 6898 4226
rect 3704 4074 4280 4076
rect 5662 4074 6238 4076
rect 3704 4070 4270 4074
rect 5662 4070 6228 4074
rect 1372 4058 1985 4064
rect 518 3972 800 3978
rect 1298 3878 1985 4058
rect 3678 3878 4270 4070
rect 5636 3878 6228 4070
rect 808 3422 1098 3428
rect 518 2750 1098 3422
rect 4364 2998 4940 3000
rect 6322 2998 6898 3000
rect 1372 2836 3350 2988
rect 3704 2848 4940 2998
rect 5662 2848 6898 2998
rect 3704 2846 4280 2848
rect 5662 2846 6238 2848
rect 3704 2842 4270 2846
rect 5662 2842 6228 2846
rect 1372 2830 1985 2836
rect 518 2744 800 2750
rect 1298 2650 1985 2830
rect 3678 2650 4270 2842
rect 5636 2650 6228 2842
rect 808 2194 1098 2200
rect 518 1522 1098 2194
rect 4364 1770 4940 1772
rect 6322 1770 6898 1772
rect 1372 1608 3350 1760
rect 3704 1620 4940 1770
rect 5662 1620 6898 1770
rect 3704 1618 4280 1620
rect 5662 1618 6238 1620
rect 3704 1614 4270 1618
rect 5662 1614 6228 1618
rect 1372 1602 1985 1608
rect 518 1516 800 1522
rect 1298 1422 1985 1602
rect 3678 1422 4270 1614
rect 5636 1422 6228 1614
rect 808 966 1098 972
rect 518 294 1098 966
rect 4364 542 4940 544
rect 1372 380 3350 532
rect 3704 392 4940 542
rect 3704 390 4280 392
rect 3704 386 4270 390
rect 1372 374 1985 380
rect 518 288 800 294
rect 1298 194 1985 374
rect 3678 194 4270 386
<< mvnmos >>
rect 1456 18826 1556 18926
rect 1744 18826 1844 18926
rect 2076 18826 2176 18926
rect 2418 18826 2518 18926
rect 2822 18826 2922 18926
rect 3166 18826 3266 18926
rect 3788 18836 3888 18936
rect 4096 18836 4196 18936
rect 4448 18838 4548 18938
rect 4756 18838 4856 18938
rect 5746 18836 5846 18936
rect 6054 18836 6154 18936
rect 6406 18838 6506 18938
rect 6714 18838 6814 18938
rect 1456 17598 1556 17698
rect 1744 17598 1844 17698
rect 2076 17598 2176 17698
rect 2418 17598 2518 17698
rect 2822 17598 2922 17698
rect 3166 17598 3266 17698
rect 3788 17608 3888 17708
rect 4096 17608 4196 17708
rect 4448 17610 4548 17710
rect 4756 17610 4856 17710
rect 5746 17608 5846 17708
rect 6054 17608 6154 17708
rect 6406 17610 6506 17710
rect 6714 17610 6814 17710
rect 1456 16370 1556 16470
rect 1744 16370 1844 16470
rect 2076 16370 2176 16470
rect 2418 16370 2518 16470
rect 2822 16370 2922 16470
rect 3166 16370 3266 16470
rect 3788 16380 3888 16480
rect 4096 16380 4196 16480
rect 4448 16382 4548 16482
rect 4756 16382 4856 16482
rect 5746 16380 5846 16480
rect 6054 16380 6154 16480
rect 6406 16382 6506 16482
rect 6714 16382 6814 16482
rect 1456 15142 1556 15242
rect 1744 15142 1844 15242
rect 2076 15142 2176 15242
rect 2418 15142 2518 15242
rect 2822 15142 2922 15242
rect 3166 15142 3266 15242
rect 3788 15152 3888 15252
rect 4096 15152 4196 15252
rect 4448 15154 4548 15254
rect 4756 15154 4856 15254
rect 5746 15152 5846 15252
rect 6054 15152 6154 15252
rect 6406 15154 6506 15254
rect 6714 15154 6814 15254
rect 1456 13914 1556 14014
rect 1744 13914 1844 14014
rect 2076 13914 2176 14014
rect 2418 13914 2518 14014
rect 2822 13914 2922 14014
rect 3166 13914 3266 14014
rect 3788 13924 3888 14024
rect 4096 13924 4196 14024
rect 4448 13926 4548 14026
rect 4756 13926 4856 14026
rect 5746 13924 5846 14024
rect 6054 13924 6154 14024
rect 6406 13926 6506 14026
rect 6714 13926 6814 14026
rect 1456 12686 1556 12786
rect 1744 12686 1844 12786
rect 2076 12686 2176 12786
rect 2418 12686 2518 12786
rect 2822 12686 2922 12786
rect 3166 12686 3266 12786
rect 3788 12696 3888 12796
rect 4096 12696 4196 12796
rect 4448 12698 4548 12798
rect 4756 12698 4856 12798
rect 5746 12696 5846 12796
rect 6054 12696 6154 12796
rect 6406 12698 6506 12798
rect 6714 12698 6814 12798
rect 1456 11458 1556 11558
rect 1744 11458 1844 11558
rect 2076 11458 2176 11558
rect 2418 11458 2518 11558
rect 2822 11458 2922 11558
rect 3166 11458 3266 11558
rect 3788 11468 3888 11568
rect 4096 11468 4196 11568
rect 4448 11470 4548 11570
rect 4756 11470 4856 11570
rect 5746 11468 5846 11568
rect 6054 11468 6154 11568
rect 6406 11470 6506 11570
rect 6714 11470 6814 11570
rect 1456 10230 1556 10330
rect 1744 10230 1844 10330
rect 2076 10230 2176 10330
rect 2418 10230 2518 10330
rect 2822 10230 2922 10330
rect 3166 10230 3266 10330
rect 3788 10240 3888 10340
rect 4096 10240 4196 10340
rect 4448 10242 4548 10342
rect 4756 10242 4856 10342
rect 5746 10240 5846 10340
rect 6054 10240 6154 10340
rect 6406 10242 6506 10342
rect 6714 10242 6814 10342
rect 1456 9002 1556 9102
rect 1744 9002 1844 9102
rect 2076 9002 2176 9102
rect 2418 9002 2518 9102
rect 2822 9002 2922 9102
rect 3166 9002 3266 9102
rect 3788 9012 3888 9112
rect 4096 9012 4196 9112
rect 4448 9014 4548 9114
rect 4756 9014 4856 9114
rect 5746 9012 5846 9112
rect 6054 9012 6154 9112
rect 6406 9014 6506 9114
rect 6714 9014 6814 9114
rect 1456 7774 1556 7874
rect 1744 7774 1844 7874
rect 2076 7774 2176 7874
rect 2418 7774 2518 7874
rect 2822 7774 2922 7874
rect 3166 7774 3266 7874
rect 3788 7784 3888 7884
rect 4096 7784 4196 7884
rect 4448 7786 4548 7886
rect 4756 7786 4856 7886
rect 5746 7784 5846 7884
rect 6054 7784 6154 7884
rect 6406 7786 6506 7886
rect 6714 7786 6814 7886
rect 1456 6546 1556 6646
rect 1744 6546 1844 6646
rect 2076 6546 2176 6646
rect 2418 6546 2518 6646
rect 2822 6546 2922 6646
rect 3166 6546 3266 6646
rect 3788 6556 3888 6656
rect 4096 6556 4196 6656
rect 4448 6558 4548 6658
rect 4756 6558 4856 6658
rect 5746 6556 5846 6656
rect 6054 6556 6154 6656
rect 6406 6558 6506 6658
rect 6714 6558 6814 6658
rect 1456 5318 1556 5418
rect 1744 5318 1844 5418
rect 2076 5318 2176 5418
rect 2418 5318 2518 5418
rect 2822 5318 2922 5418
rect 3166 5318 3266 5418
rect 3788 5328 3888 5428
rect 4096 5328 4196 5428
rect 4448 5330 4548 5430
rect 4756 5330 4856 5430
rect 5746 5328 5846 5428
rect 6054 5328 6154 5428
rect 6406 5330 6506 5430
rect 6714 5330 6814 5430
rect 1456 4090 1556 4190
rect 1744 4090 1844 4190
rect 2076 4090 2176 4190
rect 2418 4090 2518 4190
rect 2822 4090 2922 4190
rect 3166 4090 3266 4190
rect 3788 4100 3888 4200
rect 4096 4100 4196 4200
rect 4448 4102 4548 4202
rect 4756 4102 4856 4202
rect 5746 4100 5846 4200
rect 6054 4100 6154 4200
rect 6406 4102 6506 4202
rect 6714 4102 6814 4202
rect 1456 2862 1556 2962
rect 1744 2862 1844 2962
rect 2076 2862 2176 2962
rect 2418 2862 2518 2962
rect 2822 2862 2922 2962
rect 3166 2862 3266 2962
rect 3788 2872 3888 2972
rect 4096 2872 4196 2972
rect 4448 2874 4548 2974
rect 4756 2874 4856 2974
rect 5746 2872 5846 2972
rect 6054 2872 6154 2972
rect 6406 2874 6506 2974
rect 6714 2874 6814 2974
rect 1456 1634 1556 1734
rect 1744 1634 1844 1734
rect 2076 1634 2176 1734
rect 2418 1634 2518 1734
rect 2822 1634 2922 1734
rect 3166 1634 3266 1734
rect 3788 1644 3888 1744
rect 4096 1644 4196 1744
rect 4448 1646 4548 1746
rect 4756 1646 4856 1746
rect 5746 1644 5846 1744
rect 6054 1644 6154 1744
rect 6406 1646 6506 1746
rect 6714 1646 6814 1746
rect 1456 406 1556 506
rect 1744 406 1844 506
rect 2076 406 2176 506
rect 2418 406 2518 506
rect 2822 406 2922 506
rect 3166 406 3266 506
rect 3788 416 3888 516
rect 4096 416 4196 516
rect 4448 418 4548 518
rect 4756 418 4856 518
<< mvpmos >>
rect 1456 19064 1556 19264
rect 1744 19064 1844 19264
rect 2076 19064 2176 19264
rect 2418 19064 2518 19264
rect 2822 19064 2922 19264
rect 3166 19064 3266 19264
rect 3788 19074 3888 19274
rect 4096 19074 4196 19274
rect 4448 19074 4548 19274
rect 4756 19074 4856 19274
rect 5746 19074 5846 19274
rect 6054 19074 6154 19274
rect 6406 19074 6506 19274
rect 6714 19074 6814 19274
rect 1456 17836 1556 18036
rect 1744 17836 1844 18036
rect 2076 17836 2176 18036
rect 2418 17836 2518 18036
rect 2822 17836 2922 18036
rect 3166 17836 3266 18036
rect 3788 17846 3888 18046
rect 4096 17846 4196 18046
rect 4448 17846 4548 18046
rect 4756 17846 4856 18046
rect 5746 17846 5846 18046
rect 6054 17846 6154 18046
rect 6406 17846 6506 18046
rect 6714 17846 6814 18046
rect 1456 16608 1556 16808
rect 1744 16608 1844 16808
rect 2076 16608 2176 16808
rect 2418 16608 2518 16808
rect 2822 16608 2922 16808
rect 3166 16608 3266 16808
rect 3788 16618 3888 16818
rect 4096 16618 4196 16818
rect 4448 16618 4548 16818
rect 4756 16618 4856 16818
rect 5746 16618 5846 16818
rect 6054 16618 6154 16818
rect 6406 16618 6506 16818
rect 6714 16618 6814 16818
rect 1456 15380 1556 15580
rect 1744 15380 1844 15580
rect 2076 15380 2176 15580
rect 2418 15380 2518 15580
rect 2822 15380 2922 15580
rect 3166 15380 3266 15580
rect 3788 15390 3888 15590
rect 4096 15390 4196 15590
rect 4448 15390 4548 15590
rect 4756 15390 4856 15590
rect 5746 15390 5846 15590
rect 6054 15390 6154 15590
rect 6406 15390 6506 15590
rect 6714 15390 6814 15590
rect 1456 14152 1556 14352
rect 1744 14152 1844 14352
rect 2076 14152 2176 14352
rect 2418 14152 2518 14352
rect 2822 14152 2922 14352
rect 3166 14152 3266 14352
rect 3788 14162 3888 14362
rect 4096 14162 4196 14362
rect 4448 14162 4548 14362
rect 4756 14162 4856 14362
rect 5746 14162 5846 14362
rect 6054 14162 6154 14362
rect 6406 14162 6506 14362
rect 6714 14162 6814 14362
rect 1456 12924 1556 13124
rect 1744 12924 1844 13124
rect 2076 12924 2176 13124
rect 2418 12924 2518 13124
rect 2822 12924 2922 13124
rect 3166 12924 3266 13124
rect 3788 12934 3888 13134
rect 4096 12934 4196 13134
rect 4448 12934 4548 13134
rect 4756 12934 4856 13134
rect 5746 12934 5846 13134
rect 6054 12934 6154 13134
rect 6406 12934 6506 13134
rect 6714 12934 6814 13134
rect 1456 11696 1556 11896
rect 1744 11696 1844 11896
rect 2076 11696 2176 11896
rect 2418 11696 2518 11896
rect 2822 11696 2922 11896
rect 3166 11696 3266 11896
rect 3788 11706 3888 11906
rect 4096 11706 4196 11906
rect 4448 11706 4548 11906
rect 4756 11706 4856 11906
rect 5746 11706 5846 11906
rect 6054 11706 6154 11906
rect 6406 11706 6506 11906
rect 6714 11706 6814 11906
rect 1456 10468 1556 10668
rect 1744 10468 1844 10668
rect 2076 10468 2176 10668
rect 2418 10468 2518 10668
rect 2822 10468 2922 10668
rect 3166 10468 3266 10668
rect 3788 10478 3888 10678
rect 4096 10478 4196 10678
rect 4448 10478 4548 10678
rect 4756 10478 4856 10678
rect 5746 10478 5846 10678
rect 6054 10478 6154 10678
rect 6406 10478 6506 10678
rect 6714 10478 6814 10678
rect 1456 9240 1556 9440
rect 1744 9240 1844 9440
rect 2076 9240 2176 9440
rect 2418 9240 2518 9440
rect 2822 9240 2922 9440
rect 3166 9240 3266 9440
rect 3788 9250 3888 9450
rect 4096 9250 4196 9450
rect 4448 9250 4548 9450
rect 4756 9250 4856 9450
rect 5746 9250 5846 9450
rect 6054 9250 6154 9450
rect 6406 9250 6506 9450
rect 6714 9250 6814 9450
rect 1456 8012 1556 8212
rect 1744 8012 1844 8212
rect 2076 8012 2176 8212
rect 2418 8012 2518 8212
rect 2822 8012 2922 8212
rect 3166 8012 3266 8212
rect 3788 8022 3888 8222
rect 4096 8022 4196 8222
rect 4448 8022 4548 8222
rect 4756 8022 4856 8222
rect 5746 8022 5846 8222
rect 6054 8022 6154 8222
rect 6406 8022 6506 8222
rect 6714 8022 6814 8222
rect 1456 6784 1556 6984
rect 1744 6784 1844 6984
rect 2076 6784 2176 6984
rect 2418 6784 2518 6984
rect 2822 6784 2922 6984
rect 3166 6784 3266 6984
rect 3788 6794 3888 6994
rect 4096 6794 4196 6994
rect 4448 6794 4548 6994
rect 4756 6794 4856 6994
rect 5746 6794 5846 6994
rect 6054 6794 6154 6994
rect 6406 6794 6506 6994
rect 6714 6794 6814 6994
rect 1456 5556 1556 5756
rect 1744 5556 1844 5756
rect 2076 5556 2176 5756
rect 2418 5556 2518 5756
rect 2822 5556 2922 5756
rect 3166 5556 3266 5756
rect 3788 5566 3888 5766
rect 4096 5566 4196 5766
rect 4448 5566 4548 5766
rect 4756 5566 4856 5766
rect 5746 5566 5846 5766
rect 6054 5566 6154 5766
rect 6406 5566 6506 5766
rect 6714 5566 6814 5766
rect 1456 4328 1556 4528
rect 1744 4328 1844 4528
rect 2076 4328 2176 4528
rect 2418 4328 2518 4528
rect 2822 4328 2922 4528
rect 3166 4328 3266 4528
rect 3788 4338 3888 4538
rect 4096 4338 4196 4538
rect 4448 4338 4548 4538
rect 4756 4338 4856 4538
rect 5746 4338 5846 4538
rect 6054 4338 6154 4538
rect 6406 4338 6506 4538
rect 6714 4338 6814 4538
rect 1456 3100 1556 3300
rect 1744 3100 1844 3300
rect 2076 3100 2176 3300
rect 2418 3100 2518 3300
rect 2822 3100 2922 3300
rect 3166 3100 3266 3300
rect 3788 3110 3888 3310
rect 4096 3110 4196 3310
rect 4448 3110 4548 3310
rect 4756 3110 4856 3310
rect 5746 3110 5846 3310
rect 6054 3110 6154 3310
rect 6406 3110 6506 3310
rect 6714 3110 6814 3310
rect 1456 1872 1556 2072
rect 1744 1872 1844 2072
rect 2076 1872 2176 2072
rect 2418 1872 2518 2072
rect 2822 1872 2922 2072
rect 3166 1872 3266 2072
rect 3788 1882 3888 2082
rect 4096 1882 4196 2082
rect 4448 1882 4548 2082
rect 4756 1882 4856 2082
rect 5746 1882 5846 2082
rect 6054 1882 6154 2082
rect 6406 1882 6506 2082
rect 6714 1882 6814 2082
rect 1456 644 1556 844
rect 1744 644 1844 844
rect 2076 644 2176 844
rect 2418 644 2518 844
rect 2822 644 2922 844
rect 3166 644 3266 844
rect 3788 654 3888 854
rect 4096 654 4196 854
rect 4448 654 4548 854
rect 4756 654 4856 854
<< mvndiff >>
rect 544 19348 628 19360
rect 544 19314 569 19348
rect 603 19314 628 19348
rect 544 19257 628 19314
rect 544 18780 628 18837
rect 544 18746 569 18780
rect 603 18746 628 18780
rect 544 18734 628 18746
rect 690 19348 774 19360
rect 690 19314 715 19348
rect 749 19314 774 19348
rect 690 19257 774 19314
rect 690 18780 774 18837
rect 690 18746 715 18780
rect 749 18746 774 18780
rect 690 18734 774 18746
rect 834 19354 918 19366
rect 834 19320 859 19354
rect 893 19320 918 19354
rect 834 19263 918 19320
rect 834 18786 918 18843
rect 834 18752 859 18786
rect 893 18752 918 18786
rect 834 18740 918 18752
rect 988 19354 1072 19366
rect 988 19320 1013 19354
rect 1047 19320 1072 19354
rect 988 19263 1072 19320
rect 988 18786 1072 18843
rect 1398 18893 1456 18926
rect 1398 18859 1410 18893
rect 1444 18859 1456 18893
rect 1398 18826 1456 18859
rect 1556 18893 1614 18926
rect 1556 18859 1568 18893
rect 1602 18859 1614 18893
rect 1556 18826 1614 18859
rect 1686 18893 1744 18926
rect 1686 18859 1698 18893
rect 1732 18859 1744 18893
rect 1686 18826 1744 18859
rect 1844 18893 1902 18926
rect 1844 18859 1856 18893
rect 1890 18859 1902 18893
rect 1844 18826 1902 18859
rect 2018 18893 2076 18926
rect 2018 18859 2030 18893
rect 2064 18859 2076 18893
rect 2018 18826 2076 18859
rect 2176 18893 2234 18926
rect 2176 18859 2188 18893
rect 2222 18859 2234 18893
rect 2176 18826 2234 18859
rect 2360 18893 2418 18926
rect 2360 18859 2372 18893
rect 2406 18859 2418 18893
rect 2360 18826 2418 18859
rect 2518 18893 2576 18926
rect 2518 18859 2530 18893
rect 2564 18859 2576 18893
rect 2518 18826 2576 18859
rect 2764 18893 2822 18926
rect 2764 18859 2776 18893
rect 2810 18859 2822 18893
rect 2764 18826 2822 18859
rect 2922 18893 2980 18926
rect 2922 18859 2934 18893
rect 2968 18859 2980 18893
rect 2922 18826 2980 18859
rect 3108 18893 3166 18926
rect 3108 18859 3120 18893
rect 3154 18859 3166 18893
rect 3108 18826 3166 18859
rect 3266 18893 3324 18926
rect 3266 18859 3278 18893
rect 3312 18859 3324 18893
rect 3266 18826 3324 18859
rect 3730 18903 3788 18936
rect 3730 18869 3742 18903
rect 3776 18869 3788 18903
rect 3730 18836 3788 18869
rect 3888 18903 3946 18936
rect 3888 18869 3900 18903
rect 3934 18869 3946 18903
rect 3888 18836 3946 18869
rect 4038 18903 4096 18936
rect 4038 18869 4050 18903
rect 4084 18869 4096 18903
rect 4038 18836 4096 18869
rect 4196 18903 4254 18936
rect 4196 18869 4208 18903
rect 4242 18869 4254 18903
rect 4196 18836 4254 18869
rect 4390 18905 4448 18938
rect 4390 18871 4402 18905
rect 4436 18871 4448 18905
rect 4390 18838 4448 18871
rect 4548 18905 4606 18938
rect 4548 18871 4560 18905
rect 4594 18871 4606 18905
rect 4548 18838 4606 18871
rect 4698 18905 4756 18938
rect 4698 18871 4710 18905
rect 4744 18871 4756 18905
rect 4698 18838 4756 18871
rect 4856 18905 4914 18938
rect 4856 18871 4868 18905
rect 4902 18871 4914 18905
rect 4856 18838 4914 18871
rect 5688 18904 5746 18936
rect 5688 18870 5700 18904
rect 5734 18870 5746 18904
rect 5688 18836 5746 18870
rect 5846 18904 5904 18936
rect 5846 18870 5858 18904
rect 5892 18870 5904 18904
rect 5846 18836 5904 18870
rect 5996 18904 6054 18936
rect 5996 18870 6008 18904
rect 6042 18870 6054 18904
rect 5996 18836 6054 18870
rect 6154 18904 6212 18936
rect 6154 18870 6166 18904
rect 6200 18870 6212 18904
rect 6154 18836 6212 18870
rect 6348 18906 6406 18938
rect 6348 18872 6360 18906
rect 6394 18872 6406 18906
rect 6348 18838 6406 18872
rect 6506 18906 6564 18938
rect 6506 18872 6518 18906
rect 6552 18872 6564 18906
rect 6506 18838 6564 18872
rect 6656 18906 6714 18938
rect 6656 18872 6668 18906
rect 6702 18872 6714 18906
rect 6656 18838 6714 18872
rect 6814 18906 6872 18938
rect 6814 18872 6826 18906
rect 6860 18872 6872 18906
rect 6814 18838 6872 18872
rect 988 18752 1013 18786
rect 1047 18752 1072 18786
rect 988 18740 1072 18752
rect 544 18120 628 18132
rect 544 18086 569 18120
rect 603 18086 628 18120
rect 544 18029 628 18086
rect 544 17552 628 17609
rect 544 17518 569 17552
rect 603 17518 628 17552
rect 544 17506 628 17518
rect 690 18120 774 18132
rect 690 18086 715 18120
rect 749 18086 774 18120
rect 690 18029 774 18086
rect 690 17552 774 17609
rect 690 17518 715 17552
rect 749 17518 774 17552
rect 690 17506 774 17518
rect 834 18126 918 18138
rect 834 18092 859 18126
rect 893 18092 918 18126
rect 834 18035 918 18092
rect 834 17558 918 17615
rect 834 17524 859 17558
rect 893 17524 918 17558
rect 834 17512 918 17524
rect 988 18126 1072 18138
rect 988 18092 1013 18126
rect 1047 18092 1072 18126
rect 988 18035 1072 18092
rect 988 17558 1072 17615
rect 1398 17665 1456 17698
rect 1398 17631 1410 17665
rect 1444 17631 1456 17665
rect 1398 17598 1456 17631
rect 1556 17665 1614 17698
rect 1556 17631 1568 17665
rect 1602 17631 1614 17665
rect 1556 17598 1614 17631
rect 1686 17665 1744 17698
rect 1686 17631 1698 17665
rect 1732 17631 1744 17665
rect 1686 17598 1744 17631
rect 1844 17665 1902 17698
rect 1844 17631 1856 17665
rect 1890 17631 1902 17665
rect 1844 17598 1902 17631
rect 2018 17665 2076 17698
rect 2018 17631 2030 17665
rect 2064 17631 2076 17665
rect 2018 17598 2076 17631
rect 2176 17665 2234 17698
rect 2176 17631 2188 17665
rect 2222 17631 2234 17665
rect 2176 17598 2234 17631
rect 2360 17665 2418 17698
rect 2360 17631 2372 17665
rect 2406 17631 2418 17665
rect 2360 17598 2418 17631
rect 2518 17665 2576 17698
rect 2518 17631 2530 17665
rect 2564 17631 2576 17665
rect 2518 17598 2576 17631
rect 2764 17665 2822 17698
rect 2764 17631 2776 17665
rect 2810 17631 2822 17665
rect 2764 17598 2822 17631
rect 2922 17665 2980 17698
rect 2922 17631 2934 17665
rect 2968 17631 2980 17665
rect 2922 17598 2980 17631
rect 3108 17665 3166 17698
rect 3108 17631 3120 17665
rect 3154 17631 3166 17665
rect 3108 17598 3166 17631
rect 3266 17665 3324 17698
rect 3266 17631 3278 17665
rect 3312 17631 3324 17665
rect 3266 17598 3324 17631
rect 3730 17675 3788 17708
rect 3730 17641 3742 17675
rect 3776 17641 3788 17675
rect 3730 17608 3788 17641
rect 3888 17675 3946 17708
rect 3888 17641 3900 17675
rect 3934 17641 3946 17675
rect 3888 17608 3946 17641
rect 4038 17675 4096 17708
rect 4038 17641 4050 17675
rect 4084 17641 4096 17675
rect 4038 17608 4096 17641
rect 4196 17675 4254 17708
rect 4196 17641 4208 17675
rect 4242 17641 4254 17675
rect 4196 17608 4254 17641
rect 4390 17677 4448 17710
rect 4390 17643 4402 17677
rect 4436 17643 4448 17677
rect 4390 17610 4448 17643
rect 4548 17677 4606 17710
rect 4548 17643 4560 17677
rect 4594 17643 4606 17677
rect 4548 17610 4606 17643
rect 4698 17677 4756 17710
rect 4698 17643 4710 17677
rect 4744 17643 4756 17677
rect 4698 17610 4756 17643
rect 4856 17677 4914 17710
rect 4856 17643 4868 17677
rect 4902 17643 4914 17677
rect 4856 17610 4914 17643
rect 5688 17676 5746 17708
rect 5688 17642 5700 17676
rect 5734 17642 5746 17676
rect 5688 17608 5746 17642
rect 5846 17676 5904 17708
rect 5846 17642 5858 17676
rect 5892 17642 5904 17676
rect 5846 17608 5904 17642
rect 5996 17676 6054 17708
rect 5996 17642 6008 17676
rect 6042 17642 6054 17676
rect 5996 17608 6054 17642
rect 6154 17676 6212 17708
rect 6154 17642 6166 17676
rect 6200 17642 6212 17676
rect 6154 17608 6212 17642
rect 6348 17678 6406 17710
rect 6348 17644 6360 17678
rect 6394 17644 6406 17678
rect 6348 17610 6406 17644
rect 6506 17678 6564 17710
rect 6506 17644 6518 17678
rect 6552 17644 6564 17678
rect 6506 17610 6564 17644
rect 6656 17678 6714 17710
rect 6656 17644 6668 17678
rect 6702 17644 6714 17678
rect 6656 17610 6714 17644
rect 6814 17678 6872 17710
rect 6814 17644 6826 17678
rect 6860 17644 6872 17678
rect 6814 17610 6872 17644
rect 988 17524 1013 17558
rect 1047 17524 1072 17558
rect 988 17512 1072 17524
rect 544 16892 628 16904
rect 544 16858 569 16892
rect 603 16858 628 16892
rect 544 16801 628 16858
rect 544 16324 628 16381
rect 544 16290 569 16324
rect 603 16290 628 16324
rect 544 16278 628 16290
rect 690 16892 774 16904
rect 690 16858 715 16892
rect 749 16858 774 16892
rect 690 16801 774 16858
rect 690 16324 774 16381
rect 690 16290 715 16324
rect 749 16290 774 16324
rect 690 16278 774 16290
rect 834 16898 918 16910
rect 834 16864 859 16898
rect 893 16864 918 16898
rect 834 16807 918 16864
rect 834 16330 918 16387
rect 834 16296 859 16330
rect 893 16296 918 16330
rect 834 16284 918 16296
rect 988 16898 1072 16910
rect 988 16864 1013 16898
rect 1047 16864 1072 16898
rect 988 16807 1072 16864
rect 988 16330 1072 16387
rect 1398 16437 1456 16470
rect 1398 16403 1410 16437
rect 1444 16403 1456 16437
rect 1398 16370 1456 16403
rect 1556 16437 1614 16470
rect 1556 16403 1568 16437
rect 1602 16403 1614 16437
rect 1556 16370 1614 16403
rect 1686 16437 1744 16470
rect 1686 16403 1698 16437
rect 1732 16403 1744 16437
rect 1686 16370 1744 16403
rect 1844 16437 1902 16470
rect 1844 16403 1856 16437
rect 1890 16403 1902 16437
rect 1844 16370 1902 16403
rect 2018 16437 2076 16470
rect 2018 16403 2030 16437
rect 2064 16403 2076 16437
rect 2018 16370 2076 16403
rect 2176 16437 2234 16470
rect 2176 16403 2188 16437
rect 2222 16403 2234 16437
rect 2176 16370 2234 16403
rect 2360 16437 2418 16470
rect 2360 16403 2372 16437
rect 2406 16403 2418 16437
rect 2360 16370 2418 16403
rect 2518 16437 2576 16470
rect 2518 16403 2530 16437
rect 2564 16403 2576 16437
rect 2518 16370 2576 16403
rect 2764 16437 2822 16470
rect 2764 16403 2776 16437
rect 2810 16403 2822 16437
rect 2764 16370 2822 16403
rect 2922 16437 2980 16470
rect 2922 16403 2934 16437
rect 2968 16403 2980 16437
rect 2922 16370 2980 16403
rect 3108 16437 3166 16470
rect 3108 16403 3120 16437
rect 3154 16403 3166 16437
rect 3108 16370 3166 16403
rect 3266 16437 3324 16470
rect 3266 16403 3278 16437
rect 3312 16403 3324 16437
rect 3266 16370 3324 16403
rect 3730 16447 3788 16480
rect 3730 16413 3742 16447
rect 3776 16413 3788 16447
rect 3730 16380 3788 16413
rect 3888 16447 3946 16480
rect 3888 16413 3900 16447
rect 3934 16413 3946 16447
rect 3888 16380 3946 16413
rect 4038 16447 4096 16480
rect 4038 16413 4050 16447
rect 4084 16413 4096 16447
rect 4038 16380 4096 16413
rect 4196 16447 4254 16480
rect 4196 16413 4208 16447
rect 4242 16413 4254 16447
rect 4196 16380 4254 16413
rect 4390 16449 4448 16482
rect 4390 16415 4402 16449
rect 4436 16415 4448 16449
rect 4390 16382 4448 16415
rect 4548 16449 4606 16482
rect 4548 16415 4560 16449
rect 4594 16415 4606 16449
rect 4548 16382 4606 16415
rect 4698 16449 4756 16482
rect 4698 16415 4710 16449
rect 4744 16415 4756 16449
rect 4698 16382 4756 16415
rect 4856 16449 4914 16482
rect 4856 16415 4868 16449
rect 4902 16415 4914 16449
rect 4856 16382 4914 16415
rect 5688 16448 5746 16480
rect 5688 16414 5700 16448
rect 5734 16414 5746 16448
rect 5688 16380 5746 16414
rect 5846 16448 5904 16480
rect 5846 16414 5858 16448
rect 5892 16414 5904 16448
rect 5846 16380 5904 16414
rect 5996 16448 6054 16480
rect 5996 16414 6008 16448
rect 6042 16414 6054 16448
rect 5996 16380 6054 16414
rect 6154 16448 6212 16480
rect 6154 16414 6166 16448
rect 6200 16414 6212 16448
rect 6154 16380 6212 16414
rect 6348 16450 6406 16482
rect 6348 16416 6360 16450
rect 6394 16416 6406 16450
rect 6348 16382 6406 16416
rect 6506 16450 6564 16482
rect 6506 16416 6518 16450
rect 6552 16416 6564 16450
rect 6506 16382 6564 16416
rect 6656 16450 6714 16482
rect 6656 16416 6668 16450
rect 6702 16416 6714 16450
rect 6656 16382 6714 16416
rect 6814 16450 6872 16482
rect 6814 16416 6826 16450
rect 6860 16416 6872 16450
rect 6814 16382 6872 16416
rect 988 16296 1013 16330
rect 1047 16296 1072 16330
rect 988 16284 1072 16296
rect 544 15664 628 15676
rect 544 15630 569 15664
rect 603 15630 628 15664
rect 544 15573 628 15630
rect 544 15096 628 15153
rect 544 15062 569 15096
rect 603 15062 628 15096
rect 544 15050 628 15062
rect 690 15664 774 15676
rect 690 15630 715 15664
rect 749 15630 774 15664
rect 690 15573 774 15630
rect 690 15096 774 15153
rect 690 15062 715 15096
rect 749 15062 774 15096
rect 690 15050 774 15062
rect 834 15670 918 15682
rect 834 15636 859 15670
rect 893 15636 918 15670
rect 834 15579 918 15636
rect 834 15102 918 15159
rect 834 15068 859 15102
rect 893 15068 918 15102
rect 834 15056 918 15068
rect 988 15670 1072 15682
rect 988 15636 1013 15670
rect 1047 15636 1072 15670
rect 988 15579 1072 15636
rect 988 15102 1072 15159
rect 1398 15209 1456 15242
rect 1398 15175 1410 15209
rect 1444 15175 1456 15209
rect 1398 15142 1456 15175
rect 1556 15209 1614 15242
rect 1556 15175 1568 15209
rect 1602 15175 1614 15209
rect 1556 15142 1614 15175
rect 1686 15209 1744 15242
rect 1686 15175 1698 15209
rect 1732 15175 1744 15209
rect 1686 15142 1744 15175
rect 1844 15209 1902 15242
rect 1844 15175 1856 15209
rect 1890 15175 1902 15209
rect 1844 15142 1902 15175
rect 2018 15209 2076 15242
rect 2018 15175 2030 15209
rect 2064 15175 2076 15209
rect 2018 15142 2076 15175
rect 2176 15209 2234 15242
rect 2176 15175 2188 15209
rect 2222 15175 2234 15209
rect 2176 15142 2234 15175
rect 2360 15209 2418 15242
rect 2360 15175 2372 15209
rect 2406 15175 2418 15209
rect 2360 15142 2418 15175
rect 2518 15209 2576 15242
rect 2518 15175 2530 15209
rect 2564 15175 2576 15209
rect 2518 15142 2576 15175
rect 2764 15209 2822 15242
rect 2764 15175 2776 15209
rect 2810 15175 2822 15209
rect 2764 15142 2822 15175
rect 2922 15209 2980 15242
rect 2922 15175 2934 15209
rect 2968 15175 2980 15209
rect 2922 15142 2980 15175
rect 3108 15209 3166 15242
rect 3108 15175 3120 15209
rect 3154 15175 3166 15209
rect 3108 15142 3166 15175
rect 3266 15209 3324 15242
rect 3266 15175 3278 15209
rect 3312 15175 3324 15209
rect 3266 15142 3324 15175
rect 3730 15219 3788 15252
rect 3730 15185 3742 15219
rect 3776 15185 3788 15219
rect 3730 15152 3788 15185
rect 3888 15219 3946 15252
rect 3888 15185 3900 15219
rect 3934 15185 3946 15219
rect 3888 15152 3946 15185
rect 4038 15219 4096 15252
rect 4038 15185 4050 15219
rect 4084 15185 4096 15219
rect 4038 15152 4096 15185
rect 4196 15219 4254 15252
rect 4196 15185 4208 15219
rect 4242 15185 4254 15219
rect 4196 15152 4254 15185
rect 4390 15221 4448 15254
rect 4390 15187 4402 15221
rect 4436 15187 4448 15221
rect 4390 15154 4448 15187
rect 4548 15221 4606 15254
rect 4548 15187 4560 15221
rect 4594 15187 4606 15221
rect 4548 15154 4606 15187
rect 4698 15221 4756 15254
rect 4698 15187 4710 15221
rect 4744 15187 4756 15221
rect 4698 15154 4756 15187
rect 4856 15221 4914 15254
rect 4856 15187 4868 15221
rect 4902 15187 4914 15221
rect 4856 15154 4914 15187
rect 5688 15220 5746 15252
rect 5688 15186 5700 15220
rect 5734 15186 5746 15220
rect 5688 15152 5746 15186
rect 5846 15220 5904 15252
rect 5846 15186 5858 15220
rect 5892 15186 5904 15220
rect 5846 15152 5904 15186
rect 5996 15220 6054 15252
rect 5996 15186 6008 15220
rect 6042 15186 6054 15220
rect 5996 15152 6054 15186
rect 6154 15220 6212 15252
rect 6154 15186 6166 15220
rect 6200 15186 6212 15220
rect 6154 15152 6212 15186
rect 6348 15222 6406 15254
rect 6348 15188 6360 15222
rect 6394 15188 6406 15222
rect 6348 15154 6406 15188
rect 6506 15222 6564 15254
rect 6506 15188 6518 15222
rect 6552 15188 6564 15222
rect 6506 15154 6564 15188
rect 6656 15222 6714 15254
rect 6656 15188 6668 15222
rect 6702 15188 6714 15222
rect 6656 15154 6714 15188
rect 6814 15222 6872 15254
rect 6814 15188 6826 15222
rect 6860 15188 6872 15222
rect 6814 15154 6872 15188
rect 988 15068 1013 15102
rect 1047 15068 1072 15102
rect 988 15056 1072 15068
rect 544 14436 628 14448
rect 544 14402 569 14436
rect 603 14402 628 14436
rect 544 14345 628 14402
rect 544 13868 628 13925
rect 544 13834 569 13868
rect 603 13834 628 13868
rect 544 13822 628 13834
rect 690 14436 774 14448
rect 690 14402 715 14436
rect 749 14402 774 14436
rect 690 14345 774 14402
rect 690 13868 774 13925
rect 690 13834 715 13868
rect 749 13834 774 13868
rect 690 13822 774 13834
rect 834 14442 918 14454
rect 834 14408 859 14442
rect 893 14408 918 14442
rect 834 14351 918 14408
rect 834 13874 918 13931
rect 834 13840 859 13874
rect 893 13840 918 13874
rect 834 13828 918 13840
rect 988 14442 1072 14454
rect 988 14408 1013 14442
rect 1047 14408 1072 14442
rect 988 14351 1072 14408
rect 988 13874 1072 13931
rect 1398 13981 1456 14014
rect 1398 13947 1410 13981
rect 1444 13947 1456 13981
rect 1398 13914 1456 13947
rect 1556 13981 1614 14014
rect 1556 13947 1568 13981
rect 1602 13947 1614 13981
rect 1556 13914 1614 13947
rect 1686 13981 1744 14014
rect 1686 13947 1698 13981
rect 1732 13947 1744 13981
rect 1686 13914 1744 13947
rect 1844 13981 1902 14014
rect 1844 13947 1856 13981
rect 1890 13947 1902 13981
rect 1844 13914 1902 13947
rect 2018 13981 2076 14014
rect 2018 13947 2030 13981
rect 2064 13947 2076 13981
rect 2018 13914 2076 13947
rect 2176 13981 2234 14014
rect 2176 13947 2188 13981
rect 2222 13947 2234 13981
rect 2176 13914 2234 13947
rect 2360 13981 2418 14014
rect 2360 13947 2372 13981
rect 2406 13947 2418 13981
rect 2360 13914 2418 13947
rect 2518 13981 2576 14014
rect 2518 13947 2530 13981
rect 2564 13947 2576 13981
rect 2518 13914 2576 13947
rect 2764 13981 2822 14014
rect 2764 13947 2776 13981
rect 2810 13947 2822 13981
rect 2764 13914 2822 13947
rect 2922 13981 2980 14014
rect 2922 13947 2934 13981
rect 2968 13947 2980 13981
rect 2922 13914 2980 13947
rect 3108 13981 3166 14014
rect 3108 13947 3120 13981
rect 3154 13947 3166 13981
rect 3108 13914 3166 13947
rect 3266 13981 3324 14014
rect 3266 13947 3278 13981
rect 3312 13947 3324 13981
rect 3266 13914 3324 13947
rect 3730 13991 3788 14024
rect 3730 13957 3742 13991
rect 3776 13957 3788 13991
rect 3730 13924 3788 13957
rect 3888 13991 3946 14024
rect 3888 13957 3900 13991
rect 3934 13957 3946 13991
rect 3888 13924 3946 13957
rect 4038 13991 4096 14024
rect 4038 13957 4050 13991
rect 4084 13957 4096 13991
rect 4038 13924 4096 13957
rect 4196 13991 4254 14024
rect 4196 13957 4208 13991
rect 4242 13957 4254 13991
rect 4196 13924 4254 13957
rect 4390 13993 4448 14026
rect 4390 13959 4402 13993
rect 4436 13959 4448 13993
rect 4390 13926 4448 13959
rect 4548 13993 4606 14026
rect 4548 13959 4560 13993
rect 4594 13959 4606 13993
rect 4548 13926 4606 13959
rect 4698 13993 4756 14026
rect 4698 13959 4710 13993
rect 4744 13959 4756 13993
rect 4698 13926 4756 13959
rect 4856 13993 4914 14026
rect 4856 13959 4868 13993
rect 4902 13959 4914 13993
rect 4856 13926 4914 13959
rect 5688 13992 5746 14024
rect 5688 13958 5700 13992
rect 5734 13958 5746 13992
rect 5688 13924 5746 13958
rect 5846 13992 5904 14024
rect 5846 13958 5858 13992
rect 5892 13958 5904 13992
rect 5846 13924 5904 13958
rect 5996 13992 6054 14024
rect 5996 13958 6008 13992
rect 6042 13958 6054 13992
rect 5996 13924 6054 13958
rect 6154 13992 6212 14024
rect 6154 13958 6166 13992
rect 6200 13958 6212 13992
rect 6154 13924 6212 13958
rect 6348 13994 6406 14026
rect 6348 13960 6360 13994
rect 6394 13960 6406 13994
rect 6348 13926 6406 13960
rect 6506 13994 6564 14026
rect 6506 13960 6518 13994
rect 6552 13960 6564 13994
rect 6506 13926 6564 13960
rect 6656 13994 6714 14026
rect 6656 13960 6668 13994
rect 6702 13960 6714 13994
rect 6656 13926 6714 13960
rect 6814 13994 6872 14026
rect 6814 13960 6826 13994
rect 6860 13960 6872 13994
rect 6814 13926 6872 13960
rect 988 13840 1013 13874
rect 1047 13840 1072 13874
rect 988 13828 1072 13840
rect 544 13208 628 13220
rect 544 13174 569 13208
rect 603 13174 628 13208
rect 544 13117 628 13174
rect 544 12640 628 12697
rect 544 12606 569 12640
rect 603 12606 628 12640
rect 544 12594 628 12606
rect 690 13208 774 13220
rect 690 13174 715 13208
rect 749 13174 774 13208
rect 690 13117 774 13174
rect 690 12640 774 12697
rect 690 12606 715 12640
rect 749 12606 774 12640
rect 690 12594 774 12606
rect 834 13214 918 13226
rect 834 13180 859 13214
rect 893 13180 918 13214
rect 834 13123 918 13180
rect 834 12646 918 12703
rect 834 12612 859 12646
rect 893 12612 918 12646
rect 834 12600 918 12612
rect 988 13214 1072 13226
rect 988 13180 1013 13214
rect 1047 13180 1072 13214
rect 988 13123 1072 13180
rect 988 12646 1072 12703
rect 1398 12753 1456 12786
rect 1398 12719 1410 12753
rect 1444 12719 1456 12753
rect 1398 12686 1456 12719
rect 1556 12753 1614 12786
rect 1556 12719 1568 12753
rect 1602 12719 1614 12753
rect 1556 12686 1614 12719
rect 1686 12753 1744 12786
rect 1686 12719 1698 12753
rect 1732 12719 1744 12753
rect 1686 12686 1744 12719
rect 1844 12753 1902 12786
rect 1844 12719 1856 12753
rect 1890 12719 1902 12753
rect 1844 12686 1902 12719
rect 2018 12753 2076 12786
rect 2018 12719 2030 12753
rect 2064 12719 2076 12753
rect 2018 12686 2076 12719
rect 2176 12753 2234 12786
rect 2176 12719 2188 12753
rect 2222 12719 2234 12753
rect 2176 12686 2234 12719
rect 2360 12753 2418 12786
rect 2360 12719 2372 12753
rect 2406 12719 2418 12753
rect 2360 12686 2418 12719
rect 2518 12753 2576 12786
rect 2518 12719 2530 12753
rect 2564 12719 2576 12753
rect 2518 12686 2576 12719
rect 2764 12753 2822 12786
rect 2764 12719 2776 12753
rect 2810 12719 2822 12753
rect 2764 12686 2822 12719
rect 2922 12753 2980 12786
rect 2922 12719 2934 12753
rect 2968 12719 2980 12753
rect 2922 12686 2980 12719
rect 3108 12753 3166 12786
rect 3108 12719 3120 12753
rect 3154 12719 3166 12753
rect 3108 12686 3166 12719
rect 3266 12753 3324 12786
rect 3266 12719 3278 12753
rect 3312 12719 3324 12753
rect 3266 12686 3324 12719
rect 3730 12763 3788 12796
rect 3730 12729 3742 12763
rect 3776 12729 3788 12763
rect 3730 12696 3788 12729
rect 3888 12763 3946 12796
rect 3888 12729 3900 12763
rect 3934 12729 3946 12763
rect 3888 12696 3946 12729
rect 4038 12763 4096 12796
rect 4038 12729 4050 12763
rect 4084 12729 4096 12763
rect 4038 12696 4096 12729
rect 4196 12763 4254 12796
rect 4196 12729 4208 12763
rect 4242 12729 4254 12763
rect 4196 12696 4254 12729
rect 4390 12765 4448 12798
rect 4390 12731 4402 12765
rect 4436 12731 4448 12765
rect 4390 12698 4448 12731
rect 4548 12765 4606 12798
rect 4548 12731 4560 12765
rect 4594 12731 4606 12765
rect 4548 12698 4606 12731
rect 4698 12765 4756 12798
rect 4698 12731 4710 12765
rect 4744 12731 4756 12765
rect 4698 12698 4756 12731
rect 4856 12765 4914 12798
rect 4856 12731 4868 12765
rect 4902 12731 4914 12765
rect 4856 12698 4914 12731
rect 5688 12764 5746 12796
rect 5688 12730 5700 12764
rect 5734 12730 5746 12764
rect 5688 12696 5746 12730
rect 5846 12764 5904 12796
rect 5846 12730 5858 12764
rect 5892 12730 5904 12764
rect 5846 12696 5904 12730
rect 5996 12764 6054 12796
rect 5996 12730 6008 12764
rect 6042 12730 6054 12764
rect 5996 12696 6054 12730
rect 6154 12764 6212 12796
rect 6154 12730 6166 12764
rect 6200 12730 6212 12764
rect 6154 12696 6212 12730
rect 6348 12766 6406 12798
rect 6348 12732 6360 12766
rect 6394 12732 6406 12766
rect 6348 12698 6406 12732
rect 6506 12766 6564 12798
rect 6506 12732 6518 12766
rect 6552 12732 6564 12766
rect 6506 12698 6564 12732
rect 6656 12766 6714 12798
rect 6656 12732 6668 12766
rect 6702 12732 6714 12766
rect 6656 12698 6714 12732
rect 6814 12766 6872 12798
rect 6814 12732 6826 12766
rect 6860 12732 6872 12766
rect 6814 12698 6872 12732
rect 988 12612 1013 12646
rect 1047 12612 1072 12646
rect 988 12600 1072 12612
rect 544 11980 628 11992
rect 544 11946 569 11980
rect 603 11946 628 11980
rect 544 11889 628 11946
rect 544 11412 628 11469
rect 544 11378 569 11412
rect 603 11378 628 11412
rect 544 11366 628 11378
rect 690 11980 774 11992
rect 690 11946 715 11980
rect 749 11946 774 11980
rect 690 11889 774 11946
rect 690 11412 774 11469
rect 690 11378 715 11412
rect 749 11378 774 11412
rect 690 11366 774 11378
rect 834 11986 918 11998
rect 834 11952 859 11986
rect 893 11952 918 11986
rect 834 11895 918 11952
rect 834 11418 918 11475
rect 834 11384 859 11418
rect 893 11384 918 11418
rect 834 11372 918 11384
rect 988 11986 1072 11998
rect 988 11952 1013 11986
rect 1047 11952 1072 11986
rect 988 11895 1072 11952
rect 988 11418 1072 11475
rect 1398 11525 1456 11558
rect 1398 11491 1410 11525
rect 1444 11491 1456 11525
rect 1398 11458 1456 11491
rect 1556 11525 1614 11558
rect 1556 11491 1568 11525
rect 1602 11491 1614 11525
rect 1556 11458 1614 11491
rect 1686 11525 1744 11558
rect 1686 11491 1698 11525
rect 1732 11491 1744 11525
rect 1686 11458 1744 11491
rect 1844 11525 1902 11558
rect 1844 11491 1856 11525
rect 1890 11491 1902 11525
rect 1844 11458 1902 11491
rect 2018 11525 2076 11558
rect 2018 11491 2030 11525
rect 2064 11491 2076 11525
rect 2018 11458 2076 11491
rect 2176 11525 2234 11558
rect 2176 11491 2188 11525
rect 2222 11491 2234 11525
rect 2176 11458 2234 11491
rect 2360 11525 2418 11558
rect 2360 11491 2372 11525
rect 2406 11491 2418 11525
rect 2360 11458 2418 11491
rect 2518 11525 2576 11558
rect 2518 11491 2530 11525
rect 2564 11491 2576 11525
rect 2518 11458 2576 11491
rect 2764 11525 2822 11558
rect 2764 11491 2776 11525
rect 2810 11491 2822 11525
rect 2764 11458 2822 11491
rect 2922 11525 2980 11558
rect 2922 11491 2934 11525
rect 2968 11491 2980 11525
rect 2922 11458 2980 11491
rect 3108 11525 3166 11558
rect 3108 11491 3120 11525
rect 3154 11491 3166 11525
rect 3108 11458 3166 11491
rect 3266 11525 3324 11558
rect 3266 11491 3278 11525
rect 3312 11491 3324 11525
rect 3266 11458 3324 11491
rect 3730 11535 3788 11568
rect 3730 11501 3742 11535
rect 3776 11501 3788 11535
rect 3730 11468 3788 11501
rect 3888 11535 3946 11568
rect 3888 11501 3900 11535
rect 3934 11501 3946 11535
rect 3888 11468 3946 11501
rect 4038 11535 4096 11568
rect 4038 11501 4050 11535
rect 4084 11501 4096 11535
rect 4038 11468 4096 11501
rect 4196 11535 4254 11568
rect 4196 11501 4208 11535
rect 4242 11501 4254 11535
rect 4196 11468 4254 11501
rect 4390 11537 4448 11570
rect 4390 11503 4402 11537
rect 4436 11503 4448 11537
rect 4390 11470 4448 11503
rect 4548 11537 4606 11570
rect 4548 11503 4560 11537
rect 4594 11503 4606 11537
rect 4548 11470 4606 11503
rect 4698 11537 4756 11570
rect 4698 11503 4710 11537
rect 4744 11503 4756 11537
rect 4698 11470 4756 11503
rect 4856 11537 4914 11570
rect 4856 11503 4868 11537
rect 4902 11503 4914 11537
rect 4856 11470 4914 11503
rect 5688 11536 5746 11568
rect 5688 11502 5700 11536
rect 5734 11502 5746 11536
rect 5688 11468 5746 11502
rect 5846 11536 5904 11568
rect 5846 11502 5858 11536
rect 5892 11502 5904 11536
rect 5846 11468 5904 11502
rect 5996 11536 6054 11568
rect 5996 11502 6008 11536
rect 6042 11502 6054 11536
rect 5996 11468 6054 11502
rect 6154 11536 6212 11568
rect 6154 11502 6166 11536
rect 6200 11502 6212 11536
rect 6154 11468 6212 11502
rect 6348 11538 6406 11570
rect 6348 11504 6360 11538
rect 6394 11504 6406 11538
rect 6348 11470 6406 11504
rect 6506 11538 6564 11570
rect 6506 11504 6518 11538
rect 6552 11504 6564 11538
rect 6506 11470 6564 11504
rect 6656 11538 6714 11570
rect 6656 11504 6668 11538
rect 6702 11504 6714 11538
rect 6656 11470 6714 11504
rect 6814 11538 6872 11570
rect 6814 11504 6826 11538
rect 6860 11504 6872 11538
rect 6814 11470 6872 11504
rect 988 11384 1013 11418
rect 1047 11384 1072 11418
rect 988 11372 1072 11384
rect 544 10752 628 10764
rect 544 10718 569 10752
rect 603 10718 628 10752
rect 544 10661 628 10718
rect 544 10184 628 10241
rect 544 10150 569 10184
rect 603 10150 628 10184
rect 544 10138 628 10150
rect 690 10752 774 10764
rect 690 10718 715 10752
rect 749 10718 774 10752
rect 690 10661 774 10718
rect 690 10184 774 10241
rect 690 10150 715 10184
rect 749 10150 774 10184
rect 690 10138 774 10150
rect 834 10758 918 10770
rect 834 10724 859 10758
rect 893 10724 918 10758
rect 834 10667 918 10724
rect 834 10190 918 10247
rect 834 10156 859 10190
rect 893 10156 918 10190
rect 834 10144 918 10156
rect 988 10758 1072 10770
rect 988 10724 1013 10758
rect 1047 10724 1072 10758
rect 988 10667 1072 10724
rect 988 10190 1072 10247
rect 1398 10297 1456 10330
rect 1398 10263 1410 10297
rect 1444 10263 1456 10297
rect 1398 10230 1456 10263
rect 1556 10297 1614 10330
rect 1556 10263 1568 10297
rect 1602 10263 1614 10297
rect 1556 10230 1614 10263
rect 1686 10297 1744 10330
rect 1686 10263 1698 10297
rect 1732 10263 1744 10297
rect 1686 10230 1744 10263
rect 1844 10297 1902 10330
rect 1844 10263 1856 10297
rect 1890 10263 1902 10297
rect 1844 10230 1902 10263
rect 2018 10297 2076 10330
rect 2018 10263 2030 10297
rect 2064 10263 2076 10297
rect 2018 10230 2076 10263
rect 2176 10297 2234 10330
rect 2176 10263 2188 10297
rect 2222 10263 2234 10297
rect 2176 10230 2234 10263
rect 2360 10297 2418 10330
rect 2360 10263 2372 10297
rect 2406 10263 2418 10297
rect 2360 10230 2418 10263
rect 2518 10297 2576 10330
rect 2518 10263 2530 10297
rect 2564 10263 2576 10297
rect 2518 10230 2576 10263
rect 2764 10297 2822 10330
rect 2764 10263 2776 10297
rect 2810 10263 2822 10297
rect 2764 10230 2822 10263
rect 2922 10297 2980 10330
rect 2922 10263 2934 10297
rect 2968 10263 2980 10297
rect 2922 10230 2980 10263
rect 3108 10297 3166 10330
rect 3108 10263 3120 10297
rect 3154 10263 3166 10297
rect 3108 10230 3166 10263
rect 3266 10297 3324 10330
rect 3266 10263 3278 10297
rect 3312 10263 3324 10297
rect 3266 10230 3324 10263
rect 3730 10307 3788 10340
rect 3730 10273 3742 10307
rect 3776 10273 3788 10307
rect 3730 10240 3788 10273
rect 3888 10307 3946 10340
rect 3888 10273 3900 10307
rect 3934 10273 3946 10307
rect 3888 10240 3946 10273
rect 4038 10307 4096 10340
rect 4038 10273 4050 10307
rect 4084 10273 4096 10307
rect 4038 10240 4096 10273
rect 4196 10307 4254 10340
rect 4196 10273 4208 10307
rect 4242 10273 4254 10307
rect 4196 10240 4254 10273
rect 4390 10309 4448 10342
rect 4390 10275 4402 10309
rect 4436 10275 4448 10309
rect 4390 10242 4448 10275
rect 4548 10309 4606 10342
rect 4548 10275 4560 10309
rect 4594 10275 4606 10309
rect 4548 10242 4606 10275
rect 4698 10309 4756 10342
rect 4698 10275 4710 10309
rect 4744 10275 4756 10309
rect 4698 10242 4756 10275
rect 4856 10309 4914 10342
rect 4856 10275 4868 10309
rect 4902 10275 4914 10309
rect 4856 10242 4914 10275
rect 5688 10308 5746 10340
rect 5688 10274 5700 10308
rect 5734 10274 5746 10308
rect 5688 10240 5746 10274
rect 5846 10308 5904 10340
rect 5846 10274 5858 10308
rect 5892 10274 5904 10308
rect 5846 10240 5904 10274
rect 5996 10308 6054 10340
rect 5996 10274 6008 10308
rect 6042 10274 6054 10308
rect 5996 10240 6054 10274
rect 6154 10308 6212 10340
rect 6154 10274 6166 10308
rect 6200 10274 6212 10308
rect 6154 10240 6212 10274
rect 6348 10310 6406 10342
rect 6348 10276 6360 10310
rect 6394 10276 6406 10310
rect 6348 10242 6406 10276
rect 6506 10310 6564 10342
rect 6506 10276 6518 10310
rect 6552 10276 6564 10310
rect 6506 10242 6564 10276
rect 6656 10310 6714 10342
rect 6656 10276 6668 10310
rect 6702 10276 6714 10310
rect 6656 10242 6714 10276
rect 6814 10310 6872 10342
rect 6814 10276 6826 10310
rect 6860 10276 6872 10310
rect 6814 10242 6872 10276
rect 988 10156 1013 10190
rect 1047 10156 1072 10190
rect 988 10144 1072 10156
rect 544 9524 628 9536
rect 544 9490 569 9524
rect 603 9490 628 9524
rect 544 9433 628 9490
rect 544 8956 628 9013
rect 544 8922 569 8956
rect 603 8922 628 8956
rect 544 8910 628 8922
rect 690 9524 774 9536
rect 690 9490 715 9524
rect 749 9490 774 9524
rect 690 9433 774 9490
rect 690 8956 774 9013
rect 690 8922 715 8956
rect 749 8922 774 8956
rect 690 8910 774 8922
rect 834 9530 918 9542
rect 834 9496 859 9530
rect 893 9496 918 9530
rect 834 9439 918 9496
rect 834 8962 918 9019
rect 834 8928 859 8962
rect 893 8928 918 8962
rect 834 8916 918 8928
rect 988 9530 1072 9542
rect 988 9496 1013 9530
rect 1047 9496 1072 9530
rect 988 9439 1072 9496
rect 988 8962 1072 9019
rect 1398 9069 1456 9102
rect 1398 9035 1410 9069
rect 1444 9035 1456 9069
rect 1398 9002 1456 9035
rect 1556 9069 1614 9102
rect 1556 9035 1568 9069
rect 1602 9035 1614 9069
rect 1556 9002 1614 9035
rect 1686 9069 1744 9102
rect 1686 9035 1698 9069
rect 1732 9035 1744 9069
rect 1686 9002 1744 9035
rect 1844 9069 1902 9102
rect 1844 9035 1856 9069
rect 1890 9035 1902 9069
rect 1844 9002 1902 9035
rect 2018 9069 2076 9102
rect 2018 9035 2030 9069
rect 2064 9035 2076 9069
rect 2018 9002 2076 9035
rect 2176 9069 2234 9102
rect 2176 9035 2188 9069
rect 2222 9035 2234 9069
rect 2176 9002 2234 9035
rect 2360 9069 2418 9102
rect 2360 9035 2372 9069
rect 2406 9035 2418 9069
rect 2360 9002 2418 9035
rect 2518 9069 2576 9102
rect 2518 9035 2530 9069
rect 2564 9035 2576 9069
rect 2518 9002 2576 9035
rect 2764 9069 2822 9102
rect 2764 9035 2776 9069
rect 2810 9035 2822 9069
rect 2764 9002 2822 9035
rect 2922 9069 2980 9102
rect 2922 9035 2934 9069
rect 2968 9035 2980 9069
rect 2922 9002 2980 9035
rect 3108 9069 3166 9102
rect 3108 9035 3120 9069
rect 3154 9035 3166 9069
rect 3108 9002 3166 9035
rect 3266 9069 3324 9102
rect 3266 9035 3278 9069
rect 3312 9035 3324 9069
rect 3266 9002 3324 9035
rect 3730 9079 3788 9112
rect 3730 9045 3742 9079
rect 3776 9045 3788 9079
rect 3730 9012 3788 9045
rect 3888 9079 3946 9112
rect 3888 9045 3900 9079
rect 3934 9045 3946 9079
rect 3888 9012 3946 9045
rect 4038 9079 4096 9112
rect 4038 9045 4050 9079
rect 4084 9045 4096 9079
rect 4038 9012 4096 9045
rect 4196 9079 4254 9112
rect 4196 9045 4208 9079
rect 4242 9045 4254 9079
rect 4196 9012 4254 9045
rect 4390 9081 4448 9114
rect 4390 9047 4402 9081
rect 4436 9047 4448 9081
rect 4390 9014 4448 9047
rect 4548 9081 4606 9114
rect 4548 9047 4560 9081
rect 4594 9047 4606 9081
rect 4548 9014 4606 9047
rect 4698 9081 4756 9114
rect 4698 9047 4710 9081
rect 4744 9047 4756 9081
rect 4698 9014 4756 9047
rect 4856 9081 4914 9114
rect 4856 9047 4868 9081
rect 4902 9047 4914 9081
rect 4856 9014 4914 9047
rect 5688 9080 5746 9112
rect 5688 9046 5700 9080
rect 5734 9046 5746 9080
rect 5688 9012 5746 9046
rect 5846 9080 5904 9112
rect 5846 9046 5858 9080
rect 5892 9046 5904 9080
rect 5846 9012 5904 9046
rect 5996 9080 6054 9112
rect 5996 9046 6008 9080
rect 6042 9046 6054 9080
rect 5996 9012 6054 9046
rect 6154 9080 6212 9112
rect 6154 9046 6166 9080
rect 6200 9046 6212 9080
rect 6154 9012 6212 9046
rect 6348 9082 6406 9114
rect 6348 9048 6360 9082
rect 6394 9048 6406 9082
rect 6348 9014 6406 9048
rect 6506 9082 6564 9114
rect 6506 9048 6518 9082
rect 6552 9048 6564 9082
rect 6506 9014 6564 9048
rect 6656 9082 6714 9114
rect 6656 9048 6668 9082
rect 6702 9048 6714 9082
rect 6656 9014 6714 9048
rect 6814 9082 6872 9114
rect 6814 9048 6826 9082
rect 6860 9048 6872 9082
rect 6814 9014 6872 9048
rect 988 8928 1013 8962
rect 1047 8928 1072 8962
rect 988 8916 1072 8928
rect 544 8296 628 8308
rect 544 8262 569 8296
rect 603 8262 628 8296
rect 544 8205 628 8262
rect 544 7728 628 7785
rect 544 7694 569 7728
rect 603 7694 628 7728
rect 544 7682 628 7694
rect 690 8296 774 8308
rect 690 8262 715 8296
rect 749 8262 774 8296
rect 690 8205 774 8262
rect 690 7728 774 7785
rect 690 7694 715 7728
rect 749 7694 774 7728
rect 690 7682 774 7694
rect 834 8302 918 8314
rect 834 8268 859 8302
rect 893 8268 918 8302
rect 834 8211 918 8268
rect 834 7734 918 7791
rect 834 7700 859 7734
rect 893 7700 918 7734
rect 834 7688 918 7700
rect 988 8302 1072 8314
rect 988 8268 1013 8302
rect 1047 8268 1072 8302
rect 988 8211 1072 8268
rect 988 7734 1072 7791
rect 1398 7841 1456 7874
rect 1398 7807 1410 7841
rect 1444 7807 1456 7841
rect 1398 7774 1456 7807
rect 1556 7841 1614 7874
rect 1556 7807 1568 7841
rect 1602 7807 1614 7841
rect 1556 7774 1614 7807
rect 1686 7841 1744 7874
rect 1686 7807 1698 7841
rect 1732 7807 1744 7841
rect 1686 7774 1744 7807
rect 1844 7841 1902 7874
rect 1844 7807 1856 7841
rect 1890 7807 1902 7841
rect 1844 7774 1902 7807
rect 2018 7841 2076 7874
rect 2018 7807 2030 7841
rect 2064 7807 2076 7841
rect 2018 7774 2076 7807
rect 2176 7841 2234 7874
rect 2176 7807 2188 7841
rect 2222 7807 2234 7841
rect 2176 7774 2234 7807
rect 2360 7841 2418 7874
rect 2360 7807 2372 7841
rect 2406 7807 2418 7841
rect 2360 7774 2418 7807
rect 2518 7841 2576 7874
rect 2518 7807 2530 7841
rect 2564 7807 2576 7841
rect 2518 7774 2576 7807
rect 2764 7841 2822 7874
rect 2764 7807 2776 7841
rect 2810 7807 2822 7841
rect 2764 7774 2822 7807
rect 2922 7841 2980 7874
rect 2922 7807 2934 7841
rect 2968 7807 2980 7841
rect 2922 7774 2980 7807
rect 3108 7841 3166 7874
rect 3108 7807 3120 7841
rect 3154 7807 3166 7841
rect 3108 7774 3166 7807
rect 3266 7841 3324 7874
rect 3266 7807 3278 7841
rect 3312 7807 3324 7841
rect 3266 7774 3324 7807
rect 3730 7851 3788 7884
rect 3730 7817 3742 7851
rect 3776 7817 3788 7851
rect 3730 7784 3788 7817
rect 3888 7851 3946 7884
rect 3888 7817 3900 7851
rect 3934 7817 3946 7851
rect 3888 7784 3946 7817
rect 4038 7851 4096 7884
rect 4038 7817 4050 7851
rect 4084 7817 4096 7851
rect 4038 7784 4096 7817
rect 4196 7851 4254 7884
rect 4196 7817 4208 7851
rect 4242 7817 4254 7851
rect 4196 7784 4254 7817
rect 4390 7853 4448 7886
rect 4390 7819 4402 7853
rect 4436 7819 4448 7853
rect 4390 7786 4448 7819
rect 4548 7853 4606 7886
rect 4548 7819 4560 7853
rect 4594 7819 4606 7853
rect 4548 7786 4606 7819
rect 4698 7853 4756 7886
rect 4698 7819 4710 7853
rect 4744 7819 4756 7853
rect 4698 7786 4756 7819
rect 4856 7853 4914 7886
rect 4856 7819 4868 7853
rect 4902 7819 4914 7853
rect 4856 7786 4914 7819
rect 5688 7852 5746 7884
rect 5688 7818 5700 7852
rect 5734 7818 5746 7852
rect 5688 7784 5746 7818
rect 5846 7852 5904 7884
rect 5846 7818 5858 7852
rect 5892 7818 5904 7852
rect 5846 7784 5904 7818
rect 5996 7852 6054 7884
rect 5996 7818 6008 7852
rect 6042 7818 6054 7852
rect 5996 7784 6054 7818
rect 6154 7852 6212 7884
rect 6154 7818 6166 7852
rect 6200 7818 6212 7852
rect 6154 7784 6212 7818
rect 6348 7854 6406 7886
rect 6348 7820 6360 7854
rect 6394 7820 6406 7854
rect 6348 7786 6406 7820
rect 6506 7854 6564 7886
rect 6506 7820 6518 7854
rect 6552 7820 6564 7854
rect 6506 7786 6564 7820
rect 6656 7854 6714 7886
rect 6656 7820 6668 7854
rect 6702 7820 6714 7854
rect 6656 7786 6714 7820
rect 6814 7854 6872 7886
rect 6814 7820 6826 7854
rect 6860 7820 6872 7854
rect 6814 7786 6872 7820
rect 988 7700 1013 7734
rect 1047 7700 1072 7734
rect 988 7688 1072 7700
rect 544 7068 628 7080
rect 544 7034 569 7068
rect 603 7034 628 7068
rect 544 6977 628 7034
rect 544 6500 628 6557
rect 544 6466 569 6500
rect 603 6466 628 6500
rect 544 6454 628 6466
rect 690 7068 774 7080
rect 690 7034 715 7068
rect 749 7034 774 7068
rect 690 6977 774 7034
rect 690 6500 774 6557
rect 690 6466 715 6500
rect 749 6466 774 6500
rect 690 6454 774 6466
rect 834 7074 918 7086
rect 834 7040 859 7074
rect 893 7040 918 7074
rect 834 6983 918 7040
rect 834 6506 918 6563
rect 834 6472 859 6506
rect 893 6472 918 6506
rect 834 6460 918 6472
rect 988 7074 1072 7086
rect 988 7040 1013 7074
rect 1047 7040 1072 7074
rect 988 6983 1072 7040
rect 988 6506 1072 6563
rect 1398 6613 1456 6646
rect 1398 6579 1410 6613
rect 1444 6579 1456 6613
rect 1398 6546 1456 6579
rect 1556 6613 1614 6646
rect 1556 6579 1568 6613
rect 1602 6579 1614 6613
rect 1556 6546 1614 6579
rect 1686 6613 1744 6646
rect 1686 6579 1698 6613
rect 1732 6579 1744 6613
rect 1686 6546 1744 6579
rect 1844 6613 1902 6646
rect 1844 6579 1856 6613
rect 1890 6579 1902 6613
rect 1844 6546 1902 6579
rect 2018 6613 2076 6646
rect 2018 6579 2030 6613
rect 2064 6579 2076 6613
rect 2018 6546 2076 6579
rect 2176 6613 2234 6646
rect 2176 6579 2188 6613
rect 2222 6579 2234 6613
rect 2176 6546 2234 6579
rect 2360 6613 2418 6646
rect 2360 6579 2372 6613
rect 2406 6579 2418 6613
rect 2360 6546 2418 6579
rect 2518 6613 2576 6646
rect 2518 6579 2530 6613
rect 2564 6579 2576 6613
rect 2518 6546 2576 6579
rect 2764 6613 2822 6646
rect 2764 6579 2776 6613
rect 2810 6579 2822 6613
rect 2764 6546 2822 6579
rect 2922 6613 2980 6646
rect 2922 6579 2934 6613
rect 2968 6579 2980 6613
rect 2922 6546 2980 6579
rect 3108 6613 3166 6646
rect 3108 6579 3120 6613
rect 3154 6579 3166 6613
rect 3108 6546 3166 6579
rect 3266 6613 3324 6646
rect 3266 6579 3278 6613
rect 3312 6579 3324 6613
rect 3266 6546 3324 6579
rect 3730 6623 3788 6656
rect 3730 6589 3742 6623
rect 3776 6589 3788 6623
rect 3730 6556 3788 6589
rect 3888 6623 3946 6656
rect 3888 6589 3900 6623
rect 3934 6589 3946 6623
rect 3888 6556 3946 6589
rect 4038 6623 4096 6656
rect 4038 6589 4050 6623
rect 4084 6589 4096 6623
rect 4038 6556 4096 6589
rect 4196 6623 4254 6656
rect 4196 6589 4208 6623
rect 4242 6589 4254 6623
rect 4196 6556 4254 6589
rect 4390 6625 4448 6658
rect 4390 6591 4402 6625
rect 4436 6591 4448 6625
rect 4390 6558 4448 6591
rect 4548 6625 4606 6658
rect 4548 6591 4560 6625
rect 4594 6591 4606 6625
rect 4548 6558 4606 6591
rect 4698 6625 4756 6658
rect 4698 6591 4710 6625
rect 4744 6591 4756 6625
rect 4698 6558 4756 6591
rect 4856 6625 4914 6658
rect 4856 6591 4868 6625
rect 4902 6591 4914 6625
rect 4856 6558 4914 6591
rect 5688 6624 5746 6656
rect 5688 6590 5700 6624
rect 5734 6590 5746 6624
rect 5688 6556 5746 6590
rect 5846 6624 5904 6656
rect 5846 6590 5858 6624
rect 5892 6590 5904 6624
rect 5846 6556 5904 6590
rect 5996 6624 6054 6656
rect 5996 6590 6008 6624
rect 6042 6590 6054 6624
rect 5996 6556 6054 6590
rect 6154 6624 6212 6656
rect 6154 6590 6166 6624
rect 6200 6590 6212 6624
rect 6154 6556 6212 6590
rect 6348 6626 6406 6658
rect 6348 6592 6360 6626
rect 6394 6592 6406 6626
rect 6348 6558 6406 6592
rect 6506 6626 6564 6658
rect 6506 6592 6518 6626
rect 6552 6592 6564 6626
rect 6506 6558 6564 6592
rect 6656 6626 6714 6658
rect 6656 6592 6668 6626
rect 6702 6592 6714 6626
rect 6656 6558 6714 6592
rect 6814 6626 6872 6658
rect 6814 6592 6826 6626
rect 6860 6592 6872 6626
rect 6814 6558 6872 6592
rect 988 6472 1013 6506
rect 1047 6472 1072 6506
rect 988 6460 1072 6472
rect 544 5840 628 5852
rect 544 5806 569 5840
rect 603 5806 628 5840
rect 544 5749 628 5806
rect 544 5272 628 5329
rect 544 5238 569 5272
rect 603 5238 628 5272
rect 544 5226 628 5238
rect 690 5840 774 5852
rect 690 5806 715 5840
rect 749 5806 774 5840
rect 690 5749 774 5806
rect 690 5272 774 5329
rect 690 5238 715 5272
rect 749 5238 774 5272
rect 690 5226 774 5238
rect 834 5846 918 5858
rect 834 5812 859 5846
rect 893 5812 918 5846
rect 834 5755 918 5812
rect 834 5278 918 5335
rect 834 5244 859 5278
rect 893 5244 918 5278
rect 834 5232 918 5244
rect 988 5846 1072 5858
rect 988 5812 1013 5846
rect 1047 5812 1072 5846
rect 988 5755 1072 5812
rect 988 5278 1072 5335
rect 1398 5385 1456 5418
rect 1398 5351 1410 5385
rect 1444 5351 1456 5385
rect 1398 5318 1456 5351
rect 1556 5385 1614 5418
rect 1556 5351 1568 5385
rect 1602 5351 1614 5385
rect 1556 5318 1614 5351
rect 1686 5385 1744 5418
rect 1686 5351 1698 5385
rect 1732 5351 1744 5385
rect 1686 5318 1744 5351
rect 1844 5385 1902 5418
rect 1844 5351 1856 5385
rect 1890 5351 1902 5385
rect 1844 5318 1902 5351
rect 2018 5385 2076 5418
rect 2018 5351 2030 5385
rect 2064 5351 2076 5385
rect 2018 5318 2076 5351
rect 2176 5385 2234 5418
rect 2176 5351 2188 5385
rect 2222 5351 2234 5385
rect 2176 5318 2234 5351
rect 2360 5385 2418 5418
rect 2360 5351 2372 5385
rect 2406 5351 2418 5385
rect 2360 5318 2418 5351
rect 2518 5385 2576 5418
rect 2518 5351 2530 5385
rect 2564 5351 2576 5385
rect 2518 5318 2576 5351
rect 2764 5385 2822 5418
rect 2764 5351 2776 5385
rect 2810 5351 2822 5385
rect 2764 5318 2822 5351
rect 2922 5385 2980 5418
rect 2922 5351 2934 5385
rect 2968 5351 2980 5385
rect 2922 5318 2980 5351
rect 3108 5385 3166 5418
rect 3108 5351 3120 5385
rect 3154 5351 3166 5385
rect 3108 5318 3166 5351
rect 3266 5385 3324 5418
rect 3266 5351 3278 5385
rect 3312 5351 3324 5385
rect 3266 5318 3324 5351
rect 3730 5395 3788 5428
rect 3730 5361 3742 5395
rect 3776 5361 3788 5395
rect 3730 5328 3788 5361
rect 3888 5395 3946 5428
rect 3888 5361 3900 5395
rect 3934 5361 3946 5395
rect 3888 5328 3946 5361
rect 4038 5395 4096 5428
rect 4038 5361 4050 5395
rect 4084 5361 4096 5395
rect 4038 5328 4096 5361
rect 4196 5395 4254 5428
rect 4196 5361 4208 5395
rect 4242 5361 4254 5395
rect 4196 5328 4254 5361
rect 4390 5397 4448 5430
rect 4390 5363 4402 5397
rect 4436 5363 4448 5397
rect 4390 5330 4448 5363
rect 4548 5397 4606 5430
rect 4548 5363 4560 5397
rect 4594 5363 4606 5397
rect 4548 5330 4606 5363
rect 4698 5397 4756 5430
rect 4698 5363 4710 5397
rect 4744 5363 4756 5397
rect 4698 5330 4756 5363
rect 4856 5397 4914 5430
rect 4856 5363 4868 5397
rect 4902 5363 4914 5397
rect 4856 5330 4914 5363
rect 5688 5396 5746 5428
rect 5688 5362 5700 5396
rect 5734 5362 5746 5396
rect 5688 5328 5746 5362
rect 5846 5396 5904 5428
rect 5846 5362 5858 5396
rect 5892 5362 5904 5396
rect 5846 5328 5904 5362
rect 5996 5396 6054 5428
rect 5996 5362 6008 5396
rect 6042 5362 6054 5396
rect 5996 5328 6054 5362
rect 6154 5396 6212 5428
rect 6154 5362 6166 5396
rect 6200 5362 6212 5396
rect 6154 5328 6212 5362
rect 6348 5398 6406 5430
rect 6348 5364 6360 5398
rect 6394 5364 6406 5398
rect 6348 5330 6406 5364
rect 6506 5398 6564 5430
rect 6506 5364 6518 5398
rect 6552 5364 6564 5398
rect 6506 5330 6564 5364
rect 6656 5398 6714 5430
rect 6656 5364 6668 5398
rect 6702 5364 6714 5398
rect 6656 5330 6714 5364
rect 6814 5398 6872 5430
rect 6814 5364 6826 5398
rect 6860 5364 6872 5398
rect 6814 5330 6872 5364
rect 988 5244 1013 5278
rect 1047 5244 1072 5278
rect 988 5232 1072 5244
rect 544 4612 628 4624
rect 544 4578 569 4612
rect 603 4578 628 4612
rect 544 4521 628 4578
rect 544 4044 628 4101
rect 544 4010 569 4044
rect 603 4010 628 4044
rect 544 3998 628 4010
rect 690 4612 774 4624
rect 690 4578 715 4612
rect 749 4578 774 4612
rect 690 4521 774 4578
rect 690 4044 774 4101
rect 690 4010 715 4044
rect 749 4010 774 4044
rect 690 3998 774 4010
rect 834 4618 918 4630
rect 834 4584 859 4618
rect 893 4584 918 4618
rect 834 4527 918 4584
rect 834 4050 918 4107
rect 834 4016 859 4050
rect 893 4016 918 4050
rect 834 4004 918 4016
rect 988 4618 1072 4630
rect 988 4584 1013 4618
rect 1047 4584 1072 4618
rect 988 4527 1072 4584
rect 988 4050 1072 4107
rect 1398 4157 1456 4190
rect 1398 4123 1410 4157
rect 1444 4123 1456 4157
rect 1398 4090 1456 4123
rect 1556 4157 1614 4190
rect 1556 4123 1568 4157
rect 1602 4123 1614 4157
rect 1556 4090 1614 4123
rect 1686 4157 1744 4190
rect 1686 4123 1698 4157
rect 1732 4123 1744 4157
rect 1686 4090 1744 4123
rect 1844 4157 1902 4190
rect 1844 4123 1856 4157
rect 1890 4123 1902 4157
rect 1844 4090 1902 4123
rect 2018 4157 2076 4190
rect 2018 4123 2030 4157
rect 2064 4123 2076 4157
rect 2018 4090 2076 4123
rect 2176 4157 2234 4190
rect 2176 4123 2188 4157
rect 2222 4123 2234 4157
rect 2176 4090 2234 4123
rect 2360 4157 2418 4190
rect 2360 4123 2372 4157
rect 2406 4123 2418 4157
rect 2360 4090 2418 4123
rect 2518 4157 2576 4190
rect 2518 4123 2530 4157
rect 2564 4123 2576 4157
rect 2518 4090 2576 4123
rect 2764 4157 2822 4190
rect 2764 4123 2776 4157
rect 2810 4123 2822 4157
rect 2764 4090 2822 4123
rect 2922 4157 2980 4190
rect 2922 4123 2934 4157
rect 2968 4123 2980 4157
rect 2922 4090 2980 4123
rect 3108 4157 3166 4190
rect 3108 4123 3120 4157
rect 3154 4123 3166 4157
rect 3108 4090 3166 4123
rect 3266 4157 3324 4190
rect 3266 4123 3278 4157
rect 3312 4123 3324 4157
rect 3266 4090 3324 4123
rect 3730 4167 3788 4200
rect 3730 4133 3742 4167
rect 3776 4133 3788 4167
rect 3730 4100 3788 4133
rect 3888 4167 3946 4200
rect 3888 4133 3900 4167
rect 3934 4133 3946 4167
rect 3888 4100 3946 4133
rect 4038 4167 4096 4200
rect 4038 4133 4050 4167
rect 4084 4133 4096 4167
rect 4038 4100 4096 4133
rect 4196 4167 4254 4200
rect 4196 4133 4208 4167
rect 4242 4133 4254 4167
rect 4196 4100 4254 4133
rect 4390 4169 4448 4202
rect 4390 4135 4402 4169
rect 4436 4135 4448 4169
rect 4390 4102 4448 4135
rect 4548 4169 4606 4202
rect 4548 4135 4560 4169
rect 4594 4135 4606 4169
rect 4548 4102 4606 4135
rect 4698 4169 4756 4202
rect 4698 4135 4710 4169
rect 4744 4135 4756 4169
rect 4698 4102 4756 4135
rect 4856 4169 4914 4202
rect 4856 4135 4868 4169
rect 4902 4135 4914 4169
rect 4856 4102 4914 4135
rect 5688 4168 5746 4200
rect 5688 4134 5700 4168
rect 5734 4134 5746 4168
rect 5688 4100 5746 4134
rect 5846 4168 5904 4200
rect 5846 4134 5858 4168
rect 5892 4134 5904 4168
rect 5846 4100 5904 4134
rect 5996 4168 6054 4200
rect 5996 4134 6008 4168
rect 6042 4134 6054 4168
rect 5996 4100 6054 4134
rect 6154 4168 6212 4200
rect 6154 4134 6166 4168
rect 6200 4134 6212 4168
rect 6154 4100 6212 4134
rect 6348 4170 6406 4202
rect 6348 4136 6360 4170
rect 6394 4136 6406 4170
rect 6348 4102 6406 4136
rect 6506 4170 6564 4202
rect 6506 4136 6518 4170
rect 6552 4136 6564 4170
rect 6506 4102 6564 4136
rect 6656 4170 6714 4202
rect 6656 4136 6668 4170
rect 6702 4136 6714 4170
rect 6656 4102 6714 4136
rect 6814 4170 6872 4202
rect 6814 4136 6826 4170
rect 6860 4136 6872 4170
rect 6814 4102 6872 4136
rect 988 4016 1013 4050
rect 1047 4016 1072 4050
rect 988 4004 1072 4016
rect 544 3384 628 3396
rect 544 3350 569 3384
rect 603 3350 628 3384
rect 544 3293 628 3350
rect 544 2816 628 2873
rect 544 2782 569 2816
rect 603 2782 628 2816
rect 544 2770 628 2782
rect 690 3384 774 3396
rect 690 3350 715 3384
rect 749 3350 774 3384
rect 690 3293 774 3350
rect 690 2816 774 2873
rect 690 2782 715 2816
rect 749 2782 774 2816
rect 690 2770 774 2782
rect 834 3390 918 3402
rect 834 3356 859 3390
rect 893 3356 918 3390
rect 834 3299 918 3356
rect 834 2822 918 2879
rect 834 2788 859 2822
rect 893 2788 918 2822
rect 834 2776 918 2788
rect 988 3390 1072 3402
rect 988 3356 1013 3390
rect 1047 3356 1072 3390
rect 988 3299 1072 3356
rect 988 2822 1072 2879
rect 1398 2929 1456 2962
rect 1398 2895 1410 2929
rect 1444 2895 1456 2929
rect 1398 2862 1456 2895
rect 1556 2929 1614 2962
rect 1556 2895 1568 2929
rect 1602 2895 1614 2929
rect 1556 2862 1614 2895
rect 1686 2929 1744 2962
rect 1686 2895 1698 2929
rect 1732 2895 1744 2929
rect 1686 2862 1744 2895
rect 1844 2929 1902 2962
rect 1844 2895 1856 2929
rect 1890 2895 1902 2929
rect 1844 2862 1902 2895
rect 2018 2929 2076 2962
rect 2018 2895 2030 2929
rect 2064 2895 2076 2929
rect 2018 2862 2076 2895
rect 2176 2929 2234 2962
rect 2176 2895 2188 2929
rect 2222 2895 2234 2929
rect 2176 2862 2234 2895
rect 2360 2929 2418 2962
rect 2360 2895 2372 2929
rect 2406 2895 2418 2929
rect 2360 2862 2418 2895
rect 2518 2929 2576 2962
rect 2518 2895 2530 2929
rect 2564 2895 2576 2929
rect 2518 2862 2576 2895
rect 2764 2929 2822 2962
rect 2764 2895 2776 2929
rect 2810 2895 2822 2929
rect 2764 2862 2822 2895
rect 2922 2929 2980 2962
rect 2922 2895 2934 2929
rect 2968 2895 2980 2929
rect 2922 2862 2980 2895
rect 3108 2929 3166 2962
rect 3108 2895 3120 2929
rect 3154 2895 3166 2929
rect 3108 2862 3166 2895
rect 3266 2929 3324 2962
rect 3266 2895 3278 2929
rect 3312 2895 3324 2929
rect 3266 2862 3324 2895
rect 3730 2939 3788 2972
rect 3730 2905 3742 2939
rect 3776 2905 3788 2939
rect 3730 2872 3788 2905
rect 3888 2939 3946 2972
rect 3888 2905 3900 2939
rect 3934 2905 3946 2939
rect 3888 2872 3946 2905
rect 4038 2939 4096 2972
rect 4038 2905 4050 2939
rect 4084 2905 4096 2939
rect 4038 2872 4096 2905
rect 4196 2939 4254 2972
rect 4196 2905 4208 2939
rect 4242 2905 4254 2939
rect 4196 2872 4254 2905
rect 4390 2941 4448 2974
rect 4390 2907 4402 2941
rect 4436 2907 4448 2941
rect 4390 2874 4448 2907
rect 4548 2941 4606 2974
rect 4548 2907 4560 2941
rect 4594 2907 4606 2941
rect 4548 2874 4606 2907
rect 4698 2941 4756 2974
rect 4698 2907 4710 2941
rect 4744 2907 4756 2941
rect 4698 2874 4756 2907
rect 4856 2941 4914 2974
rect 4856 2907 4868 2941
rect 4902 2907 4914 2941
rect 4856 2874 4914 2907
rect 5688 2940 5746 2972
rect 5688 2906 5700 2940
rect 5734 2906 5746 2940
rect 5688 2872 5746 2906
rect 5846 2940 5904 2972
rect 5846 2906 5858 2940
rect 5892 2906 5904 2940
rect 5846 2872 5904 2906
rect 5996 2940 6054 2972
rect 5996 2906 6008 2940
rect 6042 2906 6054 2940
rect 5996 2872 6054 2906
rect 6154 2940 6212 2972
rect 6154 2906 6166 2940
rect 6200 2906 6212 2940
rect 6154 2872 6212 2906
rect 6348 2942 6406 2974
rect 6348 2908 6360 2942
rect 6394 2908 6406 2942
rect 6348 2874 6406 2908
rect 6506 2942 6564 2974
rect 6506 2908 6518 2942
rect 6552 2908 6564 2942
rect 6506 2874 6564 2908
rect 6656 2942 6714 2974
rect 6656 2908 6668 2942
rect 6702 2908 6714 2942
rect 6656 2874 6714 2908
rect 6814 2942 6872 2974
rect 6814 2908 6826 2942
rect 6860 2908 6872 2942
rect 6814 2874 6872 2908
rect 988 2788 1013 2822
rect 1047 2788 1072 2822
rect 988 2776 1072 2788
rect 544 2156 628 2168
rect 544 2122 569 2156
rect 603 2122 628 2156
rect 544 2065 628 2122
rect 544 1588 628 1645
rect 544 1554 569 1588
rect 603 1554 628 1588
rect 544 1542 628 1554
rect 690 2156 774 2168
rect 690 2122 715 2156
rect 749 2122 774 2156
rect 690 2065 774 2122
rect 690 1588 774 1645
rect 690 1554 715 1588
rect 749 1554 774 1588
rect 690 1542 774 1554
rect 834 2162 918 2174
rect 834 2128 859 2162
rect 893 2128 918 2162
rect 834 2071 918 2128
rect 834 1594 918 1651
rect 834 1560 859 1594
rect 893 1560 918 1594
rect 834 1548 918 1560
rect 988 2162 1072 2174
rect 988 2128 1013 2162
rect 1047 2128 1072 2162
rect 988 2071 1072 2128
rect 988 1594 1072 1651
rect 1398 1701 1456 1734
rect 1398 1667 1410 1701
rect 1444 1667 1456 1701
rect 1398 1634 1456 1667
rect 1556 1701 1614 1734
rect 1556 1667 1568 1701
rect 1602 1667 1614 1701
rect 1556 1634 1614 1667
rect 1686 1701 1744 1734
rect 1686 1667 1698 1701
rect 1732 1667 1744 1701
rect 1686 1634 1744 1667
rect 1844 1701 1902 1734
rect 1844 1667 1856 1701
rect 1890 1667 1902 1701
rect 1844 1634 1902 1667
rect 2018 1701 2076 1734
rect 2018 1667 2030 1701
rect 2064 1667 2076 1701
rect 2018 1634 2076 1667
rect 2176 1701 2234 1734
rect 2176 1667 2188 1701
rect 2222 1667 2234 1701
rect 2176 1634 2234 1667
rect 2360 1701 2418 1734
rect 2360 1667 2372 1701
rect 2406 1667 2418 1701
rect 2360 1634 2418 1667
rect 2518 1701 2576 1734
rect 2518 1667 2530 1701
rect 2564 1667 2576 1701
rect 2518 1634 2576 1667
rect 2764 1701 2822 1734
rect 2764 1667 2776 1701
rect 2810 1667 2822 1701
rect 2764 1634 2822 1667
rect 2922 1701 2980 1734
rect 2922 1667 2934 1701
rect 2968 1667 2980 1701
rect 2922 1634 2980 1667
rect 3108 1701 3166 1734
rect 3108 1667 3120 1701
rect 3154 1667 3166 1701
rect 3108 1634 3166 1667
rect 3266 1701 3324 1734
rect 3266 1667 3278 1701
rect 3312 1667 3324 1701
rect 3266 1634 3324 1667
rect 3730 1711 3788 1744
rect 3730 1677 3742 1711
rect 3776 1677 3788 1711
rect 3730 1644 3788 1677
rect 3888 1711 3946 1744
rect 3888 1677 3900 1711
rect 3934 1677 3946 1711
rect 3888 1644 3946 1677
rect 4038 1711 4096 1744
rect 4038 1677 4050 1711
rect 4084 1677 4096 1711
rect 4038 1644 4096 1677
rect 4196 1711 4254 1744
rect 4196 1677 4208 1711
rect 4242 1677 4254 1711
rect 4196 1644 4254 1677
rect 4390 1713 4448 1746
rect 4390 1679 4402 1713
rect 4436 1679 4448 1713
rect 4390 1646 4448 1679
rect 4548 1713 4606 1746
rect 4548 1679 4560 1713
rect 4594 1679 4606 1713
rect 4548 1646 4606 1679
rect 4698 1713 4756 1746
rect 4698 1679 4710 1713
rect 4744 1679 4756 1713
rect 4698 1646 4756 1679
rect 4856 1713 4914 1746
rect 4856 1679 4868 1713
rect 4902 1679 4914 1713
rect 4856 1646 4914 1679
rect 5688 1712 5746 1744
rect 5688 1678 5700 1712
rect 5734 1678 5746 1712
rect 5688 1644 5746 1678
rect 5846 1712 5904 1744
rect 5846 1678 5858 1712
rect 5892 1678 5904 1712
rect 5846 1644 5904 1678
rect 5996 1712 6054 1744
rect 5996 1678 6008 1712
rect 6042 1678 6054 1712
rect 5996 1644 6054 1678
rect 6154 1712 6212 1744
rect 6154 1678 6166 1712
rect 6200 1678 6212 1712
rect 6154 1644 6212 1678
rect 6348 1714 6406 1746
rect 6348 1680 6360 1714
rect 6394 1680 6406 1714
rect 6348 1646 6406 1680
rect 6506 1714 6564 1746
rect 6506 1680 6518 1714
rect 6552 1680 6564 1714
rect 6506 1646 6564 1680
rect 6656 1714 6714 1746
rect 6656 1680 6668 1714
rect 6702 1680 6714 1714
rect 6656 1646 6714 1680
rect 6814 1714 6872 1746
rect 6814 1680 6826 1714
rect 6860 1680 6872 1714
rect 6814 1646 6872 1680
rect 988 1560 1013 1594
rect 1047 1560 1072 1594
rect 988 1548 1072 1560
rect 544 928 628 940
rect 544 894 569 928
rect 603 894 628 928
rect 544 837 628 894
rect 544 360 628 417
rect 544 326 569 360
rect 603 326 628 360
rect 544 314 628 326
rect 690 928 774 940
rect 690 894 715 928
rect 749 894 774 928
rect 690 837 774 894
rect 690 360 774 417
rect 690 326 715 360
rect 749 326 774 360
rect 690 314 774 326
rect 834 934 918 946
rect 834 900 859 934
rect 893 900 918 934
rect 834 843 918 900
rect 834 366 918 423
rect 834 332 859 366
rect 893 332 918 366
rect 834 320 918 332
rect 988 934 1072 946
rect 988 900 1013 934
rect 1047 900 1072 934
rect 988 843 1072 900
rect 988 366 1072 423
rect 1398 473 1456 506
rect 1398 439 1410 473
rect 1444 439 1456 473
rect 1398 406 1456 439
rect 1556 473 1614 506
rect 1556 439 1568 473
rect 1602 439 1614 473
rect 1556 406 1614 439
rect 1686 473 1744 506
rect 1686 439 1698 473
rect 1732 439 1744 473
rect 1686 406 1744 439
rect 1844 473 1902 506
rect 1844 439 1856 473
rect 1890 439 1902 473
rect 1844 406 1902 439
rect 2018 473 2076 506
rect 2018 439 2030 473
rect 2064 439 2076 473
rect 2018 406 2076 439
rect 2176 473 2234 506
rect 2176 439 2188 473
rect 2222 439 2234 473
rect 2176 406 2234 439
rect 2360 473 2418 506
rect 2360 439 2372 473
rect 2406 439 2418 473
rect 2360 406 2418 439
rect 2518 473 2576 506
rect 2518 439 2530 473
rect 2564 439 2576 473
rect 2518 406 2576 439
rect 2764 473 2822 506
rect 2764 439 2776 473
rect 2810 439 2822 473
rect 2764 406 2822 439
rect 2922 473 2980 506
rect 2922 439 2934 473
rect 2968 439 2980 473
rect 2922 406 2980 439
rect 3108 473 3166 506
rect 3108 439 3120 473
rect 3154 439 3166 473
rect 3108 406 3166 439
rect 3266 473 3324 506
rect 3266 439 3278 473
rect 3312 439 3324 473
rect 3266 406 3324 439
rect 3730 483 3788 516
rect 3730 449 3742 483
rect 3776 449 3788 483
rect 3730 416 3788 449
rect 3888 483 3946 516
rect 3888 449 3900 483
rect 3934 449 3946 483
rect 3888 416 3946 449
rect 4038 483 4096 516
rect 4038 449 4050 483
rect 4084 449 4096 483
rect 4038 416 4096 449
rect 4196 483 4254 516
rect 4196 449 4208 483
rect 4242 449 4254 483
rect 4196 416 4254 449
rect 4390 485 4448 518
rect 4390 451 4402 485
rect 4436 451 4448 485
rect 4390 418 4448 451
rect 4548 485 4606 518
rect 4548 451 4560 485
rect 4594 451 4606 485
rect 4548 418 4606 451
rect 4698 485 4756 518
rect 4698 451 4710 485
rect 4744 451 4756 485
rect 4698 418 4756 451
rect 4856 485 4914 518
rect 4856 451 4868 485
rect 4902 451 4914 485
rect 4856 418 4914 451
rect 988 332 1013 366
rect 1047 332 1072 366
rect 988 320 1072 332
<< mvpdiff >>
rect 1398 19249 1456 19264
rect 1398 19215 1410 19249
rect 1444 19215 1456 19249
rect 1398 19181 1456 19215
rect 1398 19147 1410 19181
rect 1444 19147 1456 19181
rect 1398 19113 1456 19147
rect 1398 19079 1410 19113
rect 1444 19079 1456 19113
rect 1398 19064 1456 19079
rect 1556 19249 1614 19264
rect 1556 19215 1568 19249
rect 1602 19215 1614 19249
rect 1556 19181 1614 19215
rect 1556 19147 1568 19181
rect 1602 19147 1614 19181
rect 1556 19113 1614 19147
rect 1556 19079 1568 19113
rect 1602 19079 1614 19113
rect 1556 19064 1614 19079
rect 1686 19249 1744 19264
rect 1686 19215 1698 19249
rect 1732 19215 1744 19249
rect 1686 19181 1744 19215
rect 1686 19147 1698 19181
rect 1732 19147 1744 19181
rect 1686 19113 1744 19147
rect 1686 19079 1698 19113
rect 1732 19079 1744 19113
rect 1686 19064 1744 19079
rect 1844 19249 1902 19264
rect 1844 19215 1856 19249
rect 1890 19215 1902 19249
rect 1844 19181 1902 19215
rect 1844 19147 1856 19181
rect 1890 19147 1902 19181
rect 1844 19113 1902 19147
rect 1844 19079 1856 19113
rect 1890 19079 1902 19113
rect 1844 19064 1902 19079
rect 2018 19249 2076 19264
rect 2018 19215 2030 19249
rect 2064 19215 2076 19249
rect 2018 19181 2076 19215
rect 2018 19147 2030 19181
rect 2064 19147 2076 19181
rect 2018 19113 2076 19147
rect 2018 19079 2030 19113
rect 2064 19079 2076 19113
rect 2018 19064 2076 19079
rect 2176 19249 2234 19264
rect 2176 19215 2188 19249
rect 2222 19215 2234 19249
rect 2176 19181 2234 19215
rect 2176 19147 2188 19181
rect 2222 19147 2234 19181
rect 2176 19113 2234 19147
rect 2176 19079 2188 19113
rect 2222 19079 2234 19113
rect 2176 19064 2234 19079
rect 2360 19249 2418 19264
rect 2360 19215 2372 19249
rect 2406 19215 2418 19249
rect 2360 19181 2418 19215
rect 2360 19147 2372 19181
rect 2406 19147 2418 19181
rect 2360 19113 2418 19147
rect 2360 19079 2372 19113
rect 2406 19079 2418 19113
rect 2360 19064 2418 19079
rect 2518 19249 2576 19264
rect 2518 19215 2530 19249
rect 2564 19215 2576 19249
rect 2518 19181 2576 19215
rect 2518 19147 2530 19181
rect 2564 19147 2576 19181
rect 2518 19113 2576 19147
rect 2518 19079 2530 19113
rect 2564 19079 2576 19113
rect 2518 19064 2576 19079
rect 2764 19249 2822 19264
rect 2764 19215 2776 19249
rect 2810 19215 2822 19249
rect 2764 19181 2822 19215
rect 2764 19147 2776 19181
rect 2810 19147 2822 19181
rect 2764 19113 2822 19147
rect 2764 19079 2776 19113
rect 2810 19079 2822 19113
rect 2764 19064 2822 19079
rect 2922 19249 2980 19264
rect 2922 19215 2934 19249
rect 2968 19215 2980 19249
rect 2922 19181 2980 19215
rect 2922 19147 2934 19181
rect 2968 19147 2980 19181
rect 2922 19113 2980 19147
rect 2922 19079 2934 19113
rect 2968 19079 2980 19113
rect 2922 19064 2980 19079
rect 3108 19249 3166 19264
rect 3108 19215 3120 19249
rect 3154 19215 3166 19249
rect 3108 19181 3166 19215
rect 3108 19147 3120 19181
rect 3154 19147 3166 19181
rect 3108 19113 3166 19147
rect 3108 19079 3120 19113
rect 3154 19079 3166 19113
rect 3108 19064 3166 19079
rect 3266 19249 3324 19264
rect 3266 19215 3278 19249
rect 3312 19215 3324 19249
rect 3266 19181 3324 19215
rect 3266 19147 3278 19181
rect 3312 19147 3324 19181
rect 3266 19113 3324 19147
rect 3266 19079 3278 19113
rect 3312 19079 3324 19113
rect 3266 19064 3324 19079
rect 3730 19259 3788 19274
rect 3730 19225 3742 19259
rect 3776 19225 3788 19259
rect 3730 19191 3788 19225
rect 3730 19157 3742 19191
rect 3776 19157 3788 19191
rect 3730 19123 3788 19157
rect 3730 19089 3742 19123
rect 3776 19089 3788 19123
rect 3730 19074 3788 19089
rect 3888 19259 3946 19274
rect 3888 19225 3900 19259
rect 3934 19225 3946 19259
rect 3888 19191 3946 19225
rect 3888 19157 3900 19191
rect 3934 19157 3946 19191
rect 3888 19123 3946 19157
rect 3888 19089 3900 19123
rect 3934 19089 3946 19123
rect 3888 19074 3946 19089
rect 4038 19259 4096 19274
rect 4038 19225 4050 19259
rect 4084 19225 4096 19259
rect 4038 19191 4096 19225
rect 4038 19157 4050 19191
rect 4084 19157 4096 19191
rect 4038 19123 4096 19157
rect 4038 19089 4050 19123
rect 4084 19089 4096 19123
rect 4038 19074 4096 19089
rect 4196 19259 4254 19274
rect 4196 19225 4208 19259
rect 4242 19225 4254 19259
rect 4196 19191 4254 19225
rect 4196 19157 4208 19191
rect 4242 19157 4254 19191
rect 4196 19123 4254 19157
rect 4196 19089 4208 19123
rect 4242 19089 4254 19123
rect 4196 19074 4254 19089
rect 4390 19259 4448 19274
rect 4390 19225 4402 19259
rect 4436 19225 4448 19259
rect 4390 19191 4448 19225
rect 4390 19157 4402 19191
rect 4436 19157 4448 19191
rect 4390 19123 4448 19157
rect 4390 19089 4402 19123
rect 4436 19089 4448 19123
rect 4390 19074 4448 19089
rect 4548 19259 4606 19274
rect 4548 19225 4560 19259
rect 4594 19225 4606 19259
rect 4548 19191 4606 19225
rect 4548 19157 4560 19191
rect 4594 19157 4606 19191
rect 4548 19123 4606 19157
rect 4548 19089 4560 19123
rect 4594 19089 4606 19123
rect 4548 19074 4606 19089
rect 4698 19259 4756 19274
rect 4698 19225 4710 19259
rect 4744 19225 4756 19259
rect 4698 19191 4756 19225
rect 4698 19157 4710 19191
rect 4744 19157 4756 19191
rect 4698 19123 4756 19157
rect 4698 19089 4710 19123
rect 4744 19089 4756 19123
rect 4698 19074 4756 19089
rect 4856 19259 4914 19274
rect 4856 19225 4868 19259
rect 4902 19225 4914 19259
rect 4856 19191 4914 19225
rect 4856 19157 4868 19191
rect 4902 19157 4914 19191
rect 4856 19123 4914 19157
rect 4856 19089 4868 19123
rect 4902 19089 4914 19123
rect 4856 19074 4914 19089
rect 5688 19260 5746 19274
rect 5688 19226 5700 19260
rect 5734 19226 5746 19260
rect 5688 19192 5746 19226
rect 5688 19158 5700 19192
rect 5734 19158 5746 19192
rect 5688 19124 5746 19158
rect 5688 19090 5700 19124
rect 5734 19090 5746 19124
rect 5688 19074 5746 19090
rect 5846 19260 5904 19274
rect 5846 19226 5858 19260
rect 5892 19226 5904 19260
rect 5846 19192 5904 19226
rect 5846 19158 5858 19192
rect 5892 19158 5904 19192
rect 5846 19124 5904 19158
rect 5846 19090 5858 19124
rect 5892 19090 5904 19124
rect 5846 19074 5904 19090
rect 5996 19260 6054 19274
rect 5996 19226 6008 19260
rect 6042 19226 6054 19260
rect 5996 19192 6054 19226
rect 5996 19158 6008 19192
rect 6042 19158 6054 19192
rect 5996 19124 6054 19158
rect 5996 19090 6008 19124
rect 6042 19090 6054 19124
rect 5996 19074 6054 19090
rect 6154 19260 6212 19274
rect 6154 19226 6166 19260
rect 6200 19226 6212 19260
rect 6154 19192 6212 19226
rect 6154 19158 6166 19192
rect 6200 19158 6212 19192
rect 6154 19124 6212 19158
rect 6154 19090 6166 19124
rect 6200 19090 6212 19124
rect 6154 19074 6212 19090
rect 6348 19260 6406 19274
rect 6348 19226 6360 19260
rect 6394 19226 6406 19260
rect 6348 19192 6406 19226
rect 6348 19158 6360 19192
rect 6394 19158 6406 19192
rect 6348 19124 6406 19158
rect 6348 19090 6360 19124
rect 6394 19090 6406 19124
rect 6348 19074 6406 19090
rect 6506 19260 6564 19274
rect 6506 19226 6518 19260
rect 6552 19226 6564 19260
rect 6506 19192 6564 19226
rect 6506 19158 6518 19192
rect 6552 19158 6564 19192
rect 6506 19124 6564 19158
rect 6506 19090 6518 19124
rect 6552 19090 6564 19124
rect 6506 19074 6564 19090
rect 6656 19260 6714 19274
rect 6656 19226 6668 19260
rect 6702 19226 6714 19260
rect 6656 19192 6714 19226
rect 6656 19158 6668 19192
rect 6702 19158 6714 19192
rect 6656 19124 6714 19158
rect 6656 19090 6668 19124
rect 6702 19090 6714 19124
rect 6656 19074 6714 19090
rect 6814 19260 6872 19274
rect 6814 19226 6826 19260
rect 6860 19226 6872 19260
rect 6814 19192 6872 19226
rect 6814 19158 6826 19192
rect 6860 19158 6872 19192
rect 6814 19124 6872 19158
rect 6814 19090 6826 19124
rect 6860 19090 6872 19124
rect 6814 19074 6872 19090
rect 1398 18021 1456 18036
rect 1398 17987 1410 18021
rect 1444 17987 1456 18021
rect 1398 17953 1456 17987
rect 1398 17919 1410 17953
rect 1444 17919 1456 17953
rect 1398 17885 1456 17919
rect 1398 17851 1410 17885
rect 1444 17851 1456 17885
rect 1398 17836 1456 17851
rect 1556 18021 1614 18036
rect 1556 17987 1568 18021
rect 1602 17987 1614 18021
rect 1556 17953 1614 17987
rect 1556 17919 1568 17953
rect 1602 17919 1614 17953
rect 1556 17885 1614 17919
rect 1556 17851 1568 17885
rect 1602 17851 1614 17885
rect 1556 17836 1614 17851
rect 1686 18021 1744 18036
rect 1686 17987 1698 18021
rect 1732 17987 1744 18021
rect 1686 17953 1744 17987
rect 1686 17919 1698 17953
rect 1732 17919 1744 17953
rect 1686 17885 1744 17919
rect 1686 17851 1698 17885
rect 1732 17851 1744 17885
rect 1686 17836 1744 17851
rect 1844 18021 1902 18036
rect 1844 17987 1856 18021
rect 1890 17987 1902 18021
rect 1844 17953 1902 17987
rect 1844 17919 1856 17953
rect 1890 17919 1902 17953
rect 1844 17885 1902 17919
rect 1844 17851 1856 17885
rect 1890 17851 1902 17885
rect 1844 17836 1902 17851
rect 2018 18021 2076 18036
rect 2018 17987 2030 18021
rect 2064 17987 2076 18021
rect 2018 17953 2076 17987
rect 2018 17919 2030 17953
rect 2064 17919 2076 17953
rect 2018 17885 2076 17919
rect 2018 17851 2030 17885
rect 2064 17851 2076 17885
rect 2018 17836 2076 17851
rect 2176 18021 2234 18036
rect 2176 17987 2188 18021
rect 2222 17987 2234 18021
rect 2176 17953 2234 17987
rect 2176 17919 2188 17953
rect 2222 17919 2234 17953
rect 2176 17885 2234 17919
rect 2176 17851 2188 17885
rect 2222 17851 2234 17885
rect 2176 17836 2234 17851
rect 2360 18021 2418 18036
rect 2360 17987 2372 18021
rect 2406 17987 2418 18021
rect 2360 17953 2418 17987
rect 2360 17919 2372 17953
rect 2406 17919 2418 17953
rect 2360 17885 2418 17919
rect 2360 17851 2372 17885
rect 2406 17851 2418 17885
rect 2360 17836 2418 17851
rect 2518 18021 2576 18036
rect 2518 17987 2530 18021
rect 2564 17987 2576 18021
rect 2518 17953 2576 17987
rect 2518 17919 2530 17953
rect 2564 17919 2576 17953
rect 2518 17885 2576 17919
rect 2518 17851 2530 17885
rect 2564 17851 2576 17885
rect 2518 17836 2576 17851
rect 2764 18021 2822 18036
rect 2764 17987 2776 18021
rect 2810 17987 2822 18021
rect 2764 17953 2822 17987
rect 2764 17919 2776 17953
rect 2810 17919 2822 17953
rect 2764 17885 2822 17919
rect 2764 17851 2776 17885
rect 2810 17851 2822 17885
rect 2764 17836 2822 17851
rect 2922 18021 2980 18036
rect 2922 17987 2934 18021
rect 2968 17987 2980 18021
rect 2922 17953 2980 17987
rect 2922 17919 2934 17953
rect 2968 17919 2980 17953
rect 2922 17885 2980 17919
rect 2922 17851 2934 17885
rect 2968 17851 2980 17885
rect 2922 17836 2980 17851
rect 3108 18021 3166 18036
rect 3108 17987 3120 18021
rect 3154 17987 3166 18021
rect 3108 17953 3166 17987
rect 3108 17919 3120 17953
rect 3154 17919 3166 17953
rect 3108 17885 3166 17919
rect 3108 17851 3120 17885
rect 3154 17851 3166 17885
rect 3108 17836 3166 17851
rect 3266 18021 3324 18036
rect 3266 17987 3278 18021
rect 3312 17987 3324 18021
rect 3266 17953 3324 17987
rect 3266 17919 3278 17953
rect 3312 17919 3324 17953
rect 3266 17885 3324 17919
rect 3266 17851 3278 17885
rect 3312 17851 3324 17885
rect 3266 17836 3324 17851
rect 3730 18031 3788 18046
rect 3730 17997 3742 18031
rect 3776 17997 3788 18031
rect 3730 17963 3788 17997
rect 3730 17929 3742 17963
rect 3776 17929 3788 17963
rect 3730 17895 3788 17929
rect 3730 17861 3742 17895
rect 3776 17861 3788 17895
rect 3730 17846 3788 17861
rect 3888 18031 3946 18046
rect 3888 17997 3900 18031
rect 3934 17997 3946 18031
rect 3888 17963 3946 17997
rect 3888 17929 3900 17963
rect 3934 17929 3946 17963
rect 3888 17895 3946 17929
rect 3888 17861 3900 17895
rect 3934 17861 3946 17895
rect 3888 17846 3946 17861
rect 4038 18031 4096 18046
rect 4038 17997 4050 18031
rect 4084 17997 4096 18031
rect 4038 17963 4096 17997
rect 4038 17929 4050 17963
rect 4084 17929 4096 17963
rect 4038 17895 4096 17929
rect 4038 17861 4050 17895
rect 4084 17861 4096 17895
rect 4038 17846 4096 17861
rect 4196 18031 4254 18046
rect 4196 17997 4208 18031
rect 4242 17997 4254 18031
rect 4196 17963 4254 17997
rect 4196 17929 4208 17963
rect 4242 17929 4254 17963
rect 4196 17895 4254 17929
rect 4196 17861 4208 17895
rect 4242 17861 4254 17895
rect 4196 17846 4254 17861
rect 4390 18031 4448 18046
rect 4390 17997 4402 18031
rect 4436 17997 4448 18031
rect 4390 17963 4448 17997
rect 4390 17929 4402 17963
rect 4436 17929 4448 17963
rect 4390 17895 4448 17929
rect 4390 17861 4402 17895
rect 4436 17861 4448 17895
rect 4390 17846 4448 17861
rect 4548 18031 4606 18046
rect 4548 17997 4560 18031
rect 4594 17997 4606 18031
rect 4548 17963 4606 17997
rect 4548 17929 4560 17963
rect 4594 17929 4606 17963
rect 4548 17895 4606 17929
rect 4548 17861 4560 17895
rect 4594 17861 4606 17895
rect 4548 17846 4606 17861
rect 4698 18031 4756 18046
rect 4698 17997 4710 18031
rect 4744 17997 4756 18031
rect 4698 17963 4756 17997
rect 4698 17929 4710 17963
rect 4744 17929 4756 17963
rect 4698 17895 4756 17929
rect 4698 17861 4710 17895
rect 4744 17861 4756 17895
rect 4698 17846 4756 17861
rect 4856 18031 4914 18046
rect 4856 17997 4868 18031
rect 4902 17997 4914 18031
rect 4856 17963 4914 17997
rect 4856 17929 4868 17963
rect 4902 17929 4914 17963
rect 4856 17895 4914 17929
rect 4856 17861 4868 17895
rect 4902 17861 4914 17895
rect 4856 17846 4914 17861
rect 5688 18032 5746 18046
rect 5688 17998 5700 18032
rect 5734 17998 5746 18032
rect 5688 17964 5746 17998
rect 5688 17930 5700 17964
rect 5734 17930 5746 17964
rect 5688 17896 5746 17930
rect 5688 17862 5700 17896
rect 5734 17862 5746 17896
rect 5688 17846 5746 17862
rect 5846 18032 5904 18046
rect 5846 17998 5858 18032
rect 5892 17998 5904 18032
rect 5846 17964 5904 17998
rect 5846 17930 5858 17964
rect 5892 17930 5904 17964
rect 5846 17896 5904 17930
rect 5846 17862 5858 17896
rect 5892 17862 5904 17896
rect 5846 17846 5904 17862
rect 5996 18032 6054 18046
rect 5996 17998 6008 18032
rect 6042 17998 6054 18032
rect 5996 17964 6054 17998
rect 5996 17930 6008 17964
rect 6042 17930 6054 17964
rect 5996 17896 6054 17930
rect 5996 17862 6008 17896
rect 6042 17862 6054 17896
rect 5996 17846 6054 17862
rect 6154 18032 6212 18046
rect 6154 17998 6166 18032
rect 6200 17998 6212 18032
rect 6154 17964 6212 17998
rect 6154 17930 6166 17964
rect 6200 17930 6212 17964
rect 6154 17896 6212 17930
rect 6154 17862 6166 17896
rect 6200 17862 6212 17896
rect 6154 17846 6212 17862
rect 6348 18032 6406 18046
rect 6348 17998 6360 18032
rect 6394 17998 6406 18032
rect 6348 17964 6406 17998
rect 6348 17930 6360 17964
rect 6394 17930 6406 17964
rect 6348 17896 6406 17930
rect 6348 17862 6360 17896
rect 6394 17862 6406 17896
rect 6348 17846 6406 17862
rect 6506 18032 6564 18046
rect 6506 17998 6518 18032
rect 6552 17998 6564 18032
rect 6506 17964 6564 17998
rect 6506 17930 6518 17964
rect 6552 17930 6564 17964
rect 6506 17896 6564 17930
rect 6506 17862 6518 17896
rect 6552 17862 6564 17896
rect 6506 17846 6564 17862
rect 6656 18032 6714 18046
rect 6656 17998 6668 18032
rect 6702 17998 6714 18032
rect 6656 17964 6714 17998
rect 6656 17930 6668 17964
rect 6702 17930 6714 17964
rect 6656 17896 6714 17930
rect 6656 17862 6668 17896
rect 6702 17862 6714 17896
rect 6656 17846 6714 17862
rect 6814 18032 6872 18046
rect 6814 17998 6826 18032
rect 6860 17998 6872 18032
rect 6814 17964 6872 17998
rect 6814 17930 6826 17964
rect 6860 17930 6872 17964
rect 6814 17896 6872 17930
rect 6814 17862 6826 17896
rect 6860 17862 6872 17896
rect 6814 17846 6872 17862
rect 1398 16793 1456 16808
rect 1398 16759 1410 16793
rect 1444 16759 1456 16793
rect 1398 16725 1456 16759
rect 1398 16691 1410 16725
rect 1444 16691 1456 16725
rect 1398 16657 1456 16691
rect 1398 16623 1410 16657
rect 1444 16623 1456 16657
rect 1398 16608 1456 16623
rect 1556 16793 1614 16808
rect 1556 16759 1568 16793
rect 1602 16759 1614 16793
rect 1556 16725 1614 16759
rect 1556 16691 1568 16725
rect 1602 16691 1614 16725
rect 1556 16657 1614 16691
rect 1556 16623 1568 16657
rect 1602 16623 1614 16657
rect 1556 16608 1614 16623
rect 1686 16793 1744 16808
rect 1686 16759 1698 16793
rect 1732 16759 1744 16793
rect 1686 16725 1744 16759
rect 1686 16691 1698 16725
rect 1732 16691 1744 16725
rect 1686 16657 1744 16691
rect 1686 16623 1698 16657
rect 1732 16623 1744 16657
rect 1686 16608 1744 16623
rect 1844 16793 1902 16808
rect 1844 16759 1856 16793
rect 1890 16759 1902 16793
rect 1844 16725 1902 16759
rect 1844 16691 1856 16725
rect 1890 16691 1902 16725
rect 1844 16657 1902 16691
rect 1844 16623 1856 16657
rect 1890 16623 1902 16657
rect 1844 16608 1902 16623
rect 2018 16793 2076 16808
rect 2018 16759 2030 16793
rect 2064 16759 2076 16793
rect 2018 16725 2076 16759
rect 2018 16691 2030 16725
rect 2064 16691 2076 16725
rect 2018 16657 2076 16691
rect 2018 16623 2030 16657
rect 2064 16623 2076 16657
rect 2018 16608 2076 16623
rect 2176 16793 2234 16808
rect 2176 16759 2188 16793
rect 2222 16759 2234 16793
rect 2176 16725 2234 16759
rect 2176 16691 2188 16725
rect 2222 16691 2234 16725
rect 2176 16657 2234 16691
rect 2176 16623 2188 16657
rect 2222 16623 2234 16657
rect 2176 16608 2234 16623
rect 2360 16793 2418 16808
rect 2360 16759 2372 16793
rect 2406 16759 2418 16793
rect 2360 16725 2418 16759
rect 2360 16691 2372 16725
rect 2406 16691 2418 16725
rect 2360 16657 2418 16691
rect 2360 16623 2372 16657
rect 2406 16623 2418 16657
rect 2360 16608 2418 16623
rect 2518 16793 2576 16808
rect 2518 16759 2530 16793
rect 2564 16759 2576 16793
rect 2518 16725 2576 16759
rect 2518 16691 2530 16725
rect 2564 16691 2576 16725
rect 2518 16657 2576 16691
rect 2518 16623 2530 16657
rect 2564 16623 2576 16657
rect 2518 16608 2576 16623
rect 2764 16793 2822 16808
rect 2764 16759 2776 16793
rect 2810 16759 2822 16793
rect 2764 16725 2822 16759
rect 2764 16691 2776 16725
rect 2810 16691 2822 16725
rect 2764 16657 2822 16691
rect 2764 16623 2776 16657
rect 2810 16623 2822 16657
rect 2764 16608 2822 16623
rect 2922 16793 2980 16808
rect 2922 16759 2934 16793
rect 2968 16759 2980 16793
rect 2922 16725 2980 16759
rect 2922 16691 2934 16725
rect 2968 16691 2980 16725
rect 2922 16657 2980 16691
rect 2922 16623 2934 16657
rect 2968 16623 2980 16657
rect 2922 16608 2980 16623
rect 3108 16793 3166 16808
rect 3108 16759 3120 16793
rect 3154 16759 3166 16793
rect 3108 16725 3166 16759
rect 3108 16691 3120 16725
rect 3154 16691 3166 16725
rect 3108 16657 3166 16691
rect 3108 16623 3120 16657
rect 3154 16623 3166 16657
rect 3108 16608 3166 16623
rect 3266 16793 3324 16808
rect 3266 16759 3278 16793
rect 3312 16759 3324 16793
rect 3266 16725 3324 16759
rect 3266 16691 3278 16725
rect 3312 16691 3324 16725
rect 3266 16657 3324 16691
rect 3266 16623 3278 16657
rect 3312 16623 3324 16657
rect 3266 16608 3324 16623
rect 3730 16803 3788 16818
rect 3730 16769 3742 16803
rect 3776 16769 3788 16803
rect 3730 16735 3788 16769
rect 3730 16701 3742 16735
rect 3776 16701 3788 16735
rect 3730 16667 3788 16701
rect 3730 16633 3742 16667
rect 3776 16633 3788 16667
rect 3730 16618 3788 16633
rect 3888 16803 3946 16818
rect 3888 16769 3900 16803
rect 3934 16769 3946 16803
rect 3888 16735 3946 16769
rect 3888 16701 3900 16735
rect 3934 16701 3946 16735
rect 3888 16667 3946 16701
rect 3888 16633 3900 16667
rect 3934 16633 3946 16667
rect 3888 16618 3946 16633
rect 4038 16803 4096 16818
rect 4038 16769 4050 16803
rect 4084 16769 4096 16803
rect 4038 16735 4096 16769
rect 4038 16701 4050 16735
rect 4084 16701 4096 16735
rect 4038 16667 4096 16701
rect 4038 16633 4050 16667
rect 4084 16633 4096 16667
rect 4038 16618 4096 16633
rect 4196 16803 4254 16818
rect 4196 16769 4208 16803
rect 4242 16769 4254 16803
rect 4196 16735 4254 16769
rect 4196 16701 4208 16735
rect 4242 16701 4254 16735
rect 4196 16667 4254 16701
rect 4196 16633 4208 16667
rect 4242 16633 4254 16667
rect 4196 16618 4254 16633
rect 4390 16803 4448 16818
rect 4390 16769 4402 16803
rect 4436 16769 4448 16803
rect 4390 16735 4448 16769
rect 4390 16701 4402 16735
rect 4436 16701 4448 16735
rect 4390 16667 4448 16701
rect 4390 16633 4402 16667
rect 4436 16633 4448 16667
rect 4390 16618 4448 16633
rect 4548 16803 4606 16818
rect 4548 16769 4560 16803
rect 4594 16769 4606 16803
rect 4548 16735 4606 16769
rect 4548 16701 4560 16735
rect 4594 16701 4606 16735
rect 4548 16667 4606 16701
rect 4548 16633 4560 16667
rect 4594 16633 4606 16667
rect 4548 16618 4606 16633
rect 4698 16803 4756 16818
rect 4698 16769 4710 16803
rect 4744 16769 4756 16803
rect 4698 16735 4756 16769
rect 4698 16701 4710 16735
rect 4744 16701 4756 16735
rect 4698 16667 4756 16701
rect 4698 16633 4710 16667
rect 4744 16633 4756 16667
rect 4698 16618 4756 16633
rect 4856 16803 4914 16818
rect 4856 16769 4868 16803
rect 4902 16769 4914 16803
rect 4856 16735 4914 16769
rect 4856 16701 4868 16735
rect 4902 16701 4914 16735
rect 4856 16667 4914 16701
rect 4856 16633 4868 16667
rect 4902 16633 4914 16667
rect 4856 16618 4914 16633
rect 5688 16804 5746 16818
rect 5688 16770 5700 16804
rect 5734 16770 5746 16804
rect 5688 16736 5746 16770
rect 5688 16702 5700 16736
rect 5734 16702 5746 16736
rect 5688 16668 5746 16702
rect 5688 16634 5700 16668
rect 5734 16634 5746 16668
rect 5688 16618 5746 16634
rect 5846 16804 5904 16818
rect 5846 16770 5858 16804
rect 5892 16770 5904 16804
rect 5846 16736 5904 16770
rect 5846 16702 5858 16736
rect 5892 16702 5904 16736
rect 5846 16668 5904 16702
rect 5846 16634 5858 16668
rect 5892 16634 5904 16668
rect 5846 16618 5904 16634
rect 5996 16804 6054 16818
rect 5996 16770 6008 16804
rect 6042 16770 6054 16804
rect 5996 16736 6054 16770
rect 5996 16702 6008 16736
rect 6042 16702 6054 16736
rect 5996 16668 6054 16702
rect 5996 16634 6008 16668
rect 6042 16634 6054 16668
rect 5996 16618 6054 16634
rect 6154 16804 6212 16818
rect 6154 16770 6166 16804
rect 6200 16770 6212 16804
rect 6154 16736 6212 16770
rect 6154 16702 6166 16736
rect 6200 16702 6212 16736
rect 6154 16668 6212 16702
rect 6154 16634 6166 16668
rect 6200 16634 6212 16668
rect 6154 16618 6212 16634
rect 6348 16804 6406 16818
rect 6348 16770 6360 16804
rect 6394 16770 6406 16804
rect 6348 16736 6406 16770
rect 6348 16702 6360 16736
rect 6394 16702 6406 16736
rect 6348 16668 6406 16702
rect 6348 16634 6360 16668
rect 6394 16634 6406 16668
rect 6348 16618 6406 16634
rect 6506 16804 6564 16818
rect 6506 16770 6518 16804
rect 6552 16770 6564 16804
rect 6506 16736 6564 16770
rect 6506 16702 6518 16736
rect 6552 16702 6564 16736
rect 6506 16668 6564 16702
rect 6506 16634 6518 16668
rect 6552 16634 6564 16668
rect 6506 16618 6564 16634
rect 6656 16804 6714 16818
rect 6656 16770 6668 16804
rect 6702 16770 6714 16804
rect 6656 16736 6714 16770
rect 6656 16702 6668 16736
rect 6702 16702 6714 16736
rect 6656 16668 6714 16702
rect 6656 16634 6668 16668
rect 6702 16634 6714 16668
rect 6656 16618 6714 16634
rect 6814 16804 6872 16818
rect 6814 16770 6826 16804
rect 6860 16770 6872 16804
rect 6814 16736 6872 16770
rect 6814 16702 6826 16736
rect 6860 16702 6872 16736
rect 6814 16668 6872 16702
rect 6814 16634 6826 16668
rect 6860 16634 6872 16668
rect 6814 16618 6872 16634
rect 1398 15565 1456 15580
rect 1398 15531 1410 15565
rect 1444 15531 1456 15565
rect 1398 15497 1456 15531
rect 1398 15463 1410 15497
rect 1444 15463 1456 15497
rect 1398 15429 1456 15463
rect 1398 15395 1410 15429
rect 1444 15395 1456 15429
rect 1398 15380 1456 15395
rect 1556 15565 1614 15580
rect 1556 15531 1568 15565
rect 1602 15531 1614 15565
rect 1556 15497 1614 15531
rect 1556 15463 1568 15497
rect 1602 15463 1614 15497
rect 1556 15429 1614 15463
rect 1556 15395 1568 15429
rect 1602 15395 1614 15429
rect 1556 15380 1614 15395
rect 1686 15565 1744 15580
rect 1686 15531 1698 15565
rect 1732 15531 1744 15565
rect 1686 15497 1744 15531
rect 1686 15463 1698 15497
rect 1732 15463 1744 15497
rect 1686 15429 1744 15463
rect 1686 15395 1698 15429
rect 1732 15395 1744 15429
rect 1686 15380 1744 15395
rect 1844 15565 1902 15580
rect 1844 15531 1856 15565
rect 1890 15531 1902 15565
rect 1844 15497 1902 15531
rect 1844 15463 1856 15497
rect 1890 15463 1902 15497
rect 1844 15429 1902 15463
rect 1844 15395 1856 15429
rect 1890 15395 1902 15429
rect 1844 15380 1902 15395
rect 2018 15565 2076 15580
rect 2018 15531 2030 15565
rect 2064 15531 2076 15565
rect 2018 15497 2076 15531
rect 2018 15463 2030 15497
rect 2064 15463 2076 15497
rect 2018 15429 2076 15463
rect 2018 15395 2030 15429
rect 2064 15395 2076 15429
rect 2018 15380 2076 15395
rect 2176 15565 2234 15580
rect 2176 15531 2188 15565
rect 2222 15531 2234 15565
rect 2176 15497 2234 15531
rect 2176 15463 2188 15497
rect 2222 15463 2234 15497
rect 2176 15429 2234 15463
rect 2176 15395 2188 15429
rect 2222 15395 2234 15429
rect 2176 15380 2234 15395
rect 2360 15565 2418 15580
rect 2360 15531 2372 15565
rect 2406 15531 2418 15565
rect 2360 15497 2418 15531
rect 2360 15463 2372 15497
rect 2406 15463 2418 15497
rect 2360 15429 2418 15463
rect 2360 15395 2372 15429
rect 2406 15395 2418 15429
rect 2360 15380 2418 15395
rect 2518 15565 2576 15580
rect 2518 15531 2530 15565
rect 2564 15531 2576 15565
rect 2518 15497 2576 15531
rect 2518 15463 2530 15497
rect 2564 15463 2576 15497
rect 2518 15429 2576 15463
rect 2518 15395 2530 15429
rect 2564 15395 2576 15429
rect 2518 15380 2576 15395
rect 2764 15565 2822 15580
rect 2764 15531 2776 15565
rect 2810 15531 2822 15565
rect 2764 15497 2822 15531
rect 2764 15463 2776 15497
rect 2810 15463 2822 15497
rect 2764 15429 2822 15463
rect 2764 15395 2776 15429
rect 2810 15395 2822 15429
rect 2764 15380 2822 15395
rect 2922 15565 2980 15580
rect 2922 15531 2934 15565
rect 2968 15531 2980 15565
rect 2922 15497 2980 15531
rect 2922 15463 2934 15497
rect 2968 15463 2980 15497
rect 2922 15429 2980 15463
rect 2922 15395 2934 15429
rect 2968 15395 2980 15429
rect 2922 15380 2980 15395
rect 3108 15565 3166 15580
rect 3108 15531 3120 15565
rect 3154 15531 3166 15565
rect 3108 15497 3166 15531
rect 3108 15463 3120 15497
rect 3154 15463 3166 15497
rect 3108 15429 3166 15463
rect 3108 15395 3120 15429
rect 3154 15395 3166 15429
rect 3108 15380 3166 15395
rect 3266 15565 3324 15580
rect 3266 15531 3278 15565
rect 3312 15531 3324 15565
rect 3266 15497 3324 15531
rect 3266 15463 3278 15497
rect 3312 15463 3324 15497
rect 3266 15429 3324 15463
rect 3266 15395 3278 15429
rect 3312 15395 3324 15429
rect 3266 15380 3324 15395
rect 3730 15575 3788 15590
rect 3730 15541 3742 15575
rect 3776 15541 3788 15575
rect 3730 15507 3788 15541
rect 3730 15473 3742 15507
rect 3776 15473 3788 15507
rect 3730 15439 3788 15473
rect 3730 15405 3742 15439
rect 3776 15405 3788 15439
rect 3730 15390 3788 15405
rect 3888 15575 3946 15590
rect 3888 15541 3900 15575
rect 3934 15541 3946 15575
rect 3888 15507 3946 15541
rect 3888 15473 3900 15507
rect 3934 15473 3946 15507
rect 3888 15439 3946 15473
rect 3888 15405 3900 15439
rect 3934 15405 3946 15439
rect 3888 15390 3946 15405
rect 4038 15575 4096 15590
rect 4038 15541 4050 15575
rect 4084 15541 4096 15575
rect 4038 15507 4096 15541
rect 4038 15473 4050 15507
rect 4084 15473 4096 15507
rect 4038 15439 4096 15473
rect 4038 15405 4050 15439
rect 4084 15405 4096 15439
rect 4038 15390 4096 15405
rect 4196 15575 4254 15590
rect 4196 15541 4208 15575
rect 4242 15541 4254 15575
rect 4196 15507 4254 15541
rect 4196 15473 4208 15507
rect 4242 15473 4254 15507
rect 4196 15439 4254 15473
rect 4196 15405 4208 15439
rect 4242 15405 4254 15439
rect 4196 15390 4254 15405
rect 4390 15575 4448 15590
rect 4390 15541 4402 15575
rect 4436 15541 4448 15575
rect 4390 15507 4448 15541
rect 4390 15473 4402 15507
rect 4436 15473 4448 15507
rect 4390 15439 4448 15473
rect 4390 15405 4402 15439
rect 4436 15405 4448 15439
rect 4390 15390 4448 15405
rect 4548 15575 4606 15590
rect 4548 15541 4560 15575
rect 4594 15541 4606 15575
rect 4548 15507 4606 15541
rect 4548 15473 4560 15507
rect 4594 15473 4606 15507
rect 4548 15439 4606 15473
rect 4548 15405 4560 15439
rect 4594 15405 4606 15439
rect 4548 15390 4606 15405
rect 4698 15575 4756 15590
rect 4698 15541 4710 15575
rect 4744 15541 4756 15575
rect 4698 15507 4756 15541
rect 4698 15473 4710 15507
rect 4744 15473 4756 15507
rect 4698 15439 4756 15473
rect 4698 15405 4710 15439
rect 4744 15405 4756 15439
rect 4698 15390 4756 15405
rect 4856 15575 4914 15590
rect 4856 15541 4868 15575
rect 4902 15541 4914 15575
rect 4856 15507 4914 15541
rect 4856 15473 4868 15507
rect 4902 15473 4914 15507
rect 4856 15439 4914 15473
rect 4856 15405 4868 15439
rect 4902 15405 4914 15439
rect 4856 15390 4914 15405
rect 5688 15576 5746 15590
rect 5688 15542 5700 15576
rect 5734 15542 5746 15576
rect 5688 15508 5746 15542
rect 5688 15474 5700 15508
rect 5734 15474 5746 15508
rect 5688 15440 5746 15474
rect 5688 15406 5700 15440
rect 5734 15406 5746 15440
rect 5688 15390 5746 15406
rect 5846 15576 5904 15590
rect 5846 15542 5858 15576
rect 5892 15542 5904 15576
rect 5846 15508 5904 15542
rect 5846 15474 5858 15508
rect 5892 15474 5904 15508
rect 5846 15440 5904 15474
rect 5846 15406 5858 15440
rect 5892 15406 5904 15440
rect 5846 15390 5904 15406
rect 5996 15576 6054 15590
rect 5996 15542 6008 15576
rect 6042 15542 6054 15576
rect 5996 15508 6054 15542
rect 5996 15474 6008 15508
rect 6042 15474 6054 15508
rect 5996 15440 6054 15474
rect 5996 15406 6008 15440
rect 6042 15406 6054 15440
rect 5996 15390 6054 15406
rect 6154 15576 6212 15590
rect 6154 15542 6166 15576
rect 6200 15542 6212 15576
rect 6154 15508 6212 15542
rect 6154 15474 6166 15508
rect 6200 15474 6212 15508
rect 6154 15440 6212 15474
rect 6154 15406 6166 15440
rect 6200 15406 6212 15440
rect 6154 15390 6212 15406
rect 6348 15576 6406 15590
rect 6348 15542 6360 15576
rect 6394 15542 6406 15576
rect 6348 15508 6406 15542
rect 6348 15474 6360 15508
rect 6394 15474 6406 15508
rect 6348 15440 6406 15474
rect 6348 15406 6360 15440
rect 6394 15406 6406 15440
rect 6348 15390 6406 15406
rect 6506 15576 6564 15590
rect 6506 15542 6518 15576
rect 6552 15542 6564 15576
rect 6506 15508 6564 15542
rect 6506 15474 6518 15508
rect 6552 15474 6564 15508
rect 6506 15440 6564 15474
rect 6506 15406 6518 15440
rect 6552 15406 6564 15440
rect 6506 15390 6564 15406
rect 6656 15576 6714 15590
rect 6656 15542 6668 15576
rect 6702 15542 6714 15576
rect 6656 15508 6714 15542
rect 6656 15474 6668 15508
rect 6702 15474 6714 15508
rect 6656 15440 6714 15474
rect 6656 15406 6668 15440
rect 6702 15406 6714 15440
rect 6656 15390 6714 15406
rect 6814 15576 6872 15590
rect 6814 15542 6826 15576
rect 6860 15542 6872 15576
rect 6814 15508 6872 15542
rect 6814 15474 6826 15508
rect 6860 15474 6872 15508
rect 6814 15440 6872 15474
rect 6814 15406 6826 15440
rect 6860 15406 6872 15440
rect 6814 15390 6872 15406
rect 1398 14337 1456 14352
rect 1398 14303 1410 14337
rect 1444 14303 1456 14337
rect 1398 14269 1456 14303
rect 1398 14235 1410 14269
rect 1444 14235 1456 14269
rect 1398 14201 1456 14235
rect 1398 14167 1410 14201
rect 1444 14167 1456 14201
rect 1398 14152 1456 14167
rect 1556 14337 1614 14352
rect 1556 14303 1568 14337
rect 1602 14303 1614 14337
rect 1556 14269 1614 14303
rect 1556 14235 1568 14269
rect 1602 14235 1614 14269
rect 1556 14201 1614 14235
rect 1556 14167 1568 14201
rect 1602 14167 1614 14201
rect 1556 14152 1614 14167
rect 1686 14337 1744 14352
rect 1686 14303 1698 14337
rect 1732 14303 1744 14337
rect 1686 14269 1744 14303
rect 1686 14235 1698 14269
rect 1732 14235 1744 14269
rect 1686 14201 1744 14235
rect 1686 14167 1698 14201
rect 1732 14167 1744 14201
rect 1686 14152 1744 14167
rect 1844 14337 1902 14352
rect 1844 14303 1856 14337
rect 1890 14303 1902 14337
rect 1844 14269 1902 14303
rect 1844 14235 1856 14269
rect 1890 14235 1902 14269
rect 1844 14201 1902 14235
rect 1844 14167 1856 14201
rect 1890 14167 1902 14201
rect 1844 14152 1902 14167
rect 2018 14337 2076 14352
rect 2018 14303 2030 14337
rect 2064 14303 2076 14337
rect 2018 14269 2076 14303
rect 2018 14235 2030 14269
rect 2064 14235 2076 14269
rect 2018 14201 2076 14235
rect 2018 14167 2030 14201
rect 2064 14167 2076 14201
rect 2018 14152 2076 14167
rect 2176 14337 2234 14352
rect 2176 14303 2188 14337
rect 2222 14303 2234 14337
rect 2176 14269 2234 14303
rect 2176 14235 2188 14269
rect 2222 14235 2234 14269
rect 2176 14201 2234 14235
rect 2176 14167 2188 14201
rect 2222 14167 2234 14201
rect 2176 14152 2234 14167
rect 2360 14337 2418 14352
rect 2360 14303 2372 14337
rect 2406 14303 2418 14337
rect 2360 14269 2418 14303
rect 2360 14235 2372 14269
rect 2406 14235 2418 14269
rect 2360 14201 2418 14235
rect 2360 14167 2372 14201
rect 2406 14167 2418 14201
rect 2360 14152 2418 14167
rect 2518 14337 2576 14352
rect 2518 14303 2530 14337
rect 2564 14303 2576 14337
rect 2518 14269 2576 14303
rect 2518 14235 2530 14269
rect 2564 14235 2576 14269
rect 2518 14201 2576 14235
rect 2518 14167 2530 14201
rect 2564 14167 2576 14201
rect 2518 14152 2576 14167
rect 2764 14337 2822 14352
rect 2764 14303 2776 14337
rect 2810 14303 2822 14337
rect 2764 14269 2822 14303
rect 2764 14235 2776 14269
rect 2810 14235 2822 14269
rect 2764 14201 2822 14235
rect 2764 14167 2776 14201
rect 2810 14167 2822 14201
rect 2764 14152 2822 14167
rect 2922 14337 2980 14352
rect 2922 14303 2934 14337
rect 2968 14303 2980 14337
rect 2922 14269 2980 14303
rect 2922 14235 2934 14269
rect 2968 14235 2980 14269
rect 2922 14201 2980 14235
rect 2922 14167 2934 14201
rect 2968 14167 2980 14201
rect 2922 14152 2980 14167
rect 3108 14337 3166 14352
rect 3108 14303 3120 14337
rect 3154 14303 3166 14337
rect 3108 14269 3166 14303
rect 3108 14235 3120 14269
rect 3154 14235 3166 14269
rect 3108 14201 3166 14235
rect 3108 14167 3120 14201
rect 3154 14167 3166 14201
rect 3108 14152 3166 14167
rect 3266 14337 3324 14352
rect 3266 14303 3278 14337
rect 3312 14303 3324 14337
rect 3266 14269 3324 14303
rect 3266 14235 3278 14269
rect 3312 14235 3324 14269
rect 3266 14201 3324 14235
rect 3266 14167 3278 14201
rect 3312 14167 3324 14201
rect 3266 14152 3324 14167
rect 3730 14347 3788 14362
rect 3730 14313 3742 14347
rect 3776 14313 3788 14347
rect 3730 14279 3788 14313
rect 3730 14245 3742 14279
rect 3776 14245 3788 14279
rect 3730 14211 3788 14245
rect 3730 14177 3742 14211
rect 3776 14177 3788 14211
rect 3730 14162 3788 14177
rect 3888 14347 3946 14362
rect 3888 14313 3900 14347
rect 3934 14313 3946 14347
rect 3888 14279 3946 14313
rect 3888 14245 3900 14279
rect 3934 14245 3946 14279
rect 3888 14211 3946 14245
rect 3888 14177 3900 14211
rect 3934 14177 3946 14211
rect 3888 14162 3946 14177
rect 4038 14347 4096 14362
rect 4038 14313 4050 14347
rect 4084 14313 4096 14347
rect 4038 14279 4096 14313
rect 4038 14245 4050 14279
rect 4084 14245 4096 14279
rect 4038 14211 4096 14245
rect 4038 14177 4050 14211
rect 4084 14177 4096 14211
rect 4038 14162 4096 14177
rect 4196 14347 4254 14362
rect 4196 14313 4208 14347
rect 4242 14313 4254 14347
rect 4196 14279 4254 14313
rect 4196 14245 4208 14279
rect 4242 14245 4254 14279
rect 4196 14211 4254 14245
rect 4196 14177 4208 14211
rect 4242 14177 4254 14211
rect 4196 14162 4254 14177
rect 4390 14347 4448 14362
rect 4390 14313 4402 14347
rect 4436 14313 4448 14347
rect 4390 14279 4448 14313
rect 4390 14245 4402 14279
rect 4436 14245 4448 14279
rect 4390 14211 4448 14245
rect 4390 14177 4402 14211
rect 4436 14177 4448 14211
rect 4390 14162 4448 14177
rect 4548 14347 4606 14362
rect 4548 14313 4560 14347
rect 4594 14313 4606 14347
rect 4548 14279 4606 14313
rect 4548 14245 4560 14279
rect 4594 14245 4606 14279
rect 4548 14211 4606 14245
rect 4548 14177 4560 14211
rect 4594 14177 4606 14211
rect 4548 14162 4606 14177
rect 4698 14347 4756 14362
rect 4698 14313 4710 14347
rect 4744 14313 4756 14347
rect 4698 14279 4756 14313
rect 4698 14245 4710 14279
rect 4744 14245 4756 14279
rect 4698 14211 4756 14245
rect 4698 14177 4710 14211
rect 4744 14177 4756 14211
rect 4698 14162 4756 14177
rect 4856 14347 4914 14362
rect 4856 14313 4868 14347
rect 4902 14313 4914 14347
rect 4856 14279 4914 14313
rect 4856 14245 4868 14279
rect 4902 14245 4914 14279
rect 4856 14211 4914 14245
rect 4856 14177 4868 14211
rect 4902 14177 4914 14211
rect 4856 14162 4914 14177
rect 5688 14348 5746 14362
rect 5688 14314 5700 14348
rect 5734 14314 5746 14348
rect 5688 14280 5746 14314
rect 5688 14246 5700 14280
rect 5734 14246 5746 14280
rect 5688 14212 5746 14246
rect 5688 14178 5700 14212
rect 5734 14178 5746 14212
rect 5688 14162 5746 14178
rect 5846 14348 5904 14362
rect 5846 14314 5858 14348
rect 5892 14314 5904 14348
rect 5846 14280 5904 14314
rect 5846 14246 5858 14280
rect 5892 14246 5904 14280
rect 5846 14212 5904 14246
rect 5846 14178 5858 14212
rect 5892 14178 5904 14212
rect 5846 14162 5904 14178
rect 5996 14348 6054 14362
rect 5996 14314 6008 14348
rect 6042 14314 6054 14348
rect 5996 14280 6054 14314
rect 5996 14246 6008 14280
rect 6042 14246 6054 14280
rect 5996 14212 6054 14246
rect 5996 14178 6008 14212
rect 6042 14178 6054 14212
rect 5996 14162 6054 14178
rect 6154 14348 6212 14362
rect 6154 14314 6166 14348
rect 6200 14314 6212 14348
rect 6154 14280 6212 14314
rect 6154 14246 6166 14280
rect 6200 14246 6212 14280
rect 6154 14212 6212 14246
rect 6154 14178 6166 14212
rect 6200 14178 6212 14212
rect 6154 14162 6212 14178
rect 6348 14348 6406 14362
rect 6348 14314 6360 14348
rect 6394 14314 6406 14348
rect 6348 14280 6406 14314
rect 6348 14246 6360 14280
rect 6394 14246 6406 14280
rect 6348 14212 6406 14246
rect 6348 14178 6360 14212
rect 6394 14178 6406 14212
rect 6348 14162 6406 14178
rect 6506 14348 6564 14362
rect 6506 14314 6518 14348
rect 6552 14314 6564 14348
rect 6506 14280 6564 14314
rect 6506 14246 6518 14280
rect 6552 14246 6564 14280
rect 6506 14212 6564 14246
rect 6506 14178 6518 14212
rect 6552 14178 6564 14212
rect 6506 14162 6564 14178
rect 6656 14348 6714 14362
rect 6656 14314 6668 14348
rect 6702 14314 6714 14348
rect 6656 14280 6714 14314
rect 6656 14246 6668 14280
rect 6702 14246 6714 14280
rect 6656 14212 6714 14246
rect 6656 14178 6668 14212
rect 6702 14178 6714 14212
rect 6656 14162 6714 14178
rect 6814 14348 6872 14362
rect 6814 14314 6826 14348
rect 6860 14314 6872 14348
rect 6814 14280 6872 14314
rect 6814 14246 6826 14280
rect 6860 14246 6872 14280
rect 6814 14212 6872 14246
rect 6814 14178 6826 14212
rect 6860 14178 6872 14212
rect 6814 14162 6872 14178
rect 1398 13109 1456 13124
rect 1398 13075 1410 13109
rect 1444 13075 1456 13109
rect 1398 13041 1456 13075
rect 1398 13007 1410 13041
rect 1444 13007 1456 13041
rect 1398 12973 1456 13007
rect 1398 12939 1410 12973
rect 1444 12939 1456 12973
rect 1398 12924 1456 12939
rect 1556 13109 1614 13124
rect 1556 13075 1568 13109
rect 1602 13075 1614 13109
rect 1556 13041 1614 13075
rect 1556 13007 1568 13041
rect 1602 13007 1614 13041
rect 1556 12973 1614 13007
rect 1556 12939 1568 12973
rect 1602 12939 1614 12973
rect 1556 12924 1614 12939
rect 1686 13109 1744 13124
rect 1686 13075 1698 13109
rect 1732 13075 1744 13109
rect 1686 13041 1744 13075
rect 1686 13007 1698 13041
rect 1732 13007 1744 13041
rect 1686 12973 1744 13007
rect 1686 12939 1698 12973
rect 1732 12939 1744 12973
rect 1686 12924 1744 12939
rect 1844 13109 1902 13124
rect 1844 13075 1856 13109
rect 1890 13075 1902 13109
rect 1844 13041 1902 13075
rect 1844 13007 1856 13041
rect 1890 13007 1902 13041
rect 1844 12973 1902 13007
rect 1844 12939 1856 12973
rect 1890 12939 1902 12973
rect 1844 12924 1902 12939
rect 2018 13109 2076 13124
rect 2018 13075 2030 13109
rect 2064 13075 2076 13109
rect 2018 13041 2076 13075
rect 2018 13007 2030 13041
rect 2064 13007 2076 13041
rect 2018 12973 2076 13007
rect 2018 12939 2030 12973
rect 2064 12939 2076 12973
rect 2018 12924 2076 12939
rect 2176 13109 2234 13124
rect 2176 13075 2188 13109
rect 2222 13075 2234 13109
rect 2176 13041 2234 13075
rect 2176 13007 2188 13041
rect 2222 13007 2234 13041
rect 2176 12973 2234 13007
rect 2176 12939 2188 12973
rect 2222 12939 2234 12973
rect 2176 12924 2234 12939
rect 2360 13109 2418 13124
rect 2360 13075 2372 13109
rect 2406 13075 2418 13109
rect 2360 13041 2418 13075
rect 2360 13007 2372 13041
rect 2406 13007 2418 13041
rect 2360 12973 2418 13007
rect 2360 12939 2372 12973
rect 2406 12939 2418 12973
rect 2360 12924 2418 12939
rect 2518 13109 2576 13124
rect 2518 13075 2530 13109
rect 2564 13075 2576 13109
rect 2518 13041 2576 13075
rect 2518 13007 2530 13041
rect 2564 13007 2576 13041
rect 2518 12973 2576 13007
rect 2518 12939 2530 12973
rect 2564 12939 2576 12973
rect 2518 12924 2576 12939
rect 2764 13109 2822 13124
rect 2764 13075 2776 13109
rect 2810 13075 2822 13109
rect 2764 13041 2822 13075
rect 2764 13007 2776 13041
rect 2810 13007 2822 13041
rect 2764 12973 2822 13007
rect 2764 12939 2776 12973
rect 2810 12939 2822 12973
rect 2764 12924 2822 12939
rect 2922 13109 2980 13124
rect 2922 13075 2934 13109
rect 2968 13075 2980 13109
rect 2922 13041 2980 13075
rect 2922 13007 2934 13041
rect 2968 13007 2980 13041
rect 2922 12973 2980 13007
rect 2922 12939 2934 12973
rect 2968 12939 2980 12973
rect 2922 12924 2980 12939
rect 3108 13109 3166 13124
rect 3108 13075 3120 13109
rect 3154 13075 3166 13109
rect 3108 13041 3166 13075
rect 3108 13007 3120 13041
rect 3154 13007 3166 13041
rect 3108 12973 3166 13007
rect 3108 12939 3120 12973
rect 3154 12939 3166 12973
rect 3108 12924 3166 12939
rect 3266 13109 3324 13124
rect 3266 13075 3278 13109
rect 3312 13075 3324 13109
rect 3266 13041 3324 13075
rect 3266 13007 3278 13041
rect 3312 13007 3324 13041
rect 3266 12973 3324 13007
rect 3266 12939 3278 12973
rect 3312 12939 3324 12973
rect 3266 12924 3324 12939
rect 3730 13119 3788 13134
rect 3730 13085 3742 13119
rect 3776 13085 3788 13119
rect 3730 13051 3788 13085
rect 3730 13017 3742 13051
rect 3776 13017 3788 13051
rect 3730 12983 3788 13017
rect 3730 12949 3742 12983
rect 3776 12949 3788 12983
rect 3730 12934 3788 12949
rect 3888 13119 3946 13134
rect 3888 13085 3900 13119
rect 3934 13085 3946 13119
rect 3888 13051 3946 13085
rect 3888 13017 3900 13051
rect 3934 13017 3946 13051
rect 3888 12983 3946 13017
rect 3888 12949 3900 12983
rect 3934 12949 3946 12983
rect 3888 12934 3946 12949
rect 4038 13119 4096 13134
rect 4038 13085 4050 13119
rect 4084 13085 4096 13119
rect 4038 13051 4096 13085
rect 4038 13017 4050 13051
rect 4084 13017 4096 13051
rect 4038 12983 4096 13017
rect 4038 12949 4050 12983
rect 4084 12949 4096 12983
rect 4038 12934 4096 12949
rect 4196 13119 4254 13134
rect 4196 13085 4208 13119
rect 4242 13085 4254 13119
rect 4196 13051 4254 13085
rect 4196 13017 4208 13051
rect 4242 13017 4254 13051
rect 4196 12983 4254 13017
rect 4196 12949 4208 12983
rect 4242 12949 4254 12983
rect 4196 12934 4254 12949
rect 4390 13119 4448 13134
rect 4390 13085 4402 13119
rect 4436 13085 4448 13119
rect 4390 13051 4448 13085
rect 4390 13017 4402 13051
rect 4436 13017 4448 13051
rect 4390 12983 4448 13017
rect 4390 12949 4402 12983
rect 4436 12949 4448 12983
rect 4390 12934 4448 12949
rect 4548 13119 4606 13134
rect 4548 13085 4560 13119
rect 4594 13085 4606 13119
rect 4548 13051 4606 13085
rect 4548 13017 4560 13051
rect 4594 13017 4606 13051
rect 4548 12983 4606 13017
rect 4548 12949 4560 12983
rect 4594 12949 4606 12983
rect 4548 12934 4606 12949
rect 4698 13119 4756 13134
rect 4698 13085 4710 13119
rect 4744 13085 4756 13119
rect 4698 13051 4756 13085
rect 4698 13017 4710 13051
rect 4744 13017 4756 13051
rect 4698 12983 4756 13017
rect 4698 12949 4710 12983
rect 4744 12949 4756 12983
rect 4698 12934 4756 12949
rect 4856 13119 4914 13134
rect 4856 13085 4868 13119
rect 4902 13085 4914 13119
rect 4856 13051 4914 13085
rect 4856 13017 4868 13051
rect 4902 13017 4914 13051
rect 4856 12983 4914 13017
rect 4856 12949 4868 12983
rect 4902 12949 4914 12983
rect 4856 12934 4914 12949
rect 5688 13120 5746 13134
rect 5688 13086 5700 13120
rect 5734 13086 5746 13120
rect 5688 13052 5746 13086
rect 5688 13018 5700 13052
rect 5734 13018 5746 13052
rect 5688 12984 5746 13018
rect 5688 12950 5700 12984
rect 5734 12950 5746 12984
rect 5688 12934 5746 12950
rect 5846 13120 5904 13134
rect 5846 13086 5858 13120
rect 5892 13086 5904 13120
rect 5846 13052 5904 13086
rect 5846 13018 5858 13052
rect 5892 13018 5904 13052
rect 5846 12984 5904 13018
rect 5846 12950 5858 12984
rect 5892 12950 5904 12984
rect 5846 12934 5904 12950
rect 5996 13120 6054 13134
rect 5996 13086 6008 13120
rect 6042 13086 6054 13120
rect 5996 13052 6054 13086
rect 5996 13018 6008 13052
rect 6042 13018 6054 13052
rect 5996 12984 6054 13018
rect 5996 12950 6008 12984
rect 6042 12950 6054 12984
rect 5996 12934 6054 12950
rect 6154 13120 6212 13134
rect 6154 13086 6166 13120
rect 6200 13086 6212 13120
rect 6154 13052 6212 13086
rect 6154 13018 6166 13052
rect 6200 13018 6212 13052
rect 6154 12984 6212 13018
rect 6154 12950 6166 12984
rect 6200 12950 6212 12984
rect 6154 12934 6212 12950
rect 6348 13120 6406 13134
rect 6348 13086 6360 13120
rect 6394 13086 6406 13120
rect 6348 13052 6406 13086
rect 6348 13018 6360 13052
rect 6394 13018 6406 13052
rect 6348 12984 6406 13018
rect 6348 12950 6360 12984
rect 6394 12950 6406 12984
rect 6348 12934 6406 12950
rect 6506 13120 6564 13134
rect 6506 13086 6518 13120
rect 6552 13086 6564 13120
rect 6506 13052 6564 13086
rect 6506 13018 6518 13052
rect 6552 13018 6564 13052
rect 6506 12984 6564 13018
rect 6506 12950 6518 12984
rect 6552 12950 6564 12984
rect 6506 12934 6564 12950
rect 6656 13120 6714 13134
rect 6656 13086 6668 13120
rect 6702 13086 6714 13120
rect 6656 13052 6714 13086
rect 6656 13018 6668 13052
rect 6702 13018 6714 13052
rect 6656 12984 6714 13018
rect 6656 12950 6668 12984
rect 6702 12950 6714 12984
rect 6656 12934 6714 12950
rect 6814 13120 6872 13134
rect 6814 13086 6826 13120
rect 6860 13086 6872 13120
rect 6814 13052 6872 13086
rect 6814 13018 6826 13052
rect 6860 13018 6872 13052
rect 6814 12984 6872 13018
rect 6814 12950 6826 12984
rect 6860 12950 6872 12984
rect 6814 12934 6872 12950
rect 1398 11881 1456 11896
rect 1398 11847 1410 11881
rect 1444 11847 1456 11881
rect 1398 11813 1456 11847
rect 1398 11779 1410 11813
rect 1444 11779 1456 11813
rect 1398 11745 1456 11779
rect 1398 11711 1410 11745
rect 1444 11711 1456 11745
rect 1398 11696 1456 11711
rect 1556 11881 1614 11896
rect 1556 11847 1568 11881
rect 1602 11847 1614 11881
rect 1556 11813 1614 11847
rect 1556 11779 1568 11813
rect 1602 11779 1614 11813
rect 1556 11745 1614 11779
rect 1556 11711 1568 11745
rect 1602 11711 1614 11745
rect 1556 11696 1614 11711
rect 1686 11881 1744 11896
rect 1686 11847 1698 11881
rect 1732 11847 1744 11881
rect 1686 11813 1744 11847
rect 1686 11779 1698 11813
rect 1732 11779 1744 11813
rect 1686 11745 1744 11779
rect 1686 11711 1698 11745
rect 1732 11711 1744 11745
rect 1686 11696 1744 11711
rect 1844 11881 1902 11896
rect 1844 11847 1856 11881
rect 1890 11847 1902 11881
rect 1844 11813 1902 11847
rect 1844 11779 1856 11813
rect 1890 11779 1902 11813
rect 1844 11745 1902 11779
rect 1844 11711 1856 11745
rect 1890 11711 1902 11745
rect 1844 11696 1902 11711
rect 2018 11881 2076 11896
rect 2018 11847 2030 11881
rect 2064 11847 2076 11881
rect 2018 11813 2076 11847
rect 2018 11779 2030 11813
rect 2064 11779 2076 11813
rect 2018 11745 2076 11779
rect 2018 11711 2030 11745
rect 2064 11711 2076 11745
rect 2018 11696 2076 11711
rect 2176 11881 2234 11896
rect 2176 11847 2188 11881
rect 2222 11847 2234 11881
rect 2176 11813 2234 11847
rect 2176 11779 2188 11813
rect 2222 11779 2234 11813
rect 2176 11745 2234 11779
rect 2176 11711 2188 11745
rect 2222 11711 2234 11745
rect 2176 11696 2234 11711
rect 2360 11881 2418 11896
rect 2360 11847 2372 11881
rect 2406 11847 2418 11881
rect 2360 11813 2418 11847
rect 2360 11779 2372 11813
rect 2406 11779 2418 11813
rect 2360 11745 2418 11779
rect 2360 11711 2372 11745
rect 2406 11711 2418 11745
rect 2360 11696 2418 11711
rect 2518 11881 2576 11896
rect 2518 11847 2530 11881
rect 2564 11847 2576 11881
rect 2518 11813 2576 11847
rect 2518 11779 2530 11813
rect 2564 11779 2576 11813
rect 2518 11745 2576 11779
rect 2518 11711 2530 11745
rect 2564 11711 2576 11745
rect 2518 11696 2576 11711
rect 2764 11881 2822 11896
rect 2764 11847 2776 11881
rect 2810 11847 2822 11881
rect 2764 11813 2822 11847
rect 2764 11779 2776 11813
rect 2810 11779 2822 11813
rect 2764 11745 2822 11779
rect 2764 11711 2776 11745
rect 2810 11711 2822 11745
rect 2764 11696 2822 11711
rect 2922 11881 2980 11896
rect 2922 11847 2934 11881
rect 2968 11847 2980 11881
rect 2922 11813 2980 11847
rect 2922 11779 2934 11813
rect 2968 11779 2980 11813
rect 2922 11745 2980 11779
rect 2922 11711 2934 11745
rect 2968 11711 2980 11745
rect 2922 11696 2980 11711
rect 3108 11881 3166 11896
rect 3108 11847 3120 11881
rect 3154 11847 3166 11881
rect 3108 11813 3166 11847
rect 3108 11779 3120 11813
rect 3154 11779 3166 11813
rect 3108 11745 3166 11779
rect 3108 11711 3120 11745
rect 3154 11711 3166 11745
rect 3108 11696 3166 11711
rect 3266 11881 3324 11896
rect 3266 11847 3278 11881
rect 3312 11847 3324 11881
rect 3266 11813 3324 11847
rect 3266 11779 3278 11813
rect 3312 11779 3324 11813
rect 3266 11745 3324 11779
rect 3266 11711 3278 11745
rect 3312 11711 3324 11745
rect 3266 11696 3324 11711
rect 3730 11891 3788 11906
rect 3730 11857 3742 11891
rect 3776 11857 3788 11891
rect 3730 11823 3788 11857
rect 3730 11789 3742 11823
rect 3776 11789 3788 11823
rect 3730 11755 3788 11789
rect 3730 11721 3742 11755
rect 3776 11721 3788 11755
rect 3730 11706 3788 11721
rect 3888 11891 3946 11906
rect 3888 11857 3900 11891
rect 3934 11857 3946 11891
rect 3888 11823 3946 11857
rect 3888 11789 3900 11823
rect 3934 11789 3946 11823
rect 3888 11755 3946 11789
rect 3888 11721 3900 11755
rect 3934 11721 3946 11755
rect 3888 11706 3946 11721
rect 4038 11891 4096 11906
rect 4038 11857 4050 11891
rect 4084 11857 4096 11891
rect 4038 11823 4096 11857
rect 4038 11789 4050 11823
rect 4084 11789 4096 11823
rect 4038 11755 4096 11789
rect 4038 11721 4050 11755
rect 4084 11721 4096 11755
rect 4038 11706 4096 11721
rect 4196 11891 4254 11906
rect 4196 11857 4208 11891
rect 4242 11857 4254 11891
rect 4196 11823 4254 11857
rect 4196 11789 4208 11823
rect 4242 11789 4254 11823
rect 4196 11755 4254 11789
rect 4196 11721 4208 11755
rect 4242 11721 4254 11755
rect 4196 11706 4254 11721
rect 4390 11891 4448 11906
rect 4390 11857 4402 11891
rect 4436 11857 4448 11891
rect 4390 11823 4448 11857
rect 4390 11789 4402 11823
rect 4436 11789 4448 11823
rect 4390 11755 4448 11789
rect 4390 11721 4402 11755
rect 4436 11721 4448 11755
rect 4390 11706 4448 11721
rect 4548 11891 4606 11906
rect 4548 11857 4560 11891
rect 4594 11857 4606 11891
rect 4548 11823 4606 11857
rect 4548 11789 4560 11823
rect 4594 11789 4606 11823
rect 4548 11755 4606 11789
rect 4548 11721 4560 11755
rect 4594 11721 4606 11755
rect 4548 11706 4606 11721
rect 4698 11891 4756 11906
rect 4698 11857 4710 11891
rect 4744 11857 4756 11891
rect 4698 11823 4756 11857
rect 4698 11789 4710 11823
rect 4744 11789 4756 11823
rect 4698 11755 4756 11789
rect 4698 11721 4710 11755
rect 4744 11721 4756 11755
rect 4698 11706 4756 11721
rect 4856 11891 4914 11906
rect 4856 11857 4868 11891
rect 4902 11857 4914 11891
rect 4856 11823 4914 11857
rect 4856 11789 4868 11823
rect 4902 11789 4914 11823
rect 4856 11755 4914 11789
rect 4856 11721 4868 11755
rect 4902 11721 4914 11755
rect 4856 11706 4914 11721
rect 5688 11892 5746 11906
rect 5688 11858 5700 11892
rect 5734 11858 5746 11892
rect 5688 11824 5746 11858
rect 5688 11790 5700 11824
rect 5734 11790 5746 11824
rect 5688 11756 5746 11790
rect 5688 11722 5700 11756
rect 5734 11722 5746 11756
rect 5688 11706 5746 11722
rect 5846 11892 5904 11906
rect 5846 11858 5858 11892
rect 5892 11858 5904 11892
rect 5846 11824 5904 11858
rect 5846 11790 5858 11824
rect 5892 11790 5904 11824
rect 5846 11756 5904 11790
rect 5846 11722 5858 11756
rect 5892 11722 5904 11756
rect 5846 11706 5904 11722
rect 5996 11892 6054 11906
rect 5996 11858 6008 11892
rect 6042 11858 6054 11892
rect 5996 11824 6054 11858
rect 5996 11790 6008 11824
rect 6042 11790 6054 11824
rect 5996 11756 6054 11790
rect 5996 11722 6008 11756
rect 6042 11722 6054 11756
rect 5996 11706 6054 11722
rect 6154 11892 6212 11906
rect 6154 11858 6166 11892
rect 6200 11858 6212 11892
rect 6154 11824 6212 11858
rect 6154 11790 6166 11824
rect 6200 11790 6212 11824
rect 6154 11756 6212 11790
rect 6154 11722 6166 11756
rect 6200 11722 6212 11756
rect 6154 11706 6212 11722
rect 6348 11892 6406 11906
rect 6348 11858 6360 11892
rect 6394 11858 6406 11892
rect 6348 11824 6406 11858
rect 6348 11790 6360 11824
rect 6394 11790 6406 11824
rect 6348 11756 6406 11790
rect 6348 11722 6360 11756
rect 6394 11722 6406 11756
rect 6348 11706 6406 11722
rect 6506 11892 6564 11906
rect 6506 11858 6518 11892
rect 6552 11858 6564 11892
rect 6506 11824 6564 11858
rect 6506 11790 6518 11824
rect 6552 11790 6564 11824
rect 6506 11756 6564 11790
rect 6506 11722 6518 11756
rect 6552 11722 6564 11756
rect 6506 11706 6564 11722
rect 6656 11892 6714 11906
rect 6656 11858 6668 11892
rect 6702 11858 6714 11892
rect 6656 11824 6714 11858
rect 6656 11790 6668 11824
rect 6702 11790 6714 11824
rect 6656 11756 6714 11790
rect 6656 11722 6668 11756
rect 6702 11722 6714 11756
rect 6656 11706 6714 11722
rect 6814 11892 6872 11906
rect 6814 11858 6826 11892
rect 6860 11858 6872 11892
rect 6814 11824 6872 11858
rect 6814 11790 6826 11824
rect 6860 11790 6872 11824
rect 6814 11756 6872 11790
rect 6814 11722 6826 11756
rect 6860 11722 6872 11756
rect 6814 11706 6872 11722
rect 1398 10653 1456 10668
rect 1398 10619 1410 10653
rect 1444 10619 1456 10653
rect 1398 10585 1456 10619
rect 1398 10551 1410 10585
rect 1444 10551 1456 10585
rect 1398 10517 1456 10551
rect 1398 10483 1410 10517
rect 1444 10483 1456 10517
rect 1398 10468 1456 10483
rect 1556 10653 1614 10668
rect 1556 10619 1568 10653
rect 1602 10619 1614 10653
rect 1556 10585 1614 10619
rect 1556 10551 1568 10585
rect 1602 10551 1614 10585
rect 1556 10517 1614 10551
rect 1556 10483 1568 10517
rect 1602 10483 1614 10517
rect 1556 10468 1614 10483
rect 1686 10653 1744 10668
rect 1686 10619 1698 10653
rect 1732 10619 1744 10653
rect 1686 10585 1744 10619
rect 1686 10551 1698 10585
rect 1732 10551 1744 10585
rect 1686 10517 1744 10551
rect 1686 10483 1698 10517
rect 1732 10483 1744 10517
rect 1686 10468 1744 10483
rect 1844 10653 1902 10668
rect 1844 10619 1856 10653
rect 1890 10619 1902 10653
rect 1844 10585 1902 10619
rect 1844 10551 1856 10585
rect 1890 10551 1902 10585
rect 1844 10517 1902 10551
rect 1844 10483 1856 10517
rect 1890 10483 1902 10517
rect 1844 10468 1902 10483
rect 2018 10653 2076 10668
rect 2018 10619 2030 10653
rect 2064 10619 2076 10653
rect 2018 10585 2076 10619
rect 2018 10551 2030 10585
rect 2064 10551 2076 10585
rect 2018 10517 2076 10551
rect 2018 10483 2030 10517
rect 2064 10483 2076 10517
rect 2018 10468 2076 10483
rect 2176 10653 2234 10668
rect 2176 10619 2188 10653
rect 2222 10619 2234 10653
rect 2176 10585 2234 10619
rect 2176 10551 2188 10585
rect 2222 10551 2234 10585
rect 2176 10517 2234 10551
rect 2176 10483 2188 10517
rect 2222 10483 2234 10517
rect 2176 10468 2234 10483
rect 2360 10653 2418 10668
rect 2360 10619 2372 10653
rect 2406 10619 2418 10653
rect 2360 10585 2418 10619
rect 2360 10551 2372 10585
rect 2406 10551 2418 10585
rect 2360 10517 2418 10551
rect 2360 10483 2372 10517
rect 2406 10483 2418 10517
rect 2360 10468 2418 10483
rect 2518 10653 2576 10668
rect 2518 10619 2530 10653
rect 2564 10619 2576 10653
rect 2518 10585 2576 10619
rect 2518 10551 2530 10585
rect 2564 10551 2576 10585
rect 2518 10517 2576 10551
rect 2518 10483 2530 10517
rect 2564 10483 2576 10517
rect 2518 10468 2576 10483
rect 2764 10653 2822 10668
rect 2764 10619 2776 10653
rect 2810 10619 2822 10653
rect 2764 10585 2822 10619
rect 2764 10551 2776 10585
rect 2810 10551 2822 10585
rect 2764 10517 2822 10551
rect 2764 10483 2776 10517
rect 2810 10483 2822 10517
rect 2764 10468 2822 10483
rect 2922 10653 2980 10668
rect 2922 10619 2934 10653
rect 2968 10619 2980 10653
rect 2922 10585 2980 10619
rect 2922 10551 2934 10585
rect 2968 10551 2980 10585
rect 2922 10517 2980 10551
rect 2922 10483 2934 10517
rect 2968 10483 2980 10517
rect 2922 10468 2980 10483
rect 3108 10653 3166 10668
rect 3108 10619 3120 10653
rect 3154 10619 3166 10653
rect 3108 10585 3166 10619
rect 3108 10551 3120 10585
rect 3154 10551 3166 10585
rect 3108 10517 3166 10551
rect 3108 10483 3120 10517
rect 3154 10483 3166 10517
rect 3108 10468 3166 10483
rect 3266 10653 3324 10668
rect 3266 10619 3278 10653
rect 3312 10619 3324 10653
rect 3266 10585 3324 10619
rect 3266 10551 3278 10585
rect 3312 10551 3324 10585
rect 3266 10517 3324 10551
rect 3266 10483 3278 10517
rect 3312 10483 3324 10517
rect 3266 10468 3324 10483
rect 3730 10663 3788 10678
rect 3730 10629 3742 10663
rect 3776 10629 3788 10663
rect 3730 10595 3788 10629
rect 3730 10561 3742 10595
rect 3776 10561 3788 10595
rect 3730 10527 3788 10561
rect 3730 10493 3742 10527
rect 3776 10493 3788 10527
rect 3730 10478 3788 10493
rect 3888 10663 3946 10678
rect 3888 10629 3900 10663
rect 3934 10629 3946 10663
rect 3888 10595 3946 10629
rect 3888 10561 3900 10595
rect 3934 10561 3946 10595
rect 3888 10527 3946 10561
rect 3888 10493 3900 10527
rect 3934 10493 3946 10527
rect 3888 10478 3946 10493
rect 4038 10663 4096 10678
rect 4038 10629 4050 10663
rect 4084 10629 4096 10663
rect 4038 10595 4096 10629
rect 4038 10561 4050 10595
rect 4084 10561 4096 10595
rect 4038 10527 4096 10561
rect 4038 10493 4050 10527
rect 4084 10493 4096 10527
rect 4038 10478 4096 10493
rect 4196 10663 4254 10678
rect 4196 10629 4208 10663
rect 4242 10629 4254 10663
rect 4196 10595 4254 10629
rect 4196 10561 4208 10595
rect 4242 10561 4254 10595
rect 4196 10527 4254 10561
rect 4196 10493 4208 10527
rect 4242 10493 4254 10527
rect 4196 10478 4254 10493
rect 4390 10663 4448 10678
rect 4390 10629 4402 10663
rect 4436 10629 4448 10663
rect 4390 10595 4448 10629
rect 4390 10561 4402 10595
rect 4436 10561 4448 10595
rect 4390 10527 4448 10561
rect 4390 10493 4402 10527
rect 4436 10493 4448 10527
rect 4390 10478 4448 10493
rect 4548 10663 4606 10678
rect 4548 10629 4560 10663
rect 4594 10629 4606 10663
rect 4548 10595 4606 10629
rect 4548 10561 4560 10595
rect 4594 10561 4606 10595
rect 4548 10527 4606 10561
rect 4548 10493 4560 10527
rect 4594 10493 4606 10527
rect 4548 10478 4606 10493
rect 4698 10663 4756 10678
rect 4698 10629 4710 10663
rect 4744 10629 4756 10663
rect 4698 10595 4756 10629
rect 4698 10561 4710 10595
rect 4744 10561 4756 10595
rect 4698 10527 4756 10561
rect 4698 10493 4710 10527
rect 4744 10493 4756 10527
rect 4698 10478 4756 10493
rect 4856 10663 4914 10678
rect 4856 10629 4868 10663
rect 4902 10629 4914 10663
rect 4856 10595 4914 10629
rect 4856 10561 4868 10595
rect 4902 10561 4914 10595
rect 4856 10527 4914 10561
rect 4856 10493 4868 10527
rect 4902 10493 4914 10527
rect 4856 10478 4914 10493
rect 5688 10664 5746 10678
rect 5688 10630 5700 10664
rect 5734 10630 5746 10664
rect 5688 10596 5746 10630
rect 5688 10562 5700 10596
rect 5734 10562 5746 10596
rect 5688 10528 5746 10562
rect 5688 10494 5700 10528
rect 5734 10494 5746 10528
rect 5688 10478 5746 10494
rect 5846 10664 5904 10678
rect 5846 10630 5858 10664
rect 5892 10630 5904 10664
rect 5846 10596 5904 10630
rect 5846 10562 5858 10596
rect 5892 10562 5904 10596
rect 5846 10528 5904 10562
rect 5846 10494 5858 10528
rect 5892 10494 5904 10528
rect 5846 10478 5904 10494
rect 5996 10664 6054 10678
rect 5996 10630 6008 10664
rect 6042 10630 6054 10664
rect 5996 10596 6054 10630
rect 5996 10562 6008 10596
rect 6042 10562 6054 10596
rect 5996 10528 6054 10562
rect 5996 10494 6008 10528
rect 6042 10494 6054 10528
rect 5996 10478 6054 10494
rect 6154 10664 6212 10678
rect 6154 10630 6166 10664
rect 6200 10630 6212 10664
rect 6154 10596 6212 10630
rect 6154 10562 6166 10596
rect 6200 10562 6212 10596
rect 6154 10528 6212 10562
rect 6154 10494 6166 10528
rect 6200 10494 6212 10528
rect 6154 10478 6212 10494
rect 6348 10664 6406 10678
rect 6348 10630 6360 10664
rect 6394 10630 6406 10664
rect 6348 10596 6406 10630
rect 6348 10562 6360 10596
rect 6394 10562 6406 10596
rect 6348 10528 6406 10562
rect 6348 10494 6360 10528
rect 6394 10494 6406 10528
rect 6348 10478 6406 10494
rect 6506 10664 6564 10678
rect 6506 10630 6518 10664
rect 6552 10630 6564 10664
rect 6506 10596 6564 10630
rect 6506 10562 6518 10596
rect 6552 10562 6564 10596
rect 6506 10528 6564 10562
rect 6506 10494 6518 10528
rect 6552 10494 6564 10528
rect 6506 10478 6564 10494
rect 6656 10664 6714 10678
rect 6656 10630 6668 10664
rect 6702 10630 6714 10664
rect 6656 10596 6714 10630
rect 6656 10562 6668 10596
rect 6702 10562 6714 10596
rect 6656 10528 6714 10562
rect 6656 10494 6668 10528
rect 6702 10494 6714 10528
rect 6656 10478 6714 10494
rect 6814 10664 6872 10678
rect 6814 10630 6826 10664
rect 6860 10630 6872 10664
rect 6814 10596 6872 10630
rect 6814 10562 6826 10596
rect 6860 10562 6872 10596
rect 6814 10528 6872 10562
rect 6814 10494 6826 10528
rect 6860 10494 6872 10528
rect 6814 10478 6872 10494
rect 1398 9425 1456 9440
rect 1398 9391 1410 9425
rect 1444 9391 1456 9425
rect 1398 9357 1456 9391
rect 1398 9323 1410 9357
rect 1444 9323 1456 9357
rect 1398 9289 1456 9323
rect 1398 9255 1410 9289
rect 1444 9255 1456 9289
rect 1398 9240 1456 9255
rect 1556 9425 1614 9440
rect 1556 9391 1568 9425
rect 1602 9391 1614 9425
rect 1556 9357 1614 9391
rect 1556 9323 1568 9357
rect 1602 9323 1614 9357
rect 1556 9289 1614 9323
rect 1556 9255 1568 9289
rect 1602 9255 1614 9289
rect 1556 9240 1614 9255
rect 1686 9425 1744 9440
rect 1686 9391 1698 9425
rect 1732 9391 1744 9425
rect 1686 9357 1744 9391
rect 1686 9323 1698 9357
rect 1732 9323 1744 9357
rect 1686 9289 1744 9323
rect 1686 9255 1698 9289
rect 1732 9255 1744 9289
rect 1686 9240 1744 9255
rect 1844 9425 1902 9440
rect 1844 9391 1856 9425
rect 1890 9391 1902 9425
rect 1844 9357 1902 9391
rect 1844 9323 1856 9357
rect 1890 9323 1902 9357
rect 1844 9289 1902 9323
rect 1844 9255 1856 9289
rect 1890 9255 1902 9289
rect 1844 9240 1902 9255
rect 2018 9425 2076 9440
rect 2018 9391 2030 9425
rect 2064 9391 2076 9425
rect 2018 9357 2076 9391
rect 2018 9323 2030 9357
rect 2064 9323 2076 9357
rect 2018 9289 2076 9323
rect 2018 9255 2030 9289
rect 2064 9255 2076 9289
rect 2018 9240 2076 9255
rect 2176 9425 2234 9440
rect 2176 9391 2188 9425
rect 2222 9391 2234 9425
rect 2176 9357 2234 9391
rect 2176 9323 2188 9357
rect 2222 9323 2234 9357
rect 2176 9289 2234 9323
rect 2176 9255 2188 9289
rect 2222 9255 2234 9289
rect 2176 9240 2234 9255
rect 2360 9425 2418 9440
rect 2360 9391 2372 9425
rect 2406 9391 2418 9425
rect 2360 9357 2418 9391
rect 2360 9323 2372 9357
rect 2406 9323 2418 9357
rect 2360 9289 2418 9323
rect 2360 9255 2372 9289
rect 2406 9255 2418 9289
rect 2360 9240 2418 9255
rect 2518 9425 2576 9440
rect 2518 9391 2530 9425
rect 2564 9391 2576 9425
rect 2518 9357 2576 9391
rect 2518 9323 2530 9357
rect 2564 9323 2576 9357
rect 2518 9289 2576 9323
rect 2518 9255 2530 9289
rect 2564 9255 2576 9289
rect 2518 9240 2576 9255
rect 2764 9425 2822 9440
rect 2764 9391 2776 9425
rect 2810 9391 2822 9425
rect 2764 9357 2822 9391
rect 2764 9323 2776 9357
rect 2810 9323 2822 9357
rect 2764 9289 2822 9323
rect 2764 9255 2776 9289
rect 2810 9255 2822 9289
rect 2764 9240 2822 9255
rect 2922 9425 2980 9440
rect 2922 9391 2934 9425
rect 2968 9391 2980 9425
rect 2922 9357 2980 9391
rect 2922 9323 2934 9357
rect 2968 9323 2980 9357
rect 2922 9289 2980 9323
rect 2922 9255 2934 9289
rect 2968 9255 2980 9289
rect 2922 9240 2980 9255
rect 3108 9425 3166 9440
rect 3108 9391 3120 9425
rect 3154 9391 3166 9425
rect 3108 9357 3166 9391
rect 3108 9323 3120 9357
rect 3154 9323 3166 9357
rect 3108 9289 3166 9323
rect 3108 9255 3120 9289
rect 3154 9255 3166 9289
rect 3108 9240 3166 9255
rect 3266 9425 3324 9440
rect 3266 9391 3278 9425
rect 3312 9391 3324 9425
rect 3266 9357 3324 9391
rect 3266 9323 3278 9357
rect 3312 9323 3324 9357
rect 3266 9289 3324 9323
rect 3266 9255 3278 9289
rect 3312 9255 3324 9289
rect 3266 9240 3324 9255
rect 3730 9435 3788 9450
rect 3730 9401 3742 9435
rect 3776 9401 3788 9435
rect 3730 9367 3788 9401
rect 3730 9333 3742 9367
rect 3776 9333 3788 9367
rect 3730 9299 3788 9333
rect 3730 9265 3742 9299
rect 3776 9265 3788 9299
rect 3730 9250 3788 9265
rect 3888 9435 3946 9450
rect 3888 9401 3900 9435
rect 3934 9401 3946 9435
rect 3888 9367 3946 9401
rect 3888 9333 3900 9367
rect 3934 9333 3946 9367
rect 3888 9299 3946 9333
rect 3888 9265 3900 9299
rect 3934 9265 3946 9299
rect 3888 9250 3946 9265
rect 4038 9435 4096 9450
rect 4038 9401 4050 9435
rect 4084 9401 4096 9435
rect 4038 9367 4096 9401
rect 4038 9333 4050 9367
rect 4084 9333 4096 9367
rect 4038 9299 4096 9333
rect 4038 9265 4050 9299
rect 4084 9265 4096 9299
rect 4038 9250 4096 9265
rect 4196 9435 4254 9450
rect 4196 9401 4208 9435
rect 4242 9401 4254 9435
rect 4196 9367 4254 9401
rect 4196 9333 4208 9367
rect 4242 9333 4254 9367
rect 4196 9299 4254 9333
rect 4196 9265 4208 9299
rect 4242 9265 4254 9299
rect 4196 9250 4254 9265
rect 4390 9435 4448 9450
rect 4390 9401 4402 9435
rect 4436 9401 4448 9435
rect 4390 9367 4448 9401
rect 4390 9333 4402 9367
rect 4436 9333 4448 9367
rect 4390 9299 4448 9333
rect 4390 9265 4402 9299
rect 4436 9265 4448 9299
rect 4390 9250 4448 9265
rect 4548 9435 4606 9450
rect 4548 9401 4560 9435
rect 4594 9401 4606 9435
rect 4548 9367 4606 9401
rect 4548 9333 4560 9367
rect 4594 9333 4606 9367
rect 4548 9299 4606 9333
rect 4548 9265 4560 9299
rect 4594 9265 4606 9299
rect 4548 9250 4606 9265
rect 4698 9435 4756 9450
rect 4698 9401 4710 9435
rect 4744 9401 4756 9435
rect 4698 9367 4756 9401
rect 4698 9333 4710 9367
rect 4744 9333 4756 9367
rect 4698 9299 4756 9333
rect 4698 9265 4710 9299
rect 4744 9265 4756 9299
rect 4698 9250 4756 9265
rect 4856 9435 4914 9450
rect 4856 9401 4868 9435
rect 4902 9401 4914 9435
rect 4856 9367 4914 9401
rect 4856 9333 4868 9367
rect 4902 9333 4914 9367
rect 4856 9299 4914 9333
rect 4856 9265 4868 9299
rect 4902 9265 4914 9299
rect 4856 9250 4914 9265
rect 5688 9436 5746 9450
rect 5688 9402 5700 9436
rect 5734 9402 5746 9436
rect 5688 9368 5746 9402
rect 5688 9334 5700 9368
rect 5734 9334 5746 9368
rect 5688 9300 5746 9334
rect 5688 9266 5700 9300
rect 5734 9266 5746 9300
rect 5688 9250 5746 9266
rect 5846 9436 5904 9450
rect 5846 9402 5858 9436
rect 5892 9402 5904 9436
rect 5846 9368 5904 9402
rect 5846 9334 5858 9368
rect 5892 9334 5904 9368
rect 5846 9300 5904 9334
rect 5846 9266 5858 9300
rect 5892 9266 5904 9300
rect 5846 9250 5904 9266
rect 5996 9436 6054 9450
rect 5996 9402 6008 9436
rect 6042 9402 6054 9436
rect 5996 9368 6054 9402
rect 5996 9334 6008 9368
rect 6042 9334 6054 9368
rect 5996 9300 6054 9334
rect 5996 9266 6008 9300
rect 6042 9266 6054 9300
rect 5996 9250 6054 9266
rect 6154 9436 6212 9450
rect 6154 9402 6166 9436
rect 6200 9402 6212 9436
rect 6154 9368 6212 9402
rect 6154 9334 6166 9368
rect 6200 9334 6212 9368
rect 6154 9300 6212 9334
rect 6154 9266 6166 9300
rect 6200 9266 6212 9300
rect 6154 9250 6212 9266
rect 6348 9436 6406 9450
rect 6348 9402 6360 9436
rect 6394 9402 6406 9436
rect 6348 9368 6406 9402
rect 6348 9334 6360 9368
rect 6394 9334 6406 9368
rect 6348 9300 6406 9334
rect 6348 9266 6360 9300
rect 6394 9266 6406 9300
rect 6348 9250 6406 9266
rect 6506 9436 6564 9450
rect 6506 9402 6518 9436
rect 6552 9402 6564 9436
rect 6506 9368 6564 9402
rect 6506 9334 6518 9368
rect 6552 9334 6564 9368
rect 6506 9300 6564 9334
rect 6506 9266 6518 9300
rect 6552 9266 6564 9300
rect 6506 9250 6564 9266
rect 6656 9436 6714 9450
rect 6656 9402 6668 9436
rect 6702 9402 6714 9436
rect 6656 9368 6714 9402
rect 6656 9334 6668 9368
rect 6702 9334 6714 9368
rect 6656 9300 6714 9334
rect 6656 9266 6668 9300
rect 6702 9266 6714 9300
rect 6656 9250 6714 9266
rect 6814 9436 6872 9450
rect 6814 9402 6826 9436
rect 6860 9402 6872 9436
rect 6814 9368 6872 9402
rect 6814 9334 6826 9368
rect 6860 9334 6872 9368
rect 6814 9300 6872 9334
rect 6814 9266 6826 9300
rect 6860 9266 6872 9300
rect 6814 9250 6872 9266
rect 1398 8197 1456 8212
rect 1398 8163 1410 8197
rect 1444 8163 1456 8197
rect 1398 8129 1456 8163
rect 1398 8095 1410 8129
rect 1444 8095 1456 8129
rect 1398 8061 1456 8095
rect 1398 8027 1410 8061
rect 1444 8027 1456 8061
rect 1398 8012 1456 8027
rect 1556 8197 1614 8212
rect 1556 8163 1568 8197
rect 1602 8163 1614 8197
rect 1556 8129 1614 8163
rect 1556 8095 1568 8129
rect 1602 8095 1614 8129
rect 1556 8061 1614 8095
rect 1556 8027 1568 8061
rect 1602 8027 1614 8061
rect 1556 8012 1614 8027
rect 1686 8197 1744 8212
rect 1686 8163 1698 8197
rect 1732 8163 1744 8197
rect 1686 8129 1744 8163
rect 1686 8095 1698 8129
rect 1732 8095 1744 8129
rect 1686 8061 1744 8095
rect 1686 8027 1698 8061
rect 1732 8027 1744 8061
rect 1686 8012 1744 8027
rect 1844 8197 1902 8212
rect 1844 8163 1856 8197
rect 1890 8163 1902 8197
rect 1844 8129 1902 8163
rect 1844 8095 1856 8129
rect 1890 8095 1902 8129
rect 1844 8061 1902 8095
rect 1844 8027 1856 8061
rect 1890 8027 1902 8061
rect 1844 8012 1902 8027
rect 2018 8197 2076 8212
rect 2018 8163 2030 8197
rect 2064 8163 2076 8197
rect 2018 8129 2076 8163
rect 2018 8095 2030 8129
rect 2064 8095 2076 8129
rect 2018 8061 2076 8095
rect 2018 8027 2030 8061
rect 2064 8027 2076 8061
rect 2018 8012 2076 8027
rect 2176 8197 2234 8212
rect 2176 8163 2188 8197
rect 2222 8163 2234 8197
rect 2176 8129 2234 8163
rect 2176 8095 2188 8129
rect 2222 8095 2234 8129
rect 2176 8061 2234 8095
rect 2176 8027 2188 8061
rect 2222 8027 2234 8061
rect 2176 8012 2234 8027
rect 2360 8197 2418 8212
rect 2360 8163 2372 8197
rect 2406 8163 2418 8197
rect 2360 8129 2418 8163
rect 2360 8095 2372 8129
rect 2406 8095 2418 8129
rect 2360 8061 2418 8095
rect 2360 8027 2372 8061
rect 2406 8027 2418 8061
rect 2360 8012 2418 8027
rect 2518 8197 2576 8212
rect 2518 8163 2530 8197
rect 2564 8163 2576 8197
rect 2518 8129 2576 8163
rect 2518 8095 2530 8129
rect 2564 8095 2576 8129
rect 2518 8061 2576 8095
rect 2518 8027 2530 8061
rect 2564 8027 2576 8061
rect 2518 8012 2576 8027
rect 2764 8197 2822 8212
rect 2764 8163 2776 8197
rect 2810 8163 2822 8197
rect 2764 8129 2822 8163
rect 2764 8095 2776 8129
rect 2810 8095 2822 8129
rect 2764 8061 2822 8095
rect 2764 8027 2776 8061
rect 2810 8027 2822 8061
rect 2764 8012 2822 8027
rect 2922 8197 2980 8212
rect 2922 8163 2934 8197
rect 2968 8163 2980 8197
rect 2922 8129 2980 8163
rect 2922 8095 2934 8129
rect 2968 8095 2980 8129
rect 2922 8061 2980 8095
rect 2922 8027 2934 8061
rect 2968 8027 2980 8061
rect 2922 8012 2980 8027
rect 3108 8197 3166 8212
rect 3108 8163 3120 8197
rect 3154 8163 3166 8197
rect 3108 8129 3166 8163
rect 3108 8095 3120 8129
rect 3154 8095 3166 8129
rect 3108 8061 3166 8095
rect 3108 8027 3120 8061
rect 3154 8027 3166 8061
rect 3108 8012 3166 8027
rect 3266 8197 3324 8212
rect 3266 8163 3278 8197
rect 3312 8163 3324 8197
rect 3266 8129 3324 8163
rect 3266 8095 3278 8129
rect 3312 8095 3324 8129
rect 3266 8061 3324 8095
rect 3266 8027 3278 8061
rect 3312 8027 3324 8061
rect 3266 8012 3324 8027
rect 3730 8207 3788 8222
rect 3730 8173 3742 8207
rect 3776 8173 3788 8207
rect 3730 8139 3788 8173
rect 3730 8105 3742 8139
rect 3776 8105 3788 8139
rect 3730 8071 3788 8105
rect 3730 8037 3742 8071
rect 3776 8037 3788 8071
rect 3730 8022 3788 8037
rect 3888 8207 3946 8222
rect 3888 8173 3900 8207
rect 3934 8173 3946 8207
rect 3888 8139 3946 8173
rect 3888 8105 3900 8139
rect 3934 8105 3946 8139
rect 3888 8071 3946 8105
rect 3888 8037 3900 8071
rect 3934 8037 3946 8071
rect 3888 8022 3946 8037
rect 4038 8207 4096 8222
rect 4038 8173 4050 8207
rect 4084 8173 4096 8207
rect 4038 8139 4096 8173
rect 4038 8105 4050 8139
rect 4084 8105 4096 8139
rect 4038 8071 4096 8105
rect 4038 8037 4050 8071
rect 4084 8037 4096 8071
rect 4038 8022 4096 8037
rect 4196 8207 4254 8222
rect 4196 8173 4208 8207
rect 4242 8173 4254 8207
rect 4196 8139 4254 8173
rect 4196 8105 4208 8139
rect 4242 8105 4254 8139
rect 4196 8071 4254 8105
rect 4196 8037 4208 8071
rect 4242 8037 4254 8071
rect 4196 8022 4254 8037
rect 4390 8207 4448 8222
rect 4390 8173 4402 8207
rect 4436 8173 4448 8207
rect 4390 8139 4448 8173
rect 4390 8105 4402 8139
rect 4436 8105 4448 8139
rect 4390 8071 4448 8105
rect 4390 8037 4402 8071
rect 4436 8037 4448 8071
rect 4390 8022 4448 8037
rect 4548 8207 4606 8222
rect 4548 8173 4560 8207
rect 4594 8173 4606 8207
rect 4548 8139 4606 8173
rect 4548 8105 4560 8139
rect 4594 8105 4606 8139
rect 4548 8071 4606 8105
rect 4548 8037 4560 8071
rect 4594 8037 4606 8071
rect 4548 8022 4606 8037
rect 4698 8207 4756 8222
rect 4698 8173 4710 8207
rect 4744 8173 4756 8207
rect 4698 8139 4756 8173
rect 4698 8105 4710 8139
rect 4744 8105 4756 8139
rect 4698 8071 4756 8105
rect 4698 8037 4710 8071
rect 4744 8037 4756 8071
rect 4698 8022 4756 8037
rect 4856 8207 4914 8222
rect 4856 8173 4868 8207
rect 4902 8173 4914 8207
rect 4856 8139 4914 8173
rect 4856 8105 4868 8139
rect 4902 8105 4914 8139
rect 4856 8071 4914 8105
rect 4856 8037 4868 8071
rect 4902 8037 4914 8071
rect 4856 8022 4914 8037
rect 5688 8208 5746 8222
rect 5688 8174 5700 8208
rect 5734 8174 5746 8208
rect 5688 8140 5746 8174
rect 5688 8106 5700 8140
rect 5734 8106 5746 8140
rect 5688 8072 5746 8106
rect 5688 8038 5700 8072
rect 5734 8038 5746 8072
rect 5688 8022 5746 8038
rect 5846 8208 5904 8222
rect 5846 8174 5858 8208
rect 5892 8174 5904 8208
rect 5846 8140 5904 8174
rect 5846 8106 5858 8140
rect 5892 8106 5904 8140
rect 5846 8072 5904 8106
rect 5846 8038 5858 8072
rect 5892 8038 5904 8072
rect 5846 8022 5904 8038
rect 5996 8208 6054 8222
rect 5996 8174 6008 8208
rect 6042 8174 6054 8208
rect 5996 8140 6054 8174
rect 5996 8106 6008 8140
rect 6042 8106 6054 8140
rect 5996 8072 6054 8106
rect 5996 8038 6008 8072
rect 6042 8038 6054 8072
rect 5996 8022 6054 8038
rect 6154 8208 6212 8222
rect 6154 8174 6166 8208
rect 6200 8174 6212 8208
rect 6154 8140 6212 8174
rect 6154 8106 6166 8140
rect 6200 8106 6212 8140
rect 6154 8072 6212 8106
rect 6154 8038 6166 8072
rect 6200 8038 6212 8072
rect 6154 8022 6212 8038
rect 6348 8208 6406 8222
rect 6348 8174 6360 8208
rect 6394 8174 6406 8208
rect 6348 8140 6406 8174
rect 6348 8106 6360 8140
rect 6394 8106 6406 8140
rect 6348 8072 6406 8106
rect 6348 8038 6360 8072
rect 6394 8038 6406 8072
rect 6348 8022 6406 8038
rect 6506 8208 6564 8222
rect 6506 8174 6518 8208
rect 6552 8174 6564 8208
rect 6506 8140 6564 8174
rect 6506 8106 6518 8140
rect 6552 8106 6564 8140
rect 6506 8072 6564 8106
rect 6506 8038 6518 8072
rect 6552 8038 6564 8072
rect 6506 8022 6564 8038
rect 6656 8208 6714 8222
rect 6656 8174 6668 8208
rect 6702 8174 6714 8208
rect 6656 8140 6714 8174
rect 6656 8106 6668 8140
rect 6702 8106 6714 8140
rect 6656 8072 6714 8106
rect 6656 8038 6668 8072
rect 6702 8038 6714 8072
rect 6656 8022 6714 8038
rect 6814 8208 6872 8222
rect 6814 8174 6826 8208
rect 6860 8174 6872 8208
rect 6814 8140 6872 8174
rect 6814 8106 6826 8140
rect 6860 8106 6872 8140
rect 6814 8072 6872 8106
rect 6814 8038 6826 8072
rect 6860 8038 6872 8072
rect 6814 8022 6872 8038
rect 1398 6969 1456 6984
rect 1398 6935 1410 6969
rect 1444 6935 1456 6969
rect 1398 6901 1456 6935
rect 1398 6867 1410 6901
rect 1444 6867 1456 6901
rect 1398 6833 1456 6867
rect 1398 6799 1410 6833
rect 1444 6799 1456 6833
rect 1398 6784 1456 6799
rect 1556 6969 1614 6984
rect 1556 6935 1568 6969
rect 1602 6935 1614 6969
rect 1556 6901 1614 6935
rect 1556 6867 1568 6901
rect 1602 6867 1614 6901
rect 1556 6833 1614 6867
rect 1556 6799 1568 6833
rect 1602 6799 1614 6833
rect 1556 6784 1614 6799
rect 1686 6969 1744 6984
rect 1686 6935 1698 6969
rect 1732 6935 1744 6969
rect 1686 6901 1744 6935
rect 1686 6867 1698 6901
rect 1732 6867 1744 6901
rect 1686 6833 1744 6867
rect 1686 6799 1698 6833
rect 1732 6799 1744 6833
rect 1686 6784 1744 6799
rect 1844 6969 1902 6984
rect 1844 6935 1856 6969
rect 1890 6935 1902 6969
rect 1844 6901 1902 6935
rect 1844 6867 1856 6901
rect 1890 6867 1902 6901
rect 1844 6833 1902 6867
rect 1844 6799 1856 6833
rect 1890 6799 1902 6833
rect 1844 6784 1902 6799
rect 2018 6969 2076 6984
rect 2018 6935 2030 6969
rect 2064 6935 2076 6969
rect 2018 6901 2076 6935
rect 2018 6867 2030 6901
rect 2064 6867 2076 6901
rect 2018 6833 2076 6867
rect 2018 6799 2030 6833
rect 2064 6799 2076 6833
rect 2018 6784 2076 6799
rect 2176 6969 2234 6984
rect 2176 6935 2188 6969
rect 2222 6935 2234 6969
rect 2176 6901 2234 6935
rect 2176 6867 2188 6901
rect 2222 6867 2234 6901
rect 2176 6833 2234 6867
rect 2176 6799 2188 6833
rect 2222 6799 2234 6833
rect 2176 6784 2234 6799
rect 2360 6969 2418 6984
rect 2360 6935 2372 6969
rect 2406 6935 2418 6969
rect 2360 6901 2418 6935
rect 2360 6867 2372 6901
rect 2406 6867 2418 6901
rect 2360 6833 2418 6867
rect 2360 6799 2372 6833
rect 2406 6799 2418 6833
rect 2360 6784 2418 6799
rect 2518 6969 2576 6984
rect 2518 6935 2530 6969
rect 2564 6935 2576 6969
rect 2518 6901 2576 6935
rect 2518 6867 2530 6901
rect 2564 6867 2576 6901
rect 2518 6833 2576 6867
rect 2518 6799 2530 6833
rect 2564 6799 2576 6833
rect 2518 6784 2576 6799
rect 2764 6969 2822 6984
rect 2764 6935 2776 6969
rect 2810 6935 2822 6969
rect 2764 6901 2822 6935
rect 2764 6867 2776 6901
rect 2810 6867 2822 6901
rect 2764 6833 2822 6867
rect 2764 6799 2776 6833
rect 2810 6799 2822 6833
rect 2764 6784 2822 6799
rect 2922 6969 2980 6984
rect 2922 6935 2934 6969
rect 2968 6935 2980 6969
rect 2922 6901 2980 6935
rect 2922 6867 2934 6901
rect 2968 6867 2980 6901
rect 2922 6833 2980 6867
rect 2922 6799 2934 6833
rect 2968 6799 2980 6833
rect 2922 6784 2980 6799
rect 3108 6969 3166 6984
rect 3108 6935 3120 6969
rect 3154 6935 3166 6969
rect 3108 6901 3166 6935
rect 3108 6867 3120 6901
rect 3154 6867 3166 6901
rect 3108 6833 3166 6867
rect 3108 6799 3120 6833
rect 3154 6799 3166 6833
rect 3108 6784 3166 6799
rect 3266 6969 3324 6984
rect 3266 6935 3278 6969
rect 3312 6935 3324 6969
rect 3266 6901 3324 6935
rect 3266 6867 3278 6901
rect 3312 6867 3324 6901
rect 3266 6833 3324 6867
rect 3266 6799 3278 6833
rect 3312 6799 3324 6833
rect 3266 6784 3324 6799
rect 3730 6979 3788 6994
rect 3730 6945 3742 6979
rect 3776 6945 3788 6979
rect 3730 6911 3788 6945
rect 3730 6877 3742 6911
rect 3776 6877 3788 6911
rect 3730 6843 3788 6877
rect 3730 6809 3742 6843
rect 3776 6809 3788 6843
rect 3730 6794 3788 6809
rect 3888 6979 3946 6994
rect 3888 6945 3900 6979
rect 3934 6945 3946 6979
rect 3888 6911 3946 6945
rect 3888 6877 3900 6911
rect 3934 6877 3946 6911
rect 3888 6843 3946 6877
rect 3888 6809 3900 6843
rect 3934 6809 3946 6843
rect 3888 6794 3946 6809
rect 4038 6979 4096 6994
rect 4038 6945 4050 6979
rect 4084 6945 4096 6979
rect 4038 6911 4096 6945
rect 4038 6877 4050 6911
rect 4084 6877 4096 6911
rect 4038 6843 4096 6877
rect 4038 6809 4050 6843
rect 4084 6809 4096 6843
rect 4038 6794 4096 6809
rect 4196 6979 4254 6994
rect 4196 6945 4208 6979
rect 4242 6945 4254 6979
rect 4196 6911 4254 6945
rect 4196 6877 4208 6911
rect 4242 6877 4254 6911
rect 4196 6843 4254 6877
rect 4196 6809 4208 6843
rect 4242 6809 4254 6843
rect 4196 6794 4254 6809
rect 4390 6979 4448 6994
rect 4390 6945 4402 6979
rect 4436 6945 4448 6979
rect 4390 6911 4448 6945
rect 4390 6877 4402 6911
rect 4436 6877 4448 6911
rect 4390 6843 4448 6877
rect 4390 6809 4402 6843
rect 4436 6809 4448 6843
rect 4390 6794 4448 6809
rect 4548 6979 4606 6994
rect 4548 6945 4560 6979
rect 4594 6945 4606 6979
rect 4548 6911 4606 6945
rect 4548 6877 4560 6911
rect 4594 6877 4606 6911
rect 4548 6843 4606 6877
rect 4548 6809 4560 6843
rect 4594 6809 4606 6843
rect 4548 6794 4606 6809
rect 4698 6979 4756 6994
rect 4698 6945 4710 6979
rect 4744 6945 4756 6979
rect 4698 6911 4756 6945
rect 4698 6877 4710 6911
rect 4744 6877 4756 6911
rect 4698 6843 4756 6877
rect 4698 6809 4710 6843
rect 4744 6809 4756 6843
rect 4698 6794 4756 6809
rect 4856 6979 4914 6994
rect 4856 6945 4868 6979
rect 4902 6945 4914 6979
rect 4856 6911 4914 6945
rect 4856 6877 4868 6911
rect 4902 6877 4914 6911
rect 4856 6843 4914 6877
rect 4856 6809 4868 6843
rect 4902 6809 4914 6843
rect 4856 6794 4914 6809
rect 5688 6980 5746 6994
rect 5688 6946 5700 6980
rect 5734 6946 5746 6980
rect 5688 6912 5746 6946
rect 5688 6878 5700 6912
rect 5734 6878 5746 6912
rect 5688 6844 5746 6878
rect 5688 6810 5700 6844
rect 5734 6810 5746 6844
rect 5688 6794 5746 6810
rect 5846 6980 5904 6994
rect 5846 6946 5858 6980
rect 5892 6946 5904 6980
rect 5846 6912 5904 6946
rect 5846 6878 5858 6912
rect 5892 6878 5904 6912
rect 5846 6844 5904 6878
rect 5846 6810 5858 6844
rect 5892 6810 5904 6844
rect 5846 6794 5904 6810
rect 5996 6980 6054 6994
rect 5996 6946 6008 6980
rect 6042 6946 6054 6980
rect 5996 6912 6054 6946
rect 5996 6878 6008 6912
rect 6042 6878 6054 6912
rect 5996 6844 6054 6878
rect 5996 6810 6008 6844
rect 6042 6810 6054 6844
rect 5996 6794 6054 6810
rect 6154 6980 6212 6994
rect 6154 6946 6166 6980
rect 6200 6946 6212 6980
rect 6154 6912 6212 6946
rect 6154 6878 6166 6912
rect 6200 6878 6212 6912
rect 6154 6844 6212 6878
rect 6154 6810 6166 6844
rect 6200 6810 6212 6844
rect 6154 6794 6212 6810
rect 6348 6980 6406 6994
rect 6348 6946 6360 6980
rect 6394 6946 6406 6980
rect 6348 6912 6406 6946
rect 6348 6878 6360 6912
rect 6394 6878 6406 6912
rect 6348 6844 6406 6878
rect 6348 6810 6360 6844
rect 6394 6810 6406 6844
rect 6348 6794 6406 6810
rect 6506 6980 6564 6994
rect 6506 6946 6518 6980
rect 6552 6946 6564 6980
rect 6506 6912 6564 6946
rect 6506 6878 6518 6912
rect 6552 6878 6564 6912
rect 6506 6844 6564 6878
rect 6506 6810 6518 6844
rect 6552 6810 6564 6844
rect 6506 6794 6564 6810
rect 6656 6980 6714 6994
rect 6656 6946 6668 6980
rect 6702 6946 6714 6980
rect 6656 6912 6714 6946
rect 6656 6878 6668 6912
rect 6702 6878 6714 6912
rect 6656 6844 6714 6878
rect 6656 6810 6668 6844
rect 6702 6810 6714 6844
rect 6656 6794 6714 6810
rect 6814 6980 6872 6994
rect 6814 6946 6826 6980
rect 6860 6946 6872 6980
rect 6814 6912 6872 6946
rect 6814 6878 6826 6912
rect 6860 6878 6872 6912
rect 6814 6844 6872 6878
rect 6814 6810 6826 6844
rect 6860 6810 6872 6844
rect 6814 6794 6872 6810
rect 1398 5741 1456 5756
rect 1398 5707 1410 5741
rect 1444 5707 1456 5741
rect 1398 5673 1456 5707
rect 1398 5639 1410 5673
rect 1444 5639 1456 5673
rect 1398 5605 1456 5639
rect 1398 5571 1410 5605
rect 1444 5571 1456 5605
rect 1398 5556 1456 5571
rect 1556 5741 1614 5756
rect 1556 5707 1568 5741
rect 1602 5707 1614 5741
rect 1556 5673 1614 5707
rect 1556 5639 1568 5673
rect 1602 5639 1614 5673
rect 1556 5605 1614 5639
rect 1556 5571 1568 5605
rect 1602 5571 1614 5605
rect 1556 5556 1614 5571
rect 1686 5741 1744 5756
rect 1686 5707 1698 5741
rect 1732 5707 1744 5741
rect 1686 5673 1744 5707
rect 1686 5639 1698 5673
rect 1732 5639 1744 5673
rect 1686 5605 1744 5639
rect 1686 5571 1698 5605
rect 1732 5571 1744 5605
rect 1686 5556 1744 5571
rect 1844 5741 1902 5756
rect 1844 5707 1856 5741
rect 1890 5707 1902 5741
rect 1844 5673 1902 5707
rect 1844 5639 1856 5673
rect 1890 5639 1902 5673
rect 1844 5605 1902 5639
rect 1844 5571 1856 5605
rect 1890 5571 1902 5605
rect 1844 5556 1902 5571
rect 2018 5741 2076 5756
rect 2018 5707 2030 5741
rect 2064 5707 2076 5741
rect 2018 5673 2076 5707
rect 2018 5639 2030 5673
rect 2064 5639 2076 5673
rect 2018 5605 2076 5639
rect 2018 5571 2030 5605
rect 2064 5571 2076 5605
rect 2018 5556 2076 5571
rect 2176 5741 2234 5756
rect 2176 5707 2188 5741
rect 2222 5707 2234 5741
rect 2176 5673 2234 5707
rect 2176 5639 2188 5673
rect 2222 5639 2234 5673
rect 2176 5605 2234 5639
rect 2176 5571 2188 5605
rect 2222 5571 2234 5605
rect 2176 5556 2234 5571
rect 2360 5741 2418 5756
rect 2360 5707 2372 5741
rect 2406 5707 2418 5741
rect 2360 5673 2418 5707
rect 2360 5639 2372 5673
rect 2406 5639 2418 5673
rect 2360 5605 2418 5639
rect 2360 5571 2372 5605
rect 2406 5571 2418 5605
rect 2360 5556 2418 5571
rect 2518 5741 2576 5756
rect 2518 5707 2530 5741
rect 2564 5707 2576 5741
rect 2518 5673 2576 5707
rect 2518 5639 2530 5673
rect 2564 5639 2576 5673
rect 2518 5605 2576 5639
rect 2518 5571 2530 5605
rect 2564 5571 2576 5605
rect 2518 5556 2576 5571
rect 2764 5741 2822 5756
rect 2764 5707 2776 5741
rect 2810 5707 2822 5741
rect 2764 5673 2822 5707
rect 2764 5639 2776 5673
rect 2810 5639 2822 5673
rect 2764 5605 2822 5639
rect 2764 5571 2776 5605
rect 2810 5571 2822 5605
rect 2764 5556 2822 5571
rect 2922 5741 2980 5756
rect 2922 5707 2934 5741
rect 2968 5707 2980 5741
rect 2922 5673 2980 5707
rect 2922 5639 2934 5673
rect 2968 5639 2980 5673
rect 2922 5605 2980 5639
rect 2922 5571 2934 5605
rect 2968 5571 2980 5605
rect 2922 5556 2980 5571
rect 3108 5741 3166 5756
rect 3108 5707 3120 5741
rect 3154 5707 3166 5741
rect 3108 5673 3166 5707
rect 3108 5639 3120 5673
rect 3154 5639 3166 5673
rect 3108 5605 3166 5639
rect 3108 5571 3120 5605
rect 3154 5571 3166 5605
rect 3108 5556 3166 5571
rect 3266 5741 3324 5756
rect 3266 5707 3278 5741
rect 3312 5707 3324 5741
rect 3266 5673 3324 5707
rect 3266 5639 3278 5673
rect 3312 5639 3324 5673
rect 3266 5605 3324 5639
rect 3266 5571 3278 5605
rect 3312 5571 3324 5605
rect 3266 5556 3324 5571
rect 3730 5751 3788 5766
rect 3730 5717 3742 5751
rect 3776 5717 3788 5751
rect 3730 5683 3788 5717
rect 3730 5649 3742 5683
rect 3776 5649 3788 5683
rect 3730 5615 3788 5649
rect 3730 5581 3742 5615
rect 3776 5581 3788 5615
rect 3730 5566 3788 5581
rect 3888 5751 3946 5766
rect 3888 5717 3900 5751
rect 3934 5717 3946 5751
rect 3888 5683 3946 5717
rect 3888 5649 3900 5683
rect 3934 5649 3946 5683
rect 3888 5615 3946 5649
rect 3888 5581 3900 5615
rect 3934 5581 3946 5615
rect 3888 5566 3946 5581
rect 4038 5751 4096 5766
rect 4038 5717 4050 5751
rect 4084 5717 4096 5751
rect 4038 5683 4096 5717
rect 4038 5649 4050 5683
rect 4084 5649 4096 5683
rect 4038 5615 4096 5649
rect 4038 5581 4050 5615
rect 4084 5581 4096 5615
rect 4038 5566 4096 5581
rect 4196 5751 4254 5766
rect 4196 5717 4208 5751
rect 4242 5717 4254 5751
rect 4196 5683 4254 5717
rect 4196 5649 4208 5683
rect 4242 5649 4254 5683
rect 4196 5615 4254 5649
rect 4196 5581 4208 5615
rect 4242 5581 4254 5615
rect 4196 5566 4254 5581
rect 4390 5751 4448 5766
rect 4390 5717 4402 5751
rect 4436 5717 4448 5751
rect 4390 5683 4448 5717
rect 4390 5649 4402 5683
rect 4436 5649 4448 5683
rect 4390 5615 4448 5649
rect 4390 5581 4402 5615
rect 4436 5581 4448 5615
rect 4390 5566 4448 5581
rect 4548 5751 4606 5766
rect 4548 5717 4560 5751
rect 4594 5717 4606 5751
rect 4548 5683 4606 5717
rect 4548 5649 4560 5683
rect 4594 5649 4606 5683
rect 4548 5615 4606 5649
rect 4548 5581 4560 5615
rect 4594 5581 4606 5615
rect 4548 5566 4606 5581
rect 4698 5751 4756 5766
rect 4698 5717 4710 5751
rect 4744 5717 4756 5751
rect 4698 5683 4756 5717
rect 4698 5649 4710 5683
rect 4744 5649 4756 5683
rect 4698 5615 4756 5649
rect 4698 5581 4710 5615
rect 4744 5581 4756 5615
rect 4698 5566 4756 5581
rect 4856 5751 4914 5766
rect 4856 5717 4868 5751
rect 4902 5717 4914 5751
rect 4856 5683 4914 5717
rect 4856 5649 4868 5683
rect 4902 5649 4914 5683
rect 4856 5615 4914 5649
rect 4856 5581 4868 5615
rect 4902 5581 4914 5615
rect 4856 5566 4914 5581
rect 5688 5752 5746 5766
rect 5688 5718 5700 5752
rect 5734 5718 5746 5752
rect 5688 5684 5746 5718
rect 5688 5650 5700 5684
rect 5734 5650 5746 5684
rect 5688 5616 5746 5650
rect 5688 5582 5700 5616
rect 5734 5582 5746 5616
rect 5688 5566 5746 5582
rect 5846 5752 5904 5766
rect 5846 5718 5858 5752
rect 5892 5718 5904 5752
rect 5846 5684 5904 5718
rect 5846 5650 5858 5684
rect 5892 5650 5904 5684
rect 5846 5616 5904 5650
rect 5846 5582 5858 5616
rect 5892 5582 5904 5616
rect 5846 5566 5904 5582
rect 5996 5752 6054 5766
rect 5996 5718 6008 5752
rect 6042 5718 6054 5752
rect 5996 5684 6054 5718
rect 5996 5650 6008 5684
rect 6042 5650 6054 5684
rect 5996 5616 6054 5650
rect 5996 5582 6008 5616
rect 6042 5582 6054 5616
rect 5996 5566 6054 5582
rect 6154 5752 6212 5766
rect 6154 5718 6166 5752
rect 6200 5718 6212 5752
rect 6154 5684 6212 5718
rect 6154 5650 6166 5684
rect 6200 5650 6212 5684
rect 6154 5616 6212 5650
rect 6154 5582 6166 5616
rect 6200 5582 6212 5616
rect 6154 5566 6212 5582
rect 6348 5752 6406 5766
rect 6348 5718 6360 5752
rect 6394 5718 6406 5752
rect 6348 5684 6406 5718
rect 6348 5650 6360 5684
rect 6394 5650 6406 5684
rect 6348 5616 6406 5650
rect 6348 5582 6360 5616
rect 6394 5582 6406 5616
rect 6348 5566 6406 5582
rect 6506 5752 6564 5766
rect 6506 5718 6518 5752
rect 6552 5718 6564 5752
rect 6506 5684 6564 5718
rect 6506 5650 6518 5684
rect 6552 5650 6564 5684
rect 6506 5616 6564 5650
rect 6506 5582 6518 5616
rect 6552 5582 6564 5616
rect 6506 5566 6564 5582
rect 6656 5752 6714 5766
rect 6656 5718 6668 5752
rect 6702 5718 6714 5752
rect 6656 5684 6714 5718
rect 6656 5650 6668 5684
rect 6702 5650 6714 5684
rect 6656 5616 6714 5650
rect 6656 5582 6668 5616
rect 6702 5582 6714 5616
rect 6656 5566 6714 5582
rect 6814 5752 6872 5766
rect 6814 5718 6826 5752
rect 6860 5718 6872 5752
rect 6814 5684 6872 5718
rect 6814 5650 6826 5684
rect 6860 5650 6872 5684
rect 6814 5616 6872 5650
rect 6814 5582 6826 5616
rect 6860 5582 6872 5616
rect 6814 5566 6872 5582
rect 1398 4513 1456 4528
rect 1398 4479 1410 4513
rect 1444 4479 1456 4513
rect 1398 4445 1456 4479
rect 1398 4411 1410 4445
rect 1444 4411 1456 4445
rect 1398 4377 1456 4411
rect 1398 4343 1410 4377
rect 1444 4343 1456 4377
rect 1398 4328 1456 4343
rect 1556 4513 1614 4528
rect 1556 4479 1568 4513
rect 1602 4479 1614 4513
rect 1556 4445 1614 4479
rect 1556 4411 1568 4445
rect 1602 4411 1614 4445
rect 1556 4377 1614 4411
rect 1556 4343 1568 4377
rect 1602 4343 1614 4377
rect 1556 4328 1614 4343
rect 1686 4513 1744 4528
rect 1686 4479 1698 4513
rect 1732 4479 1744 4513
rect 1686 4445 1744 4479
rect 1686 4411 1698 4445
rect 1732 4411 1744 4445
rect 1686 4377 1744 4411
rect 1686 4343 1698 4377
rect 1732 4343 1744 4377
rect 1686 4328 1744 4343
rect 1844 4513 1902 4528
rect 1844 4479 1856 4513
rect 1890 4479 1902 4513
rect 1844 4445 1902 4479
rect 1844 4411 1856 4445
rect 1890 4411 1902 4445
rect 1844 4377 1902 4411
rect 1844 4343 1856 4377
rect 1890 4343 1902 4377
rect 1844 4328 1902 4343
rect 2018 4513 2076 4528
rect 2018 4479 2030 4513
rect 2064 4479 2076 4513
rect 2018 4445 2076 4479
rect 2018 4411 2030 4445
rect 2064 4411 2076 4445
rect 2018 4377 2076 4411
rect 2018 4343 2030 4377
rect 2064 4343 2076 4377
rect 2018 4328 2076 4343
rect 2176 4513 2234 4528
rect 2176 4479 2188 4513
rect 2222 4479 2234 4513
rect 2176 4445 2234 4479
rect 2176 4411 2188 4445
rect 2222 4411 2234 4445
rect 2176 4377 2234 4411
rect 2176 4343 2188 4377
rect 2222 4343 2234 4377
rect 2176 4328 2234 4343
rect 2360 4513 2418 4528
rect 2360 4479 2372 4513
rect 2406 4479 2418 4513
rect 2360 4445 2418 4479
rect 2360 4411 2372 4445
rect 2406 4411 2418 4445
rect 2360 4377 2418 4411
rect 2360 4343 2372 4377
rect 2406 4343 2418 4377
rect 2360 4328 2418 4343
rect 2518 4513 2576 4528
rect 2518 4479 2530 4513
rect 2564 4479 2576 4513
rect 2518 4445 2576 4479
rect 2518 4411 2530 4445
rect 2564 4411 2576 4445
rect 2518 4377 2576 4411
rect 2518 4343 2530 4377
rect 2564 4343 2576 4377
rect 2518 4328 2576 4343
rect 2764 4513 2822 4528
rect 2764 4479 2776 4513
rect 2810 4479 2822 4513
rect 2764 4445 2822 4479
rect 2764 4411 2776 4445
rect 2810 4411 2822 4445
rect 2764 4377 2822 4411
rect 2764 4343 2776 4377
rect 2810 4343 2822 4377
rect 2764 4328 2822 4343
rect 2922 4513 2980 4528
rect 2922 4479 2934 4513
rect 2968 4479 2980 4513
rect 2922 4445 2980 4479
rect 2922 4411 2934 4445
rect 2968 4411 2980 4445
rect 2922 4377 2980 4411
rect 2922 4343 2934 4377
rect 2968 4343 2980 4377
rect 2922 4328 2980 4343
rect 3108 4513 3166 4528
rect 3108 4479 3120 4513
rect 3154 4479 3166 4513
rect 3108 4445 3166 4479
rect 3108 4411 3120 4445
rect 3154 4411 3166 4445
rect 3108 4377 3166 4411
rect 3108 4343 3120 4377
rect 3154 4343 3166 4377
rect 3108 4328 3166 4343
rect 3266 4513 3324 4528
rect 3266 4479 3278 4513
rect 3312 4479 3324 4513
rect 3266 4445 3324 4479
rect 3266 4411 3278 4445
rect 3312 4411 3324 4445
rect 3266 4377 3324 4411
rect 3266 4343 3278 4377
rect 3312 4343 3324 4377
rect 3266 4328 3324 4343
rect 3730 4523 3788 4538
rect 3730 4489 3742 4523
rect 3776 4489 3788 4523
rect 3730 4455 3788 4489
rect 3730 4421 3742 4455
rect 3776 4421 3788 4455
rect 3730 4387 3788 4421
rect 3730 4353 3742 4387
rect 3776 4353 3788 4387
rect 3730 4338 3788 4353
rect 3888 4523 3946 4538
rect 3888 4489 3900 4523
rect 3934 4489 3946 4523
rect 3888 4455 3946 4489
rect 3888 4421 3900 4455
rect 3934 4421 3946 4455
rect 3888 4387 3946 4421
rect 3888 4353 3900 4387
rect 3934 4353 3946 4387
rect 3888 4338 3946 4353
rect 4038 4523 4096 4538
rect 4038 4489 4050 4523
rect 4084 4489 4096 4523
rect 4038 4455 4096 4489
rect 4038 4421 4050 4455
rect 4084 4421 4096 4455
rect 4038 4387 4096 4421
rect 4038 4353 4050 4387
rect 4084 4353 4096 4387
rect 4038 4338 4096 4353
rect 4196 4523 4254 4538
rect 4196 4489 4208 4523
rect 4242 4489 4254 4523
rect 4196 4455 4254 4489
rect 4196 4421 4208 4455
rect 4242 4421 4254 4455
rect 4196 4387 4254 4421
rect 4196 4353 4208 4387
rect 4242 4353 4254 4387
rect 4196 4338 4254 4353
rect 4390 4523 4448 4538
rect 4390 4489 4402 4523
rect 4436 4489 4448 4523
rect 4390 4455 4448 4489
rect 4390 4421 4402 4455
rect 4436 4421 4448 4455
rect 4390 4387 4448 4421
rect 4390 4353 4402 4387
rect 4436 4353 4448 4387
rect 4390 4338 4448 4353
rect 4548 4523 4606 4538
rect 4548 4489 4560 4523
rect 4594 4489 4606 4523
rect 4548 4455 4606 4489
rect 4548 4421 4560 4455
rect 4594 4421 4606 4455
rect 4548 4387 4606 4421
rect 4548 4353 4560 4387
rect 4594 4353 4606 4387
rect 4548 4338 4606 4353
rect 4698 4523 4756 4538
rect 4698 4489 4710 4523
rect 4744 4489 4756 4523
rect 4698 4455 4756 4489
rect 4698 4421 4710 4455
rect 4744 4421 4756 4455
rect 4698 4387 4756 4421
rect 4698 4353 4710 4387
rect 4744 4353 4756 4387
rect 4698 4338 4756 4353
rect 4856 4523 4914 4538
rect 4856 4489 4868 4523
rect 4902 4489 4914 4523
rect 4856 4455 4914 4489
rect 4856 4421 4868 4455
rect 4902 4421 4914 4455
rect 4856 4387 4914 4421
rect 4856 4353 4868 4387
rect 4902 4353 4914 4387
rect 4856 4338 4914 4353
rect 5688 4524 5746 4538
rect 5688 4490 5700 4524
rect 5734 4490 5746 4524
rect 5688 4456 5746 4490
rect 5688 4422 5700 4456
rect 5734 4422 5746 4456
rect 5688 4388 5746 4422
rect 5688 4354 5700 4388
rect 5734 4354 5746 4388
rect 5688 4338 5746 4354
rect 5846 4524 5904 4538
rect 5846 4490 5858 4524
rect 5892 4490 5904 4524
rect 5846 4456 5904 4490
rect 5846 4422 5858 4456
rect 5892 4422 5904 4456
rect 5846 4388 5904 4422
rect 5846 4354 5858 4388
rect 5892 4354 5904 4388
rect 5846 4338 5904 4354
rect 5996 4524 6054 4538
rect 5996 4490 6008 4524
rect 6042 4490 6054 4524
rect 5996 4456 6054 4490
rect 5996 4422 6008 4456
rect 6042 4422 6054 4456
rect 5996 4388 6054 4422
rect 5996 4354 6008 4388
rect 6042 4354 6054 4388
rect 5996 4338 6054 4354
rect 6154 4524 6212 4538
rect 6154 4490 6166 4524
rect 6200 4490 6212 4524
rect 6154 4456 6212 4490
rect 6154 4422 6166 4456
rect 6200 4422 6212 4456
rect 6154 4388 6212 4422
rect 6154 4354 6166 4388
rect 6200 4354 6212 4388
rect 6154 4338 6212 4354
rect 6348 4524 6406 4538
rect 6348 4490 6360 4524
rect 6394 4490 6406 4524
rect 6348 4456 6406 4490
rect 6348 4422 6360 4456
rect 6394 4422 6406 4456
rect 6348 4388 6406 4422
rect 6348 4354 6360 4388
rect 6394 4354 6406 4388
rect 6348 4338 6406 4354
rect 6506 4524 6564 4538
rect 6506 4490 6518 4524
rect 6552 4490 6564 4524
rect 6506 4456 6564 4490
rect 6506 4422 6518 4456
rect 6552 4422 6564 4456
rect 6506 4388 6564 4422
rect 6506 4354 6518 4388
rect 6552 4354 6564 4388
rect 6506 4338 6564 4354
rect 6656 4524 6714 4538
rect 6656 4490 6668 4524
rect 6702 4490 6714 4524
rect 6656 4456 6714 4490
rect 6656 4422 6668 4456
rect 6702 4422 6714 4456
rect 6656 4388 6714 4422
rect 6656 4354 6668 4388
rect 6702 4354 6714 4388
rect 6656 4338 6714 4354
rect 6814 4524 6872 4538
rect 6814 4490 6826 4524
rect 6860 4490 6872 4524
rect 6814 4456 6872 4490
rect 6814 4422 6826 4456
rect 6860 4422 6872 4456
rect 6814 4388 6872 4422
rect 6814 4354 6826 4388
rect 6860 4354 6872 4388
rect 6814 4338 6872 4354
rect 1398 3285 1456 3300
rect 1398 3251 1410 3285
rect 1444 3251 1456 3285
rect 1398 3217 1456 3251
rect 1398 3183 1410 3217
rect 1444 3183 1456 3217
rect 1398 3149 1456 3183
rect 1398 3115 1410 3149
rect 1444 3115 1456 3149
rect 1398 3100 1456 3115
rect 1556 3285 1614 3300
rect 1556 3251 1568 3285
rect 1602 3251 1614 3285
rect 1556 3217 1614 3251
rect 1556 3183 1568 3217
rect 1602 3183 1614 3217
rect 1556 3149 1614 3183
rect 1556 3115 1568 3149
rect 1602 3115 1614 3149
rect 1556 3100 1614 3115
rect 1686 3285 1744 3300
rect 1686 3251 1698 3285
rect 1732 3251 1744 3285
rect 1686 3217 1744 3251
rect 1686 3183 1698 3217
rect 1732 3183 1744 3217
rect 1686 3149 1744 3183
rect 1686 3115 1698 3149
rect 1732 3115 1744 3149
rect 1686 3100 1744 3115
rect 1844 3285 1902 3300
rect 1844 3251 1856 3285
rect 1890 3251 1902 3285
rect 1844 3217 1902 3251
rect 1844 3183 1856 3217
rect 1890 3183 1902 3217
rect 1844 3149 1902 3183
rect 1844 3115 1856 3149
rect 1890 3115 1902 3149
rect 1844 3100 1902 3115
rect 2018 3285 2076 3300
rect 2018 3251 2030 3285
rect 2064 3251 2076 3285
rect 2018 3217 2076 3251
rect 2018 3183 2030 3217
rect 2064 3183 2076 3217
rect 2018 3149 2076 3183
rect 2018 3115 2030 3149
rect 2064 3115 2076 3149
rect 2018 3100 2076 3115
rect 2176 3285 2234 3300
rect 2176 3251 2188 3285
rect 2222 3251 2234 3285
rect 2176 3217 2234 3251
rect 2176 3183 2188 3217
rect 2222 3183 2234 3217
rect 2176 3149 2234 3183
rect 2176 3115 2188 3149
rect 2222 3115 2234 3149
rect 2176 3100 2234 3115
rect 2360 3285 2418 3300
rect 2360 3251 2372 3285
rect 2406 3251 2418 3285
rect 2360 3217 2418 3251
rect 2360 3183 2372 3217
rect 2406 3183 2418 3217
rect 2360 3149 2418 3183
rect 2360 3115 2372 3149
rect 2406 3115 2418 3149
rect 2360 3100 2418 3115
rect 2518 3285 2576 3300
rect 2518 3251 2530 3285
rect 2564 3251 2576 3285
rect 2518 3217 2576 3251
rect 2518 3183 2530 3217
rect 2564 3183 2576 3217
rect 2518 3149 2576 3183
rect 2518 3115 2530 3149
rect 2564 3115 2576 3149
rect 2518 3100 2576 3115
rect 2764 3285 2822 3300
rect 2764 3251 2776 3285
rect 2810 3251 2822 3285
rect 2764 3217 2822 3251
rect 2764 3183 2776 3217
rect 2810 3183 2822 3217
rect 2764 3149 2822 3183
rect 2764 3115 2776 3149
rect 2810 3115 2822 3149
rect 2764 3100 2822 3115
rect 2922 3285 2980 3300
rect 2922 3251 2934 3285
rect 2968 3251 2980 3285
rect 2922 3217 2980 3251
rect 2922 3183 2934 3217
rect 2968 3183 2980 3217
rect 2922 3149 2980 3183
rect 2922 3115 2934 3149
rect 2968 3115 2980 3149
rect 2922 3100 2980 3115
rect 3108 3285 3166 3300
rect 3108 3251 3120 3285
rect 3154 3251 3166 3285
rect 3108 3217 3166 3251
rect 3108 3183 3120 3217
rect 3154 3183 3166 3217
rect 3108 3149 3166 3183
rect 3108 3115 3120 3149
rect 3154 3115 3166 3149
rect 3108 3100 3166 3115
rect 3266 3285 3324 3300
rect 3266 3251 3278 3285
rect 3312 3251 3324 3285
rect 3266 3217 3324 3251
rect 3266 3183 3278 3217
rect 3312 3183 3324 3217
rect 3266 3149 3324 3183
rect 3266 3115 3278 3149
rect 3312 3115 3324 3149
rect 3266 3100 3324 3115
rect 3730 3295 3788 3310
rect 3730 3261 3742 3295
rect 3776 3261 3788 3295
rect 3730 3227 3788 3261
rect 3730 3193 3742 3227
rect 3776 3193 3788 3227
rect 3730 3159 3788 3193
rect 3730 3125 3742 3159
rect 3776 3125 3788 3159
rect 3730 3110 3788 3125
rect 3888 3295 3946 3310
rect 3888 3261 3900 3295
rect 3934 3261 3946 3295
rect 3888 3227 3946 3261
rect 3888 3193 3900 3227
rect 3934 3193 3946 3227
rect 3888 3159 3946 3193
rect 3888 3125 3900 3159
rect 3934 3125 3946 3159
rect 3888 3110 3946 3125
rect 4038 3295 4096 3310
rect 4038 3261 4050 3295
rect 4084 3261 4096 3295
rect 4038 3227 4096 3261
rect 4038 3193 4050 3227
rect 4084 3193 4096 3227
rect 4038 3159 4096 3193
rect 4038 3125 4050 3159
rect 4084 3125 4096 3159
rect 4038 3110 4096 3125
rect 4196 3295 4254 3310
rect 4196 3261 4208 3295
rect 4242 3261 4254 3295
rect 4196 3227 4254 3261
rect 4196 3193 4208 3227
rect 4242 3193 4254 3227
rect 4196 3159 4254 3193
rect 4196 3125 4208 3159
rect 4242 3125 4254 3159
rect 4196 3110 4254 3125
rect 4390 3295 4448 3310
rect 4390 3261 4402 3295
rect 4436 3261 4448 3295
rect 4390 3227 4448 3261
rect 4390 3193 4402 3227
rect 4436 3193 4448 3227
rect 4390 3159 4448 3193
rect 4390 3125 4402 3159
rect 4436 3125 4448 3159
rect 4390 3110 4448 3125
rect 4548 3295 4606 3310
rect 4548 3261 4560 3295
rect 4594 3261 4606 3295
rect 4548 3227 4606 3261
rect 4548 3193 4560 3227
rect 4594 3193 4606 3227
rect 4548 3159 4606 3193
rect 4548 3125 4560 3159
rect 4594 3125 4606 3159
rect 4548 3110 4606 3125
rect 4698 3295 4756 3310
rect 4698 3261 4710 3295
rect 4744 3261 4756 3295
rect 4698 3227 4756 3261
rect 4698 3193 4710 3227
rect 4744 3193 4756 3227
rect 4698 3159 4756 3193
rect 4698 3125 4710 3159
rect 4744 3125 4756 3159
rect 4698 3110 4756 3125
rect 4856 3295 4914 3310
rect 4856 3261 4868 3295
rect 4902 3261 4914 3295
rect 4856 3227 4914 3261
rect 4856 3193 4868 3227
rect 4902 3193 4914 3227
rect 4856 3159 4914 3193
rect 4856 3125 4868 3159
rect 4902 3125 4914 3159
rect 4856 3110 4914 3125
rect 5688 3296 5746 3310
rect 5688 3262 5700 3296
rect 5734 3262 5746 3296
rect 5688 3228 5746 3262
rect 5688 3194 5700 3228
rect 5734 3194 5746 3228
rect 5688 3160 5746 3194
rect 5688 3126 5700 3160
rect 5734 3126 5746 3160
rect 5688 3110 5746 3126
rect 5846 3296 5904 3310
rect 5846 3262 5858 3296
rect 5892 3262 5904 3296
rect 5846 3228 5904 3262
rect 5846 3194 5858 3228
rect 5892 3194 5904 3228
rect 5846 3160 5904 3194
rect 5846 3126 5858 3160
rect 5892 3126 5904 3160
rect 5846 3110 5904 3126
rect 5996 3296 6054 3310
rect 5996 3262 6008 3296
rect 6042 3262 6054 3296
rect 5996 3228 6054 3262
rect 5996 3194 6008 3228
rect 6042 3194 6054 3228
rect 5996 3160 6054 3194
rect 5996 3126 6008 3160
rect 6042 3126 6054 3160
rect 5996 3110 6054 3126
rect 6154 3296 6212 3310
rect 6154 3262 6166 3296
rect 6200 3262 6212 3296
rect 6154 3228 6212 3262
rect 6154 3194 6166 3228
rect 6200 3194 6212 3228
rect 6154 3160 6212 3194
rect 6154 3126 6166 3160
rect 6200 3126 6212 3160
rect 6154 3110 6212 3126
rect 6348 3296 6406 3310
rect 6348 3262 6360 3296
rect 6394 3262 6406 3296
rect 6348 3228 6406 3262
rect 6348 3194 6360 3228
rect 6394 3194 6406 3228
rect 6348 3160 6406 3194
rect 6348 3126 6360 3160
rect 6394 3126 6406 3160
rect 6348 3110 6406 3126
rect 6506 3296 6564 3310
rect 6506 3262 6518 3296
rect 6552 3262 6564 3296
rect 6506 3228 6564 3262
rect 6506 3194 6518 3228
rect 6552 3194 6564 3228
rect 6506 3160 6564 3194
rect 6506 3126 6518 3160
rect 6552 3126 6564 3160
rect 6506 3110 6564 3126
rect 6656 3296 6714 3310
rect 6656 3262 6668 3296
rect 6702 3262 6714 3296
rect 6656 3228 6714 3262
rect 6656 3194 6668 3228
rect 6702 3194 6714 3228
rect 6656 3160 6714 3194
rect 6656 3126 6668 3160
rect 6702 3126 6714 3160
rect 6656 3110 6714 3126
rect 6814 3296 6872 3310
rect 6814 3262 6826 3296
rect 6860 3262 6872 3296
rect 6814 3228 6872 3262
rect 6814 3194 6826 3228
rect 6860 3194 6872 3228
rect 6814 3160 6872 3194
rect 6814 3126 6826 3160
rect 6860 3126 6872 3160
rect 6814 3110 6872 3126
rect 1398 2057 1456 2072
rect 1398 2023 1410 2057
rect 1444 2023 1456 2057
rect 1398 1989 1456 2023
rect 1398 1955 1410 1989
rect 1444 1955 1456 1989
rect 1398 1921 1456 1955
rect 1398 1887 1410 1921
rect 1444 1887 1456 1921
rect 1398 1872 1456 1887
rect 1556 2057 1614 2072
rect 1556 2023 1568 2057
rect 1602 2023 1614 2057
rect 1556 1989 1614 2023
rect 1556 1955 1568 1989
rect 1602 1955 1614 1989
rect 1556 1921 1614 1955
rect 1556 1887 1568 1921
rect 1602 1887 1614 1921
rect 1556 1872 1614 1887
rect 1686 2057 1744 2072
rect 1686 2023 1698 2057
rect 1732 2023 1744 2057
rect 1686 1989 1744 2023
rect 1686 1955 1698 1989
rect 1732 1955 1744 1989
rect 1686 1921 1744 1955
rect 1686 1887 1698 1921
rect 1732 1887 1744 1921
rect 1686 1872 1744 1887
rect 1844 2057 1902 2072
rect 1844 2023 1856 2057
rect 1890 2023 1902 2057
rect 1844 1989 1902 2023
rect 1844 1955 1856 1989
rect 1890 1955 1902 1989
rect 1844 1921 1902 1955
rect 1844 1887 1856 1921
rect 1890 1887 1902 1921
rect 1844 1872 1902 1887
rect 2018 2057 2076 2072
rect 2018 2023 2030 2057
rect 2064 2023 2076 2057
rect 2018 1989 2076 2023
rect 2018 1955 2030 1989
rect 2064 1955 2076 1989
rect 2018 1921 2076 1955
rect 2018 1887 2030 1921
rect 2064 1887 2076 1921
rect 2018 1872 2076 1887
rect 2176 2057 2234 2072
rect 2176 2023 2188 2057
rect 2222 2023 2234 2057
rect 2176 1989 2234 2023
rect 2176 1955 2188 1989
rect 2222 1955 2234 1989
rect 2176 1921 2234 1955
rect 2176 1887 2188 1921
rect 2222 1887 2234 1921
rect 2176 1872 2234 1887
rect 2360 2057 2418 2072
rect 2360 2023 2372 2057
rect 2406 2023 2418 2057
rect 2360 1989 2418 2023
rect 2360 1955 2372 1989
rect 2406 1955 2418 1989
rect 2360 1921 2418 1955
rect 2360 1887 2372 1921
rect 2406 1887 2418 1921
rect 2360 1872 2418 1887
rect 2518 2057 2576 2072
rect 2518 2023 2530 2057
rect 2564 2023 2576 2057
rect 2518 1989 2576 2023
rect 2518 1955 2530 1989
rect 2564 1955 2576 1989
rect 2518 1921 2576 1955
rect 2518 1887 2530 1921
rect 2564 1887 2576 1921
rect 2518 1872 2576 1887
rect 2764 2057 2822 2072
rect 2764 2023 2776 2057
rect 2810 2023 2822 2057
rect 2764 1989 2822 2023
rect 2764 1955 2776 1989
rect 2810 1955 2822 1989
rect 2764 1921 2822 1955
rect 2764 1887 2776 1921
rect 2810 1887 2822 1921
rect 2764 1872 2822 1887
rect 2922 2057 2980 2072
rect 2922 2023 2934 2057
rect 2968 2023 2980 2057
rect 2922 1989 2980 2023
rect 2922 1955 2934 1989
rect 2968 1955 2980 1989
rect 2922 1921 2980 1955
rect 2922 1887 2934 1921
rect 2968 1887 2980 1921
rect 2922 1872 2980 1887
rect 3108 2057 3166 2072
rect 3108 2023 3120 2057
rect 3154 2023 3166 2057
rect 3108 1989 3166 2023
rect 3108 1955 3120 1989
rect 3154 1955 3166 1989
rect 3108 1921 3166 1955
rect 3108 1887 3120 1921
rect 3154 1887 3166 1921
rect 3108 1872 3166 1887
rect 3266 2057 3324 2072
rect 3266 2023 3278 2057
rect 3312 2023 3324 2057
rect 3266 1989 3324 2023
rect 3266 1955 3278 1989
rect 3312 1955 3324 1989
rect 3266 1921 3324 1955
rect 3266 1887 3278 1921
rect 3312 1887 3324 1921
rect 3266 1872 3324 1887
rect 3730 2067 3788 2082
rect 3730 2033 3742 2067
rect 3776 2033 3788 2067
rect 3730 1999 3788 2033
rect 3730 1965 3742 1999
rect 3776 1965 3788 1999
rect 3730 1931 3788 1965
rect 3730 1897 3742 1931
rect 3776 1897 3788 1931
rect 3730 1882 3788 1897
rect 3888 2067 3946 2082
rect 3888 2033 3900 2067
rect 3934 2033 3946 2067
rect 3888 1999 3946 2033
rect 3888 1965 3900 1999
rect 3934 1965 3946 1999
rect 3888 1931 3946 1965
rect 3888 1897 3900 1931
rect 3934 1897 3946 1931
rect 3888 1882 3946 1897
rect 4038 2067 4096 2082
rect 4038 2033 4050 2067
rect 4084 2033 4096 2067
rect 4038 1999 4096 2033
rect 4038 1965 4050 1999
rect 4084 1965 4096 1999
rect 4038 1931 4096 1965
rect 4038 1897 4050 1931
rect 4084 1897 4096 1931
rect 4038 1882 4096 1897
rect 4196 2067 4254 2082
rect 4196 2033 4208 2067
rect 4242 2033 4254 2067
rect 4196 1999 4254 2033
rect 4196 1965 4208 1999
rect 4242 1965 4254 1999
rect 4196 1931 4254 1965
rect 4196 1897 4208 1931
rect 4242 1897 4254 1931
rect 4196 1882 4254 1897
rect 4390 2067 4448 2082
rect 4390 2033 4402 2067
rect 4436 2033 4448 2067
rect 4390 1999 4448 2033
rect 4390 1965 4402 1999
rect 4436 1965 4448 1999
rect 4390 1931 4448 1965
rect 4390 1897 4402 1931
rect 4436 1897 4448 1931
rect 4390 1882 4448 1897
rect 4548 2067 4606 2082
rect 4548 2033 4560 2067
rect 4594 2033 4606 2067
rect 4548 1999 4606 2033
rect 4548 1965 4560 1999
rect 4594 1965 4606 1999
rect 4548 1931 4606 1965
rect 4548 1897 4560 1931
rect 4594 1897 4606 1931
rect 4548 1882 4606 1897
rect 4698 2067 4756 2082
rect 4698 2033 4710 2067
rect 4744 2033 4756 2067
rect 4698 1999 4756 2033
rect 4698 1965 4710 1999
rect 4744 1965 4756 1999
rect 4698 1931 4756 1965
rect 4698 1897 4710 1931
rect 4744 1897 4756 1931
rect 4698 1882 4756 1897
rect 4856 2067 4914 2082
rect 4856 2033 4868 2067
rect 4902 2033 4914 2067
rect 4856 1999 4914 2033
rect 4856 1965 4868 1999
rect 4902 1965 4914 1999
rect 4856 1931 4914 1965
rect 4856 1897 4868 1931
rect 4902 1897 4914 1931
rect 4856 1882 4914 1897
rect 5688 2068 5746 2082
rect 5688 2034 5700 2068
rect 5734 2034 5746 2068
rect 5688 2000 5746 2034
rect 5688 1966 5700 2000
rect 5734 1966 5746 2000
rect 5688 1932 5746 1966
rect 5688 1898 5700 1932
rect 5734 1898 5746 1932
rect 5688 1882 5746 1898
rect 5846 2068 5904 2082
rect 5846 2034 5858 2068
rect 5892 2034 5904 2068
rect 5846 2000 5904 2034
rect 5846 1966 5858 2000
rect 5892 1966 5904 2000
rect 5846 1932 5904 1966
rect 5846 1898 5858 1932
rect 5892 1898 5904 1932
rect 5846 1882 5904 1898
rect 5996 2068 6054 2082
rect 5996 2034 6008 2068
rect 6042 2034 6054 2068
rect 5996 2000 6054 2034
rect 5996 1966 6008 2000
rect 6042 1966 6054 2000
rect 5996 1932 6054 1966
rect 5996 1898 6008 1932
rect 6042 1898 6054 1932
rect 5996 1882 6054 1898
rect 6154 2068 6212 2082
rect 6154 2034 6166 2068
rect 6200 2034 6212 2068
rect 6154 2000 6212 2034
rect 6154 1966 6166 2000
rect 6200 1966 6212 2000
rect 6154 1932 6212 1966
rect 6154 1898 6166 1932
rect 6200 1898 6212 1932
rect 6154 1882 6212 1898
rect 6348 2068 6406 2082
rect 6348 2034 6360 2068
rect 6394 2034 6406 2068
rect 6348 2000 6406 2034
rect 6348 1966 6360 2000
rect 6394 1966 6406 2000
rect 6348 1932 6406 1966
rect 6348 1898 6360 1932
rect 6394 1898 6406 1932
rect 6348 1882 6406 1898
rect 6506 2068 6564 2082
rect 6506 2034 6518 2068
rect 6552 2034 6564 2068
rect 6506 2000 6564 2034
rect 6506 1966 6518 2000
rect 6552 1966 6564 2000
rect 6506 1932 6564 1966
rect 6506 1898 6518 1932
rect 6552 1898 6564 1932
rect 6506 1882 6564 1898
rect 6656 2068 6714 2082
rect 6656 2034 6668 2068
rect 6702 2034 6714 2068
rect 6656 2000 6714 2034
rect 6656 1966 6668 2000
rect 6702 1966 6714 2000
rect 6656 1932 6714 1966
rect 6656 1898 6668 1932
rect 6702 1898 6714 1932
rect 6656 1882 6714 1898
rect 6814 2068 6872 2082
rect 6814 2034 6826 2068
rect 6860 2034 6872 2068
rect 6814 2000 6872 2034
rect 6814 1966 6826 2000
rect 6860 1966 6872 2000
rect 6814 1932 6872 1966
rect 6814 1898 6826 1932
rect 6860 1898 6872 1932
rect 6814 1882 6872 1898
rect 1398 829 1456 844
rect 1398 795 1410 829
rect 1444 795 1456 829
rect 1398 761 1456 795
rect 1398 727 1410 761
rect 1444 727 1456 761
rect 1398 693 1456 727
rect 1398 659 1410 693
rect 1444 659 1456 693
rect 1398 644 1456 659
rect 1556 829 1614 844
rect 1556 795 1568 829
rect 1602 795 1614 829
rect 1556 761 1614 795
rect 1556 727 1568 761
rect 1602 727 1614 761
rect 1556 693 1614 727
rect 1556 659 1568 693
rect 1602 659 1614 693
rect 1556 644 1614 659
rect 1686 829 1744 844
rect 1686 795 1698 829
rect 1732 795 1744 829
rect 1686 761 1744 795
rect 1686 727 1698 761
rect 1732 727 1744 761
rect 1686 693 1744 727
rect 1686 659 1698 693
rect 1732 659 1744 693
rect 1686 644 1744 659
rect 1844 829 1902 844
rect 1844 795 1856 829
rect 1890 795 1902 829
rect 1844 761 1902 795
rect 1844 727 1856 761
rect 1890 727 1902 761
rect 1844 693 1902 727
rect 1844 659 1856 693
rect 1890 659 1902 693
rect 1844 644 1902 659
rect 2018 829 2076 844
rect 2018 795 2030 829
rect 2064 795 2076 829
rect 2018 761 2076 795
rect 2018 727 2030 761
rect 2064 727 2076 761
rect 2018 693 2076 727
rect 2018 659 2030 693
rect 2064 659 2076 693
rect 2018 644 2076 659
rect 2176 829 2234 844
rect 2176 795 2188 829
rect 2222 795 2234 829
rect 2176 761 2234 795
rect 2176 727 2188 761
rect 2222 727 2234 761
rect 2176 693 2234 727
rect 2176 659 2188 693
rect 2222 659 2234 693
rect 2176 644 2234 659
rect 2360 829 2418 844
rect 2360 795 2372 829
rect 2406 795 2418 829
rect 2360 761 2418 795
rect 2360 727 2372 761
rect 2406 727 2418 761
rect 2360 693 2418 727
rect 2360 659 2372 693
rect 2406 659 2418 693
rect 2360 644 2418 659
rect 2518 829 2576 844
rect 2518 795 2530 829
rect 2564 795 2576 829
rect 2518 761 2576 795
rect 2518 727 2530 761
rect 2564 727 2576 761
rect 2518 693 2576 727
rect 2518 659 2530 693
rect 2564 659 2576 693
rect 2518 644 2576 659
rect 2764 829 2822 844
rect 2764 795 2776 829
rect 2810 795 2822 829
rect 2764 761 2822 795
rect 2764 727 2776 761
rect 2810 727 2822 761
rect 2764 693 2822 727
rect 2764 659 2776 693
rect 2810 659 2822 693
rect 2764 644 2822 659
rect 2922 829 2980 844
rect 2922 795 2934 829
rect 2968 795 2980 829
rect 2922 761 2980 795
rect 2922 727 2934 761
rect 2968 727 2980 761
rect 2922 693 2980 727
rect 2922 659 2934 693
rect 2968 659 2980 693
rect 2922 644 2980 659
rect 3108 829 3166 844
rect 3108 795 3120 829
rect 3154 795 3166 829
rect 3108 761 3166 795
rect 3108 727 3120 761
rect 3154 727 3166 761
rect 3108 693 3166 727
rect 3108 659 3120 693
rect 3154 659 3166 693
rect 3108 644 3166 659
rect 3266 829 3324 844
rect 3266 795 3278 829
rect 3312 795 3324 829
rect 3266 761 3324 795
rect 3266 727 3278 761
rect 3312 727 3324 761
rect 3266 693 3324 727
rect 3266 659 3278 693
rect 3312 659 3324 693
rect 3266 644 3324 659
rect 3730 839 3788 854
rect 3730 805 3742 839
rect 3776 805 3788 839
rect 3730 771 3788 805
rect 3730 737 3742 771
rect 3776 737 3788 771
rect 3730 703 3788 737
rect 3730 669 3742 703
rect 3776 669 3788 703
rect 3730 654 3788 669
rect 3888 839 3946 854
rect 3888 805 3900 839
rect 3934 805 3946 839
rect 3888 771 3946 805
rect 3888 737 3900 771
rect 3934 737 3946 771
rect 3888 703 3946 737
rect 3888 669 3900 703
rect 3934 669 3946 703
rect 3888 654 3946 669
rect 4038 839 4096 854
rect 4038 805 4050 839
rect 4084 805 4096 839
rect 4038 771 4096 805
rect 4038 737 4050 771
rect 4084 737 4096 771
rect 4038 703 4096 737
rect 4038 669 4050 703
rect 4084 669 4096 703
rect 4038 654 4096 669
rect 4196 839 4254 854
rect 4196 805 4208 839
rect 4242 805 4254 839
rect 4196 771 4254 805
rect 4196 737 4208 771
rect 4242 737 4254 771
rect 4196 703 4254 737
rect 4196 669 4208 703
rect 4242 669 4254 703
rect 4196 654 4254 669
rect 4390 839 4448 854
rect 4390 805 4402 839
rect 4436 805 4448 839
rect 4390 771 4448 805
rect 4390 737 4402 771
rect 4436 737 4448 771
rect 4390 703 4448 737
rect 4390 669 4402 703
rect 4436 669 4448 703
rect 4390 654 4448 669
rect 4548 839 4606 854
rect 4548 805 4560 839
rect 4594 805 4606 839
rect 4548 771 4606 805
rect 4548 737 4560 771
rect 4594 737 4606 771
rect 4548 703 4606 737
rect 4548 669 4560 703
rect 4594 669 4606 703
rect 4548 654 4606 669
rect 4698 839 4756 854
rect 4698 805 4710 839
rect 4744 805 4756 839
rect 4698 771 4756 805
rect 4698 737 4710 771
rect 4744 737 4756 771
rect 4698 703 4756 737
rect 4698 669 4710 703
rect 4744 669 4756 703
rect 4698 654 4756 669
rect 4856 839 4914 854
rect 4856 805 4868 839
rect 4902 805 4914 839
rect 4856 771 4914 805
rect 4856 737 4868 771
rect 4902 737 4914 771
rect 4856 703 4914 737
rect 4856 669 4868 703
rect 4902 669 4914 703
rect 4856 654 4914 669
<< mvndiffc >>
rect 569 19314 603 19348
rect 569 18746 603 18780
rect 715 19314 749 19348
rect 715 18746 749 18780
rect 859 19320 893 19354
rect 859 18752 893 18786
rect 1013 19320 1047 19354
rect 1410 18859 1444 18893
rect 1568 18859 1602 18893
rect 1698 18859 1732 18893
rect 1856 18859 1890 18893
rect 2030 18859 2064 18893
rect 2188 18859 2222 18893
rect 2372 18859 2406 18893
rect 2530 18859 2564 18893
rect 2776 18859 2810 18893
rect 2934 18859 2968 18893
rect 3120 18859 3154 18893
rect 3278 18859 3312 18893
rect 3742 18869 3776 18903
rect 3900 18869 3934 18903
rect 4050 18869 4084 18903
rect 4208 18869 4242 18903
rect 4402 18871 4436 18905
rect 4560 18871 4594 18905
rect 4710 18871 4744 18905
rect 4868 18871 4902 18905
rect 5700 18870 5734 18904
rect 5858 18870 5892 18904
rect 6008 18870 6042 18904
rect 6166 18870 6200 18904
rect 6360 18872 6394 18906
rect 6518 18872 6552 18906
rect 6668 18872 6702 18906
rect 6826 18872 6860 18906
rect 1013 18752 1047 18786
rect 569 18086 603 18120
rect 569 17518 603 17552
rect 715 18086 749 18120
rect 715 17518 749 17552
rect 859 18092 893 18126
rect 859 17524 893 17558
rect 1013 18092 1047 18126
rect 1410 17631 1444 17665
rect 1568 17631 1602 17665
rect 1698 17631 1732 17665
rect 1856 17631 1890 17665
rect 2030 17631 2064 17665
rect 2188 17631 2222 17665
rect 2372 17631 2406 17665
rect 2530 17631 2564 17665
rect 2776 17631 2810 17665
rect 2934 17631 2968 17665
rect 3120 17631 3154 17665
rect 3278 17631 3312 17665
rect 3742 17641 3776 17675
rect 3900 17641 3934 17675
rect 4050 17641 4084 17675
rect 4208 17641 4242 17675
rect 4402 17643 4436 17677
rect 4560 17643 4594 17677
rect 4710 17643 4744 17677
rect 4868 17643 4902 17677
rect 5700 17642 5734 17676
rect 5858 17642 5892 17676
rect 6008 17642 6042 17676
rect 6166 17642 6200 17676
rect 6360 17644 6394 17678
rect 6518 17644 6552 17678
rect 6668 17644 6702 17678
rect 6826 17644 6860 17678
rect 1013 17524 1047 17558
rect 569 16858 603 16892
rect 569 16290 603 16324
rect 715 16858 749 16892
rect 715 16290 749 16324
rect 859 16864 893 16898
rect 859 16296 893 16330
rect 1013 16864 1047 16898
rect 1410 16403 1444 16437
rect 1568 16403 1602 16437
rect 1698 16403 1732 16437
rect 1856 16403 1890 16437
rect 2030 16403 2064 16437
rect 2188 16403 2222 16437
rect 2372 16403 2406 16437
rect 2530 16403 2564 16437
rect 2776 16403 2810 16437
rect 2934 16403 2968 16437
rect 3120 16403 3154 16437
rect 3278 16403 3312 16437
rect 3742 16413 3776 16447
rect 3900 16413 3934 16447
rect 4050 16413 4084 16447
rect 4208 16413 4242 16447
rect 4402 16415 4436 16449
rect 4560 16415 4594 16449
rect 4710 16415 4744 16449
rect 4868 16415 4902 16449
rect 5700 16414 5734 16448
rect 5858 16414 5892 16448
rect 6008 16414 6042 16448
rect 6166 16414 6200 16448
rect 6360 16416 6394 16450
rect 6518 16416 6552 16450
rect 6668 16416 6702 16450
rect 6826 16416 6860 16450
rect 1013 16296 1047 16330
rect 569 15630 603 15664
rect 569 15062 603 15096
rect 715 15630 749 15664
rect 715 15062 749 15096
rect 859 15636 893 15670
rect 859 15068 893 15102
rect 1013 15636 1047 15670
rect 1410 15175 1444 15209
rect 1568 15175 1602 15209
rect 1698 15175 1732 15209
rect 1856 15175 1890 15209
rect 2030 15175 2064 15209
rect 2188 15175 2222 15209
rect 2372 15175 2406 15209
rect 2530 15175 2564 15209
rect 2776 15175 2810 15209
rect 2934 15175 2968 15209
rect 3120 15175 3154 15209
rect 3278 15175 3312 15209
rect 3742 15185 3776 15219
rect 3900 15185 3934 15219
rect 4050 15185 4084 15219
rect 4208 15185 4242 15219
rect 4402 15187 4436 15221
rect 4560 15187 4594 15221
rect 4710 15187 4744 15221
rect 4868 15187 4902 15221
rect 5700 15186 5734 15220
rect 5858 15186 5892 15220
rect 6008 15186 6042 15220
rect 6166 15186 6200 15220
rect 6360 15188 6394 15222
rect 6518 15188 6552 15222
rect 6668 15188 6702 15222
rect 6826 15188 6860 15222
rect 1013 15068 1047 15102
rect 569 14402 603 14436
rect 569 13834 603 13868
rect 715 14402 749 14436
rect 715 13834 749 13868
rect 859 14408 893 14442
rect 859 13840 893 13874
rect 1013 14408 1047 14442
rect 1410 13947 1444 13981
rect 1568 13947 1602 13981
rect 1698 13947 1732 13981
rect 1856 13947 1890 13981
rect 2030 13947 2064 13981
rect 2188 13947 2222 13981
rect 2372 13947 2406 13981
rect 2530 13947 2564 13981
rect 2776 13947 2810 13981
rect 2934 13947 2968 13981
rect 3120 13947 3154 13981
rect 3278 13947 3312 13981
rect 3742 13957 3776 13991
rect 3900 13957 3934 13991
rect 4050 13957 4084 13991
rect 4208 13957 4242 13991
rect 4402 13959 4436 13993
rect 4560 13959 4594 13993
rect 4710 13959 4744 13993
rect 4868 13959 4902 13993
rect 5700 13958 5734 13992
rect 5858 13958 5892 13992
rect 6008 13958 6042 13992
rect 6166 13958 6200 13992
rect 6360 13960 6394 13994
rect 6518 13960 6552 13994
rect 6668 13960 6702 13994
rect 6826 13960 6860 13994
rect 1013 13840 1047 13874
rect 569 13174 603 13208
rect 569 12606 603 12640
rect 715 13174 749 13208
rect 715 12606 749 12640
rect 859 13180 893 13214
rect 859 12612 893 12646
rect 1013 13180 1047 13214
rect 1410 12719 1444 12753
rect 1568 12719 1602 12753
rect 1698 12719 1732 12753
rect 1856 12719 1890 12753
rect 2030 12719 2064 12753
rect 2188 12719 2222 12753
rect 2372 12719 2406 12753
rect 2530 12719 2564 12753
rect 2776 12719 2810 12753
rect 2934 12719 2968 12753
rect 3120 12719 3154 12753
rect 3278 12719 3312 12753
rect 3742 12729 3776 12763
rect 3900 12729 3934 12763
rect 4050 12729 4084 12763
rect 4208 12729 4242 12763
rect 4402 12731 4436 12765
rect 4560 12731 4594 12765
rect 4710 12731 4744 12765
rect 4868 12731 4902 12765
rect 5700 12730 5734 12764
rect 5858 12730 5892 12764
rect 6008 12730 6042 12764
rect 6166 12730 6200 12764
rect 6360 12732 6394 12766
rect 6518 12732 6552 12766
rect 6668 12732 6702 12766
rect 6826 12732 6860 12766
rect 1013 12612 1047 12646
rect 569 11946 603 11980
rect 569 11378 603 11412
rect 715 11946 749 11980
rect 715 11378 749 11412
rect 859 11952 893 11986
rect 859 11384 893 11418
rect 1013 11952 1047 11986
rect 1410 11491 1444 11525
rect 1568 11491 1602 11525
rect 1698 11491 1732 11525
rect 1856 11491 1890 11525
rect 2030 11491 2064 11525
rect 2188 11491 2222 11525
rect 2372 11491 2406 11525
rect 2530 11491 2564 11525
rect 2776 11491 2810 11525
rect 2934 11491 2968 11525
rect 3120 11491 3154 11525
rect 3278 11491 3312 11525
rect 3742 11501 3776 11535
rect 3900 11501 3934 11535
rect 4050 11501 4084 11535
rect 4208 11501 4242 11535
rect 4402 11503 4436 11537
rect 4560 11503 4594 11537
rect 4710 11503 4744 11537
rect 4868 11503 4902 11537
rect 5700 11502 5734 11536
rect 5858 11502 5892 11536
rect 6008 11502 6042 11536
rect 6166 11502 6200 11536
rect 6360 11504 6394 11538
rect 6518 11504 6552 11538
rect 6668 11504 6702 11538
rect 6826 11504 6860 11538
rect 1013 11384 1047 11418
rect 569 10718 603 10752
rect 569 10150 603 10184
rect 715 10718 749 10752
rect 715 10150 749 10184
rect 859 10724 893 10758
rect 859 10156 893 10190
rect 1013 10724 1047 10758
rect 1410 10263 1444 10297
rect 1568 10263 1602 10297
rect 1698 10263 1732 10297
rect 1856 10263 1890 10297
rect 2030 10263 2064 10297
rect 2188 10263 2222 10297
rect 2372 10263 2406 10297
rect 2530 10263 2564 10297
rect 2776 10263 2810 10297
rect 2934 10263 2968 10297
rect 3120 10263 3154 10297
rect 3278 10263 3312 10297
rect 3742 10273 3776 10307
rect 3900 10273 3934 10307
rect 4050 10273 4084 10307
rect 4208 10273 4242 10307
rect 4402 10275 4436 10309
rect 4560 10275 4594 10309
rect 4710 10275 4744 10309
rect 4868 10275 4902 10309
rect 5700 10274 5734 10308
rect 5858 10274 5892 10308
rect 6008 10274 6042 10308
rect 6166 10274 6200 10308
rect 6360 10276 6394 10310
rect 6518 10276 6552 10310
rect 6668 10276 6702 10310
rect 6826 10276 6860 10310
rect 1013 10156 1047 10190
rect 569 9490 603 9524
rect 569 8922 603 8956
rect 715 9490 749 9524
rect 715 8922 749 8956
rect 859 9496 893 9530
rect 859 8928 893 8962
rect 1013 9496 1047 9530
rect 1410 9035 1444 9069
rect 1568 9035 1602 9069
rect 1698 9035 1732 9069
rect 1856 9035 1890 9069
rect 2030 9035 2064 9069
rect 2188 9035 2222 9069
rect 2372 9035 2406 9069
rect 2530 9035 2564 9069
rect 2776 9035 2810 9069
rect 2934 9035 2968 9069
rect 3120 9035 3154 9069
rect 3278 9035 3312 9069
rect 3742 9045 3776 9079
rect 3900 9045 3934 9079
rect 4050 9045 4084 9079
rect 4208 9045 4242 9079
rect 4402 9047 4436 9081
rect 4560 9047 4594 9081
rect 4710 9047 4744 9081
rect 4868 9047 4902 9081
rect 5700 9046 5734 9080
rect 5858 9046 5892 9080
rect 6008 9046 6042 9080
rect 6166 9046 6200 9080
rect 6360 9048 6394 9082
rect 6518 9048 6552 9082
rect 6668 9048 6702 9082
rect 6826 9048 6860 9082
rect 1013 8928 1047 8962
rect 569 8262 603 8296
rect 569 7694 603 7728
rect 715 8262 749 8296
rect 715 7694 749 7728
rect 859 8268 893 8302
rect 859 7700 893 7734
rect 1013 8268 1047 8302
rect 1410 7807 1444 7841
rect 1568 7807 1602 7841
rect 1698 7807 1732 7841
rect 1856 7807 1890 7841
rect 2030 7807 2064 7841
rect 2188 7807 2222 7841
rect 2372 7807 2406 7841
rect 2530 7807 2564 7841
rect 2776 7807 2810 7841
rect 2934 7807 2968 7841
rect 3120 7807 3154 7841
rect 3278 7807 3312 7841
rect 3742 7817 3776 7851
rect 3900 7817 3934 7851
rect 4050 7817 4084 7851
rect 4208 7817 4242 7851
rect 4402 7819 4436 7853
rect 4560 7819 4594 7853
rect 4710 7819 4744 7853
rect 4868 7819 4902 7853
rect 5700 7818 5734 7852
rect 5858 7818 5892 7852
rect 6008 7818 6042 7852
rect 6166 7818 6200 7852
rect 6360 7820 6394 7854
rect 6518 7820 6552 7854
rect 6668 7820 6702 7854
rect 6826 7820 6860 7854
rect 1013 7700 1047 7734
rect 569 7034 603 7068
rect 569 6466 603 6500
rect 715 7034 749 7068
rect 715 6466 749 6500
rect 859 7040 893 7074
rect 859 6472 893 6506
rect 1013 7040 1047 7074
rect 1410 6579 1444 6613
rect 1568 6579 1602 6613
rect 1698 6579 1732 6613
rect 1856 6579 1890 6613
rect 2030 6579 2064 6613
rect 2188 6579 2222 6613
rect 2372 6579 2406 6613
rect 2530 6579 2564 6613
rect 2776 6579 2810 6613
rect 2934 6579 2968 6613
rect 3120 6579 3154 6613
rect 3278 6579 3312 6613
rect 3742 6589 3776 6623
rect 3900 6589 3934 6623
rect 4050 6589 4084 6623
rect 4208 6589 4242 6623
rect 4402 6591 4436 6625
rect 4560 6591 4594 6625
rect 4710 6591 4744 6625
rect 4868 6591 4902 6625
rect 5700 6590 5734 6624
rect 5858 6590 5892 6624
rect 6008 6590 6042 6624
rect 6166 6590 6200 6624
rect 6360 6592 6394 6626
rect 6518 6592 6552 6626
rect 6668 6592 6702 6626
rect 6826 6592 6860 6626
rect 1013 6472 1047 6506
rect 569 5806 603 5840
rect 569 5238 603 5272
rect 715 5806 749 5840
rect 715 5238 749 5272
rect 859 5812 893 5846
rect 859 5244 893 5278
rect 1013 5812 1047 5846
rect 1410 5351 1444 5385
rect 1568 5351 1602 5385
rect 1698 5351 1732 5385
rect 1856 5351 1890 5385
rect 2030 5351 2064 5385
rect 2188 5351 2222 5385
rect 2372 5351 2406 5385
rect 2530 5351 2564 5385
rect 2776 5351 2810 5385
rect 2934 5351 2968 5385
rect 3120 5351 3154 5385
rect 3278 5351 3312 5385
rect 3742 5361 3776 5395
rect 3900 5361 3934 5395
rect 4050 5361 4084 5395
rect 4208 5361 4242 5395
rect 4402 5363 4436 5397
rect 4560 5363 4594 5397
rect 4710 5363 4744 5397
rect 4868 5363 4902 5397
rect 5700 5362 5734 5396
rect 5858 5362 5892 5396
rect 6008 5362 6042 5396
rect 6166 5362 6200 5396
rect 6360 5364 6394 5398
rect 6518 5364 6552 5398
rect 6668 5364 6702 5398
rect 6826 5364 6860 5398
rect 1013 5244 1047 5278
rect 569 4578 603 4612
rect 569 4010 603 4044
rect 715 4578 749 4612
rect 715 4010 749 4044
rect 859 4584 893 4618
rect 859 4016 893 4050
rect 1013 4584 1047 4618
rect 1410 4123 1444 4157
rect 1568 4123 1602 4157
rect 1698 4123 1732 4157
rect 1856 4123 1890 4157
rect 2030 4123 2064 4157
rect 2188 4123 2222 4157
rect 2372 4123 2406 4157
rect 2530 4123 2564 4157
rect 2776 4123 2810 4157
rect 2934 4123 2968 4157
rect 3120 4123 3154 4157
rect 3278 4123 3312 4157
rect 3742 4133 3776 4167
rect 3900 4133 3934 4167
rect 4050 4133 4084 4167
rect 4208 4133 4242 4167
rect 4402 4135 4436 4169
rect 4560 4135 4594 4169
rect 4710 4135 4744 4169
rect 4868 4135 4902 4169
rect 5700 4134 5734 4168
rect 5858 4134 5892 4168
rect 6008 4134 6042 4168
rect 6166 4134 6200 4168
rect 6360 4136 6394 4170
rect 6518 4136 6552 4170
rect 6668 4136 6702 4170
rect 6826 4136 6860 4170
rect 1013 4016 1047 4050
rect 569 3350 603 3384
rect 569 2782 603 2816
rect 715 3350 749 3384
rect 715 2782 749 2816
rect 859 3356 893 3390
rect 859 2788 893 2822
rect 1013 3356 1047 3390
rect 1410 2895 1444 2929
rect 1568 2895 1602 2929
rect 1698 2895 1732 2929
rect 1856 2895 1890 2929
rect 2030 2895 2064 2929
rect 2188 2895 2222 2929
rect 2372 2895 2406 2929
rect 2530 2895 2564 2929
rect 2776 2895 2810 2929
rect 2934 2895 2968 2929
rect 3120 2895 3154 2929
rect 3278 2895 3312 2929
rect 3742 2905 3776 2939
rect 3900 2905 3934 2939
rect 4050 2905 4084 2939
rect 4208 2905 4242 2939
rect 4402 2907 4436 2941
rect 4560 2907 4594 2941
rect 4710 2907 4744 2941
rect 4868 2907 4902 2941
rect 5700 2906 5734 2940
rect 5858 2906 5892 2940
rect 6008 2906 6042 2940
rect 6166 2906 6200 2940
rect 6360 2908 6394 2942
rect 6518 2908 6552 2942
rect 6668 2908 6702 2942
rect 6826 2908 6860 2942
rect 1013 2788 1047 2822
rect 569 2122 603 2156
rect 569 1554 603 1588
rect 715 2122 749 2156
rect 715 1554 749 1588
rect 859 2128 893 2162
rect 859 1560 893 1594
rect 1013 2128 1047 2162
rect 1410 1667 1444 1701
rect 1568 1667 1602 1701
rect 1698 1667 1732 1701
rect 1856 1667 1890 1701
rect 2030 1667 2064 1701
rect 2188 1667 2222 1701
rect 2372 1667 2406 1701
rect 2530 1667 2564 1701
rect 2776 1667 2810 1701
rect 2934 1667 2968 1701
rect 3120 1667 3154 1701
rect 3278 1667 3312 1701
rect 3742 1677 3776 1711
rect 3900 1677 3934 1711
rect 4050 1677 4084 1711
rect 4208 1677 4242 1711
rect 4402 1679 4436 1713
rect 4560 1679 4594 1713
rect 4710 1679 4744 1713
rect 4868 1679 4902 1713
rect 5700 1678 5734 1712
rect 5858 1678 5892 1712
rect 6008 1678 6042 1712
rect 6166 1678 6200 1712
rect 6360 1680 6394 1714
rect 6518 1680 6552 1714
rect 6668 1680 6702 1714
rect 6826 1680 6860 1714
rect 1013 1560 1047 1594
rect 569 894 603 928
rect 569 326 603 360
rect 715 894 749 928
rect 715 326 749 360
rect 859 900 893 934
rect 859 332 893 366
rect 1013 900 1047 934
rect 1410 439 1444 473
rect 1568 439 1602 473
rect 1698 439 1732 473
rect 1856 439 1890 473
rect 2030 439 2064 473
rect 2188 439 2222 473
rect 2372 439 2406 473
rect 2530 439 2564 473
rect 2776 439 2810 473
rect 2934 439 2968 473
rect 3120 439 3154 473
rect 3278 439 3312 473
rect 3742 449 3776 483
rect 3900 449 3934 483
rect 4050 449 4084 483
rect 4208 449 4242 483
rect 4402 451 4436 485
rect 4560 451 4594 485
rect 4710 451 4744 485
rect 4868 451 4902 485
rect 1013 332 1047 366
<< mvpdiffc >>
rect 1410 19215 1444 19249
rect 1410 19147 1444 19181
rect 1410 19079 1444 19113
rect 1568 19215 1602 19249
rect 1568 19147 1602 19181
rect 1568 19079 1602 19113
rect 1698 19215 1732 19249
rect 1698 19147 1732 19181
rect 1698 19079 1732 19113
rect 1856 19215 1890 19249
rect 1856 19147 1890 19181
rect 1856 19079 1890 19113
rect 2030 19215 2064 19249
rect 2030 19147 2064 19181
rect 2030 19079 2064 19113
rect 2188 19215 2222 19249
rect 2188 19147 2222 19181
rect 2188 19079 2222 19113
rect 2372 19215 2406 19249
rect 2372 19147 2406 19181
rect 2372 19079 2406 19113
rect 2530 19215 2564 19249
rect 2530 19147 2564 19181
rect 2530 19079 2564 19113
rect 2776 19215 2810 19249
rect 2776 19147 2810 19181
rect 2776 19079 2810 19113
rect 2934 19215 2968 19249
rect 2934 19147 2968 19181
rect 2934 19079 2968 19113
rect 3120 19215 3154 19249
rect 3120 19147 3154 19181
rect 3120 19079 3154 19113
rect 3278 19215 3312 19249
rect 3278 19147 3312 19181
rect 3278 19079 3312 19113
rect 3742 19225 3776 19259
rect 3742 19157 3776 19191
rect 3742 19089 3776 19123
rect 3900 19225 3934 19259
rect 3900 19157 3934 19191
rect 3900 19089 3934 19123
rect 4050 19225 4084 19259
rect 4050 19157 4084 19191
rect 4050 19089 4084 19123
rect 4208 19225 4242 19259
rect 4208 19157 4242 19191
rect 4208 19089 4242 19123
rect 4402 19225 4436 19259
rect 4402 19157 4436 19191
rect 4402 19089 4436 19123
rect 4560 19225 4594 19259
rect 4560 19157 4594 19191
rect 4560 19089 4594 19123
rect 4710 19225 4744 19259
rect 4710 19157 4744 19191
rect 4710 19089 4744 19123
rect 4868 19225 4902 19259
rect 4868 19157 4902 19191
rect 4868 19089 4902 19123
rect 5700 19226 5734 19260
rect 5700 19158 5734 19192
rect 5700 19090 5734 19124
rect 5858 19226 5892 19260
rect 5858 19158 5892 19192
rect 5858 19090 5892 19124
rect 6008 19226 6042 19260
rect 6008 19158 6042 19192
rect 6008 19090 6042 19124
rect 6166 19226 6200 19260
rect 6166 19158 6200 19192
rect 6166 19090 6200 19124
rect 6360 19226 6394 19260
rect 6360 19158 6394 19192
rect 6360 19090 6394 19124
rect 6518 19226 6552 19260
rect 6518 19158 6552 19192
rect 6518 19090 6552 19124
rect 6668 19226 6702 19260
rect 6668 19158 6702 19192
rect 6668 19090 6702 19124
rect 6826 19226 6860 19260
rect 6826 19158 6860 19192
rect 6826 19090 6860 19124
rect 1410 17987 1444 18021
rect 1410 17919 1444 17953
rect 1410 17851 1444 17885
rect 1568 17987 1602 18021
rect 1568 17919 1602 17953
rect 1568 17851 1602 17885
rect 1698 17987 1732 18021
rect 1698 17919 1732 17953
rect 1698 17851 1732 17885
rect 1856 17987 1890 18021
rect 1856 17919 1890 17953
rect 1856 17851 1890 17885
rect 2030 17987 2064 18021
rect 2030 17919 2064 17953
rect 2030 17851 2064 17885
rect 2188 17987 2222 18021
rect 2188 17919 2222 17953
rect 2188 17851 2222 17885
rect 2372 17987 2406 18021
rect 2372 17919 2406 17953
rect 2372 17851 2406 17885
rect 2530 17987 2564 18021
rect 2530 17919 2564 17953
rect 2530 17851 2564 17885
rect 2776 17987 2810 18021
rect 2776 17919 2810 17953
rect 2776 17851 2810 17885
rect 2934 17987 2968 18021
rect 2934 17919 2968 17953
rect 2934 17851 2968 17885
rect 3120 17987 3154 18021
rect 3120 17919 3154 17953
rect 3120 17851 3154 17885
rect 3278 17987 3312 18021
rect 3278 17919 3312 17953
rect 3278 17851 3312 17885
rect 3742 17997 3776 18031
rect 3742 17929 3776 17963
rect 3742 17861 3776 17895
rect 3900 17997 3934 18031
rect 3900 17929 3934 17963
rect 3900 17861 3934 17895
rect 4050 17997 4084 18031
rect 4050 17929 4084 17963
rect 4050 17861 4084 17895
rect 4208 17997 4242 18031
rect 4208 17929 4242 17963
rect 4208 17861 4242 17895
rect 4402 17997 4436 18031
rect 4402 17929 4436 17963
rect 4402 17861 4436 17895
rect 4560 17997 4594 18031
rect 4560 17929 4594 17963
rect 4560 17861 4594 17895
rect 4710 17997 4744 18031
rect 4710 17929 4744 17963
rect 4710 17861 4744 17895
rect 4868 17997 4902 18031
rect 4868 17929 4902 17963
rect 4868 17861 4902 17895
rect 5700 17998 5734 18032
rect 5700 17930 5734 17964
rect 5700 17862 5734 17896
rect 5858 17998 5892 18032
rect 5858 17930 5892 17964
rect 5858 17862 5892 17896
rect 6008 17998 6042 18032
rect 6008 17930 6042 17964
rect 6008 17862 6042 17896
rect 6166 17998 6200 18032
rect 6166 17930 6200 17964
rect 6166 17862 6200 17896
rect 6360 17998 6394 18032
rect 6360 17930 6394 17964
rect 6360 17862 6394 17896
rect 6518 17998 6552 18032
rect 6518 17930 6552 17964
rect 6518 17862 6552 17896
rect 6668 17998 6702 18032
rect 6668 17930 6702 17964
rect 6668 17862 6702 17896
rect 6826 17998 6860 18032
rect 6826 17930 6860 17964
rect 6826 17862 6860 17896
rect 1410 16759 1444 16793
rect 1410 16691 1444 16725
rect 1410 16623 1444 16657
rect 1568 16759 1602 16793
rect 1568 16691 1602 16725
rect 1568 16623 1602 16657
rect 1698 16759 1732 16793
rect 1698 16691 1732 16725
rect 1698 16623 1732 16657
rect 1856 16759 1890 16793
rect 1856 16691 1890 16725
rect 1856 16623 1890 16657
rect 2030 16759 2064 16793
rect 2030 16691 2064 16725
rect 2030 16623 2064 16657
rect 2188 16759 2222 16793
rect 2188 16691 2222 16725
rect 2188 16623 2222 16657
rect 2372 16759 2406 16793
rect 2372 16691 2406 16725
rect 2372 16623 2406 16657
rect 2530 16759 2564 16793
rect 2530 16691 2564 16725
rect 2530 16623 2564 16657
rect 2776 16759 2810 16793
rect 2776 16691 2810 16725
rect 2776 16623 2810 16657
rect 2934 16759 2968 16793
rect 2934 16691 2968 16725
rect 2934 16623 2968 16657
rect 3120 16759 3154 16793
rect 3120 16691 3154 16725
rect 3120 16623 3154 16657
rect 3278 16759 3312 16793
rect 3278 16691 3312 16725
rect 3278 16623 3312 16657
rect 3742 16769 3776 16803
rect 3742 16701 3776 16735
rect 3742 16633 3776 16667
rect 3900 16769 3934 16803
rect 3900 16701 3934 16735
rect 3900 16633 3934 16667
rect 4050 16769 4084 16803
rect 4050 16701 4084 16735
rect 4050 16633 4084 16667
rect 4208 16769 4242 16803
rect 4208 16701 4242 16735
rect 4208 16633 4242 16667
rect 4402 16769 4436 16803
rect 4402 16701 4436 16735
rect 4402 16633 4436 16667
rect 4560 16769 4594 16803
rect 4560 16701 4594 16735
rect 4560 16633 4594 16667
rect 4710 16769 4744 16803
rect 4710 16701 4744 16735
rect 4710 16633 4744 16667
rect 4868 16769 4902 16803
rect 4868 16701 4902 16735
rect 4868 16633 4902 16667
rect 5700 16770 5734 16804
rect 5700 16702 5734 16736
rect 5700 16634 5734 16668
rect 5858 16770 5892 16804
rect 5858 16702 5892 16736
rect 5858 16634 5892 16668
rect 6008 16770 6042 16804
rect 6008 16702 6042 16736
rect 6008 16634 6042 16668
rect 6166 16770 6200 16804
rect 6166 16702 6200 16736
rect 6166 16634 6200 16668
rect 6360 16770 6394 16804
rect 6360 16702 6394 16736
rect 6360 16634 6394 16668
rect 6518 16770 6552 16804
rect 6518 16702 6552 16736
rect 6518 16634 6552 16668
rect 6668 16770 6702 16804
rect 6668 16702 6702 16736
rect 6668 16634 6702 16668
rect 6826 16770 6860 16804
rect 6826 16702 6860 16736
rect 6826 16634 6860 16668
rect 1410 15531 1444 15565
rect 1410 15463 1444 15497
rect 1410 15395 1444 15429
rect 1568 15531 1602 15565
rect 1568 15463 1602 15497
rect 1568 15395 1602 15429
rect 1698 15531 1732 15565
rect 1698 15463 1732 15497
rect 1698 15395 1732 15429
rect 1856 15531 1890 15565
rect 1856 15463 1890 15497
rect 1856 15395 1890 15429
rect 2030 15531 2064 15565
rect 2030 15463 2064 15497
rect 2030 15395 2064 15429
rect 2188 15531 2222 15565
rect 2188 15463 2222 15497
rect 2188 15395 2222 15429
rect 2372 15531 2406 15565
rect 2372 15463 2406 15497
rect 2372 15395 2406 15429
rect 2530 15531 2564 15565
rect 2530 15463 2564 15497
rect 2530 15395 2564 15429
rect 2776 15531 2810 15565
rect 2776 15463 2810 15497
rect 2776 15395 2810 15429
rect 2934 15531 2968 15565
rect 2934 15463 2968 15497
rect 2934 15395 2968 15429
rect 3120 15531 3154 15565
rect 3120 15463 3154 15497
rect 3120 15395 3154 15429
rect 3278 15531 3312 15565
rect 3278 15463 3312 15497
rect 3278 15395 3312 15429
rect 3742 15541 3776 15575
rect 3742 15473 3776 15507
rect 3742 15405 3776 15439
rect 3900 15541 3934 15575
rect 3900 15473 3934 15507
rect 3900 15405 3934 15439
rect 4050 15541 4084 15575
rect 4050 15473 4084 15507
rect 4050 15405 4084 15439
rect 4208 15541 4242 15575
rect 4208 15473 4242 15507
rect 4208 15405 4242 15439
rect 4402 15541 4436 15575
rect 4402 15473 4436 15507
rect 4402 15405 4436 15439
rect 4560 15541 4594 15575
rect 4560 15473 4594 15507
rect 4560 15405 4594 15439
rect 4710 15541 4744 15575
rect 4710 15473 4744 15507
rect 4710 15405 4744 15439
rect 4868 15541 4902 15575
rect 4868 15473 4902 15507
rect 4868 15405 4902 15439
rect 5700 15542 5734 15576
rect 5700 15474 5734 15508
rect 5700 15406 5734 15440
rect 5858 15542 5892 15576
rect 5858 15474 5892 15508
rect 5858 15406 5892 15440
rect 6008 15542 6042 15576
rect 6008 15474 6042 15508
rect 6008 15406 6042 15440
rect 6166 15542 6200 15576
rect 6166 15474 6200 15508
rect 6166 15406 6200 15440
rect 6360 15542 6394 15576
rect 6360 15474 6394 15508
rect 6360 15406 6394 15440
rect 6518 15542 6552 15576
rect 6518 15474 6552 15508
rect 6518 15406 6552 15440
rect 6668 15542 6702 15576
rect 6668 15474 6702 15508
rect 6668 15406 6702 15440
rect 6826 15542 6860 15576
rect 6826 15474 6860 15508
rect 6826 15406 6860 15440
rect 1410 14303 1444 14337
rect 1410 14235 1444 14269
rect 1410 14167 1444 14201
rect 1568 14303 1602 14337
rect 1568 14235 1602 14269
rect 1568 14167 1602 14201
rect 1698 14303 1732 14337
rect 1698 14235 1732 14269
rect 1698 14167 1732 14201
rect 1856 14303 1890 14337
rect 1856 14235 1890 14269
rect 1856 14167 1890 14201
rect 2030 14303 2064 14337
rect 2030 14235 2064 14269
rect 2030 14167 2064 14201
rect 2188 14303 2222 14337
rect 2188 14235 2222 14269
rect 2188 14167 2222 14201
rect 2372 14303 2406 14337
rect 2372 14235 2406 14269
rect 2372 14167 2406 14201
rect 2530 14303 2564 14337
rect 2530 14235 2564 14269
rect 2530 14167 2564 14201
rect 2776 14303 2810 14337
rect 2776 14235 2810 14269
rect 2776 14167 2810 14201
rect 2934 14303 2968 14337
rect 2934 14235 2968 14269
rect 2934 14167 2968 14201
rect 3120 14303 3154 14337
rect 3120 14235 3154 14269
rect 3120 14167 3154 14201
rect 3278 14303 3312 14337
rect 3278 14235 3312 14269
rect 3278 14167 3312 14201
rect 3742 14313 3776 14347
rect 3742 14245 3776 14279
rect 3742 14177 3776 14211
rect 3900 14313 3934 14347
rect 3900 14245 3934 14279
rect 3900 14177 3934 14211
rect 4050 14313 4084 14347
rect 4050 14245 4084 14279
rect 4050 14177 4084 14211
rect 4208 14313 4242 14347
rect 4208 14245 4242 14279
rect 4208 14177 4242 14211
rect 4402 14313 4436 14347
rect 4402 14245 4436 14279
rect 4402 14177 4436 14211
rect 4560 14313 4594 14347
rect 4560 14245 4594 14279
rect 4560 14177 4594 14211
rect 4710 14313 4744 14347
rect 4710 14245 4744 14279
rect 4710 14177 4744 14211
rect 4868 14313 4902 14347
rect 4868 14245 4902 14279
rect 4868 14177 4902 14211
rect 5700 14314 5734 14348
rect 5700 14246 5734 14280
rect 5700 14178 5734 14212
rect 5858 14314 5892 14348
rect 5858 14246 5892 14280
rect 5858 14178 5892 14212
rect 6008 14314 6042 14348
rect 6008 14246 6042 14280
rect 6008 14178 6042 14212
rect 6166 14314 6200 14348
rect 6166 14246 6200 14280
rect 6166 14178 6200 14212
rect 6360 14314 6394 14348
rect 6360 14246 6394 14280
rect 6360 14178 6394 14212
rect 6518 14314 6552 14348
rect 6518 14246 6552 14280
rect 6518 14178 6552 14212
rect 6668 14314 6702 14348
rect 6668 14246 6702 14280
rect 6668 14178 6702 14212
rect 6826 14314 6860 14348
rect 6826 14246 6860 14280
rect 6826 14178 6860 14212
rect 1410 13075 1444 13109
rect 1410 13007 1444 13041
rect 1410 12939 1444 12973
rect 1568 13075 1602 13109
rect 1568 13007 1602 13041
rect 1568 12939 1602 12973
rect 1698 13075 1732 13109
rect 1698 13007 1732 13041
rect 1698 12939 1732 12973
rect 1856 13075 1890 13109
rect 1856 13007 1890 13041
rect 1856 12939 1890 12973
rect 2030 13075 2064 13109
rect 2030 13007 2064 13041
rect 2030 12939 2064 12973
rect 2188 13075 2222 13109
rect 2188 13007 2222 13041
rect 2188 12939 2222 12973
rect 2372 13075 2406 13109
rect 2372 13007 2406 13041
rect 2372 12939 2406 12973
rect 2530 13075 2564 13109
rect 2530 13007 2564 13041
rect 2530 12939 2564 12973
rect 2776 13075 2810 13109
rect 2776 13007 2810 13041
rect 2776 12939 2810 12973
rect 2934 13075 2968 13109
rect 2934 13007 2968 13041
rect 2934 12939 2968 12973
rect 3120 13075 3154 13109
rect 3120 13007 3154 13041
rect 3120 12939 3154 12973
rect 3278 13075 3312 13109
rect 3278 13007 3312 13041
rect 3278 12939 3312 12973
rect 3742 13085 3776 13119
rect 3742 13017 3776 13051
rect 3742 12949 3776 12983
rect 3900 13085 3934 13119
rect 3900 13017 3934 13051
rect 3900 12949 3934 12983
rect 4050 13085 4084 13119
rect 4050 13017 4084 13051
rect 4050 12949 4084 12983
rect 4208 13085 4242 13119
rect 4208 13017 4242 13051
rect 4208 12949 4242 12983
rect 4402 13085 4436 13119
rect 4402 13017 4436 13051
rect 4402 12949 4436 12983
rect 4560 13085 4594 13119
rect 4560 13017 4594 13051
rect 4560 12949 4594 12983
rect 4710 13085 4744 13119
rect 4710 13017 4744 13051
rect 4710 12949 4744 12983
rect 4868 13085 4902 13119
rect 4868 13017 4902 13051
rect 4868 12949 4902 12983
rect 5700 13086 5734 13120
rect 5700 13018 5734 13052
rect 5700 12950 5734 12984
rect 5858 13086 5892 13120
rect 5858 13018 5892 13052
rect 5858 12950 5892 12984
rect 6008 13086 6042 13120
rect 6008 13018 6042 13052
rect 6008 12950 6042 12984
rect 6166 13086 6200 13120
rect 6166 13018 6200 13052
rect 6166 12950 6200 12984
rect 6360 13086 6394 13120
rect 6360 13018 6394 13052
rect 6360 12950 6394 12984
rect 6518 13086 6552 13120
rect 6518 13018 6552 13052
rect 6518 12950 6552 12984
rect 6668 13086 6702 13120
rect 6668 13018 6702 13052
rect 6668 12950 6702 12984
rect 6826 13086 6860 13120
rect 6826 13018 6860 13052
rect 6826 12950 6860 12984
rect 1410 11847 1444 11881
rect 1410 11779 1444 11813
rect 1410 11711 1444 11745
rect 1568 11847 1602 11881
rect 1568 11779 1602 11813
rect 1568 11711 1602 11745
rect 1698 11847 1732 11881
rect 1698 11779 1732 11813
rect 1698 11711 1732 11745
rect 1856 11847 1890 11881
rect 1856 11779 1890 11813
rect 1856 11711 1890 11745
rect 2030 11847 2064 11881
rect 2030 11779 2064 11813
rect 2030 11711 2064 11745
rect 2188 11847 2222 11881
rect 2188 11779 2222 11813
rect 2188 11711 2222 11745
rect 2372 11847 2406 11881
rect 2372 11779 2406 11813
rect 2372 11711 2406 11745
rect 2530 11847 2564 11881
rect 2530 11779 2564 11813
rect 2530 11711 2564 11745
rect 2776 11847 2810 11881
rect 2776 11779 2810 11813
rect 2776 11711 2810 11745
rect 2934 11847 2968 11881
rect 2934 11779 2968 11813
rect 2934 11711 2968 11745
rect 3120 11847 3154 11881
rect 3120 11779 3154 11813
rect 3120 11711 3154 11745
rect 3278 11847 3312 11881
rect 3278 11779 3312 11813
rect 3278 11711 3312 11745
rect 3742 11857 3776 11891
rect 3742 11789 3776 11823
rect 3742 11721 3776 11755
rect 3900 11857 3934 11891
rect 3900 11789 3934 11823
rect 3900 11721 3934 11755
rect 4050 11857 4084 11891
rect 4050 11789 4084 11823
rect 4050 11721 4084 11755
rect 4208 11857 4242 11891
rect 4208 11789 4242 11823
rect 4208 11721 4242 11755
rect 4402 11857 4436 11891
rect 4402 11789 4436 11823
rect 4402 11721 4436 11755
rect 4560 11857 4594 11891
rect 4560 11789 4594 11823
rect 4560 11721 4594 11755
rect 4710 11857 4744 11891
rect 4710 11789 4744 11823
rect 4710 11721 4744 11755
rect 4868 11857 4902 11891
rect 4868 11789 4902 11823
rect 4868 11721 4902 11755
rect 5700 11858 5734 11892
rect 5700 11790 5734 11824
rect 5700 11722 5734 11756
rect 5858 11858 5892 11892
rect 5858 11790 5892 11824
rect 5858 11722 5892 11756
rect 6008 11858 6042 11892
rect 6008 11790 6042 11824
rect 6008 11722 6042 11756
rect 6166 11858 6200 11892
rect 6166 11790 6200 11824
rect 6166 11722 6200 11756
rect 6360 11858 6394 11892
rect 6360 11790 6394 11824
rect 6360 11722 6394 11756
rect 6518 11858 6552 11892
rect 6518 11790 6552 11824
rect 6518 11722 6552 11756
rect 6668 11858 6702 11892
rect 6668 11790 6702 11824
rect 6668 11722 6702 11756
rect 6826 11858 6860 11892
rect 6826 11790 6860 11824
rect 6826 11722 6860 11756
rect 1410 10619 1444 10653
rect 1410 10551 1444 10585
rect 1410 10483 1444 10517
rect 1568 10619 1602 10653
rect 1568 10551 1602 10585
rect 1568 10483 1602 10517
rect 1698 10619 1732 10653
rect 1698 10551 1732 10585
rect 1698 10483 1732 10517
rect 1856 10619 1890 10653
rect 1856 10551 1890 10585
rect 1856 10483 1890 10517
rect 2030 10619 2064 10653
rect 2030 10551 2064 10585
rect 2030 10483 2064 10517
rect 2188 10619 2222 10653
rect 2188 10551 2222 10585
rect 2188 10483 2222 10517
rect 2372 10619 2406 10653
rect 2372 10551 2406 10585
rect 2372 10483 2406 10517
rect 2530 10619 2564 10653
rect 2530 10551 2564 10585
rect 2530 10483 2564 10517
rect 2776 10619 2810 10653
rect 2776 10551 2810 10585
rect 2776 10483 2810 10517
rect 2934 10619 2968 10653
rect 2934 10551 2968 10585
rect 2934 10483 2968 10517
rect 3120 10619 3154 10653
rect 3120 10551 3154 10585
rect 3120 10483 3154 10517
rect 3278 10619 3312 10653
rect 3278 10551 3312 10585
rect 3278 10483 3312 10517
rect 3742 10629 3776 10663
rect 3742 10561 3776 10595
rect 3742 10493 3776 10527
rect 3900 10629 3934 10663
rect 3900 10561 3934 10595
rect 3900 10493 3934 10527
rect 4050 10629 4084 10663
rect 4050 10561 4084 10595
rect 4050 10493 4084 10527
rect 4208 10629 4242 10663
rect 4208 10561 4242 10595
rect 4208 10493 4242 10527
rect 4402 10629 4436 10663
rect 4402 10561 4436 10595
rect 4402 10493 4436 10527
rect 4560 10629 4594 10663
rect 4560 10561 4594 10595
rect 4560 10493 4594 10527
rect 4710 10629 4744 10663
rect 4710 10561 4744 10595
rect 4710 10493 4744 10527
rect 4868 10629 4902 10663
rect 4868 10561 4902 10595
rect 4868 10493 4902 10527
rect 5700 10630 5734 10664
rect 5700 10562 5734 10596
rect 5700 10494 5734 10528
rect 5858 10630 5892 10664
rect 5858 10562 5892 10596
rect 5858 10494 5892 10528
rect 6008 10630 6042 10664
rect 6008 10562 6042 10596
rect 6008 10494 6042 10528
rect 6166 10630 6200 10664
rect 6166 10562 6200 10596
rect 6166 10494 6200 10528
rect 6360 10630 6394 10664
rect 6360 10562 6394 10596
rect 6360 10494 6394 10528
rect 6518 10630 6552 10664
rect 6518 10562 6552 10596
rect 6518 10494 6552 10528
rect 6668 10630 6702 10664
rect 6668 10562 6702 10596
rect 6668 10494 6702 10528
rect 6826 10630 6860 10664
rect 6826 10562 6860 10596
rect 6826 10494 6860 10528
rect 1410 9391 1444 9425
rect 1410 9323 1444 9357
rect 1410 9255 1444 9289
rect 1568 9391 1602 9425
rect 1568 9323 1602 9357
rect 1568 9255 1602 9289
rect 1698 9391 1732 9425
rect 1698 9323 1732 9357
rect 1698 9255 1732 9289
rect 1856 9391 1890 9425
rect 1856 9323 1890 9357
rect 1856 9255 1890 9289
rect 2030 9391 2064 9425
rect 2030 9323 2064 9357
rect 2030 9255 2064 9289
rect 2188 9391 2222 9425
rect 2188 9323 2222 9357
rect 2188 9255 2222 9289
rect 2372 9391 2406 9425
rect 2372 9323 2406 9357
rect 2372 9255 2406 9289
rect 2530 9391 2564 9425
rect 2530 9323 2564 9357
rect 2530 9255 2564 9289
rect 2776 9391 2810 9425
rect 2776 9323 2810 9357
rect 2776 9255 2810 9289
rect 2934 9391 2968 9425
rect 2934 9323 2968 9357
rect 2934 9255 2968 9289
rect 3120 9391 3154 9425
rect 3120 9323 3154 9357
rect 3120 9255 3154 9289
rect 3278 9391 3312 9425
rect 3278 9323 3312 9357
rect 3278 9255 3312 9289
rect 3742 9401 3776 9435
rect 3742 9333 3776 9367
rect 3742 9265 3776 9299
rect 3900 9401 3934 9435
rect 3900 9333 3934 9367
rect 3900 9265 3934 9299
rect 4050 9401 4084 9435
rect 4050 9333 4084 9367
rect 4050 9265 4084 9299
rect 4208 9401 4242 9435
rect 4208 9333 4242 9367
rect 4208 9265 4242 9299
rect 4402 9401 4436 9435
rect 4402 9333 4436 9367
rect 4402 9265 4436 9299
rect 4560 9401 4594 9435
rect 4560 9333 4594 9367
rect 4560 9265 4594 9299
rect 4710 9401 4744 9435
rect 4710 9333 4744 9367
rect 4710 9265 4744 9299
rect 4868 9401 4902 9435
rect 4868 9333 4902 9367
rect 4868 9265 4902 9299
rect 5700 9402 5734 9436
rect 5700 9334 5734 9368
rect 5700 9266 5734 9300
rect 5858 9402 5892 9436
rect 5858 9334 5892 9368
rect 5858 9266 5892 9300
rect 6008 9402 6042 9436
rect 6008 9334 6042 9368
rect 6008 9266 6042 9300
rect 6166 9402 6200 9436
rect 6166 9334 6200 9368
rect 6166 9266 6200 9300
rect 6360 9402 6394 9436
rect 6360 9334 6394 9368
rect 6360 9266 6394 9300
rect 6518 9402 6552 9436
rect 6518 9334 6552 9368
rect 6518 9266 6552 9300
rect 6668 9402 6702 9436
rect 6668 9334 6702 9368
rect 6668 9266 6702 9300
rect 6826 9402 6860 9436
rect 6826 9334 6860 9368
rect 6826 9266 6860 9300
rect 1410 8163 1444 8197
rect 1410 8095 1444 8129
rect 1410 8027 1444 8061
rect 1568 8163 1602 8197
rect 1568 8095 1602 8129
rect 1568 8027 1602 8061
rect 1698 8163 1732 8197
rect 1698 8095 1732 8129
rect 1698 8027 1732 8061
rect 1856 8163 1890 8197
rect 1856 8095 1890 8129
rect 1856 8027 1890 8061
rect 2030 8163 2064 8197
rect 2030 8095 2064 8129
rect 2030 8027 2064 8061
rect 2188 8163 2222 8197
rect 2188 8095 2222 8129
rect 2188 8027 2222 8061
rect 2372 8163 2406 8197
rect 2372 8095 2406 8129
rect 2372 8027 2406 8061
rect 2530 8163 2564 8197
rect 2530 8095 2564 8129
rect 2530 8027 2564 8061
rect 2776 8163 2810 8197
rect 2776 8095 2810 8129
rect 2776 8027 2810 8061
rect 2934 8163 2968 8197
rect 2934 8095 2968 8129
rect 2934 8027 2968 8061
rect 3120 8163 3154 8197
rect 3120 8095 3154 8129
rect 3120 8027 3154 8061
rect 3278 8163 3312 8197
rect 3278 8095 3312 8129
rect 3278 8027 3312 8061
rect 3742 8173 3776 8207
rect 3742 8105 3776 8139
rect 3742 8037 3776 8071
rect 3900 8173 3934 8207
rect 3900 8105 3934 8139
rect 3900 8037 3934 8071
rect 4050 8173 4084 8207
rect 4050 8105 4084 8139
rect 4050 8037 4084 8071
rect 4208 8173 4242 8207
rect 4208 8105 4242 8139
rect 4208 8037 4242 8071
rect 4402 8173 4436 8207
rect 4402 8105 4436 8139
rect 4402 8037 4436 8071
rect 4560 8173 4594 8207
rect 4560 8105 4594 8139
rect 4560 8037 4594 8071
rect 4710 8173 4744 8207
rect 4710 8105 4744 8139
rect 4710 8037 4744 8071
rect 4868 8173 4902 8207
rect 4868 8105 4902 8139
rect 4868 8037 4902 8071
rect 5700 8174 5734 8208
rect 5700 8106 5734 8140
rect 5700 8038 5734 8072
rect 5858 8174 5892 8208
rect 5858 8106 5892 8140
rect 5858 8038 5892 8072
rect 6008 8174 6042 8208
rect 6008 8106 6042 8140
rect 6008 8038 6042 8072
rect 6166 8174 6200 8208
rect 6166 8106 6200 8140
rect 6166 8038 6200 8072
rect 6360 8174 6394 8208
rect 6360 8106 6394 8140
rect 6360 8038 6394 8072
rect 6518 8174 6552 8208
rect 6518 8106 6552 8140
rect 6518 8038 6552 8072
rect 6668 8174 6702 8208
rect 6668 8106 6702 8140
rect 6668 8038 6702 8072
rect 6826 8174 6860 8208
rect 6826 8106 6860 8140
rect 6826 8038 6860 8072
rect 1410 6935 1444 6969
rect 1410 6867 1444 6901
rect 1410 6799 1444 6833
rect 1568 6935 1602 6969
rect 1568 6867 1602 6901
rect 1568 6799 1602 6833
rect 1698 6935 1732 6969
rect 1698 6867 1732 6901
rect 1698 6799 1732 6833
rect 1856 6935 1890 6969
rect 1856 6867 1890 6901
rect 1856 6799 1890 6833
rect 2030 6935 2064 6969
rect 2030 6867 2064 6901
rect 2030 6799 2064 6833
rect 2188 6935 2222 6969
rect 2188 6867 2222 6901
rect 2188 6799 2222 6833
rect 2372 6935 2406 6969
rect 2372 6867 2406 6901
rect 2372 6799 2406 6833
rect 2530 6935 2564 6969
rect 2530 6867 2564 6901
rect 2530 6799 2564 6833
rect 2776 6935 2810 6969
rect 2776 6867 2810 6901
rect 2776 6799 2810 6833
rect 2934 6935 2968 6969
rect 2934 6867 2968 6901
rect 2934 6799 2968 6833
rect 3120 6935 3154 6969
rect 3120 6867 3154 6901
rect 3120 6799 3154 6833
rect 3278 6935 3312 6969
rect 3278 6867 3312 6901
rect 3278 6799 3312 6833
rect 3742 6945 3776 6979
rect 3742 6877 3776 6911
rect 3742 6809 3776 6843
rect 3900 6945 3934 6979
rect 3900 6877 3934 6911
rect 3900 6809 3934 6843
rect 4050 6945 4084 6979
rect 4050 6877 4084 6911
rect 4050 6809 4084 6843
rect 4208 6945 4242 6979
rect 4208 6877 4242 6911
rect 4208 6809 4242 6843
rect 4402 6945 4436 6979
rect 4402 6877 4436 6911
rect 4402 6809 4436 6843
rect 4560 6945 4594 6979
rect 4560 6877 4594 6911
rect 4560 6809 4594 6843
rect 4710 6945 4744 6979
rect 4710 6877 4744 6911
rect 4710 6809 4744 6843
rect 4868 6945 4902 6979
rect 4868 6877 4902 6911
rect 4868 6809 4902 6843
rect 5700 6946 5734 6980
rect 5700 6878 5734 6912
rect 5700 6810 5734 6844
rect 5858 6946 5892 6980
rect 5858 6878 5892 6912
rect 5858 6810 5892 6844
rect 6008 6946 6042 6980
rect 6008 6878 6042 6912
rect 6008 6810 6042 6844
rect 6166 6946 6200 6980
rect 6166 6878 6200 6912
rect 6166 6810 6200 6844
rect 6360 6946 6394 6980
rect 6360 6878 6394 6912
rect 6360 6810 6394 6844
rect 6518 6946 6552 6980
rect 6518 6878 6552 6912
rect 6518 6810 6552 6844
rect 6668 6946 6702 6980
rect 6668 6878 6702 6912
rect 6668 6810 6702 6844
rect 6826 6946 6860 6980
rect 6826 6878 6860 6912
rect 6826 6810 6860 6844
rect 1410 5707 1444 5741
rect 1410 5639 1444 5673
rect 1410 5571 1444 5605
rect 1568 5707 1602 5741
rect 1568 5639 1602 5673
rect 1568 5571 1602 5605
rect 1698 5707 1732 5741
rect 1698 5639 1732 5673
rect 1698 5571 1732 5605
rect 1856 5707 1890 5741
rect 1856 5639 1890 5673
rect 1856 5571 1890 5605
rect 2030 5707 2064 5741
rect 2030 5639 2064 5673
rect 2030 5571 2064 5605
rect 2188 5707 2222 5741
rect 2188 5639 2222 5673
rect 2188 5571 2222 5605
rect 2372 5707 2406 5741
rect 2372 5639 2406 5673
rect 2372 5571 2406 5605
rect 2530 5707 2564 5741
rect 2530 5639 2564 5673
rect 2530 5571 2564 5605
rect 2776 5707 2810 5741
rect 2776 5639 2810 5673
rect 2776 5571 2810 5605
rect 2934 5707 2968 5741
rect 2934 5639 2968 5673
rect 2934 5571 2968 5605
rect 3120 5707 3154 5741
rect 3120 5639 3154 5673
rect 3120 5571 3154 5605
rect 3278 5707 3312 5741
rect 3278 5639 3312 5673
rect 3278 5571 3312 5605
rect 3742 5717 3776 5751
rect 3742 5649 3776 5683
rect 3742 5581 3776 5615
rect 3900 5717 3934 5751
rect 3900 5649 3934 5683
rect 3900 5581 3934 5615
rect 4050 5717 4084 5751
rect 4050 5649 4084 5683
rect 4050 5581 4084 5615
rect 4208 5717 4242 5751
rect 4208 5649 4242 5683
rect 4208 5581 4242 5615
rect 4402 5717 4436 5751
rect 4402 5649 4436 5683
rect 4402 5581 4436 5615
rect 4560 5717 4594 5751
rect 4560 5649 4594 5683
rect 4560 5581 4594 5615
rect 4710 5717 4744 5751
rect 4710 5649 4744 5683
rect 4710 5581 4744 5615
rect 4868 5717 4902 5751
rect 4868 5649 4902 5683
rect 4868 5581 4902 5615
rect 5700 5718 5734 5752
rect 5700 5650 5734 5684
rect 5700 5582 5734 5616
rect 5858 5718 5892 5752
rect 5858 5650 5892 5684
rect 5858 5582 5892 5616
rect 6008 5718 6042 5752
rect 6008 5650 6042 5684
rect 6008 5582 6042 5616
rect 6166 5718 6200 5752
rect 6166 5650 6200 5684
rect 6166 5582 6200 5616
rect 6360 5718 6394 5752
rect 6360 5650 6394 5684
rect 6360 5582 6394 5616
rect 6518 5718 6552 5752
rect 6518 5650 6552 5684
rect 6518 5582 6552 5616
rect 6668 5718 6702 5752
rect 6668 5650 6702 5684
rect 6668 5582 6702 5616
rect 6826 5718 6860 5752
rect 6826 5650 6860 5684
rect 6826 5582 6860 5616
rect 1410 4479 1444 4513
rect 1410 4411 1444 4445
rect 1410 4343 1444 4377
rect 1568 4479 1602 4513
rect 1568 4411 1602 4445
rect 1568 4343 1602 4377
rect 1698 4479 1732 4513
rect 1698 4411 1732 4445
rect 1698 4343 1732 4377
rect 1856 4479 1890 4513
rect 1856 4411 1890 4445
rect 1856 4343 1890 4377
rect 2030 4479 2064 4513
rect 2030 4411 2064 4445
rect 2030 4343 2064 4377
rect 2188 4479 2222 4513
rect 2188 4411 2222 4445
rect 2188 4343 2222 4377
rect 2372 4479 2406 4513
rect 2372 4411 2406 4445
rect 2372 4343 2406 4377
rect 2530 4479 2564 4513
rect 2530 4411 2564 4445
rect 2530 4343 2564 4377
rect 2776 4479 2810 4513
rect 2776 4411 2810 4445
rect 2776 4343 2810 4377
rect 2934 4479 2968 4513
rect 2934 4411 2968 4445
rect 2934 4343 2968 4377
rect 3120 4479 3154 4513
rect 3120 4411 3154 4445
rect 3120 4343 3154 4377
rect 3278 4479 3312 4513
rect 3278 4411 3312 4445
rect 3278 4343 3312 4377
rect 3742 4489 3776 4523
rect 3742 4421 3776 4455
rect 3742 4353 3776 4387
rect 3900 4489 3934 4523
rect 3900 4421 3934 4455
rect 3900 4353 3934 4387
rect 4050 4489 4084 4523
rect 4050 4421 4084 4455
rect 4050 4353 4084 4387
rect 4208 4489 4242 4523
rect 4208 4421 4242 4455
rect 4208 4353 4242 4387
rect 4402 4489 4436 4523
rect 4402 4421 4436 4455
rect 4402 4353 4436 4387
rect 4560 4489 4594 4523
rect 4560 4421 4594 4455
rect 4560 4353 4594 4387
rect 4710 4489 4744 4523
rect 4710 4421 4744 4455
rect 4710 4353 4744 4387
rect 4868 4489 4902 4523
rect 4868 4421 4902 4455
rect 4868 4353 4902 4387
rect 5700 4490 5734 4524
rect 5700 4422 5734 4456
rect 5700 4354 5734 4388
rect 5858 4490 5892 4524
rect 5858 4422 5892 4456
rect 5858 4354 5892 4388
rect 6008 4490 6042 4524
rect 6008 4422 6042 4456
rect 6008 4354 6042 4388
rect 6166 4490 6200 4524
rect 6166 4422 6200 4456
rect 6166 4354 6200 4388
rect 6360 4490 6394 4524
rect 6360 4422 6394 4456
rect 6360 4354 6394 4388
rect 6518 4490 6552 4524
rect 6518 4422 6552 4456
rect 6518 4354 6552 4388
rect 6668 4490 6702 4524
rect 6668 4422 6702 4456
rect 6668 4354 6702 4388
rect 6826 4490 6860 4524
rect 6826 4422 6860 4456
rect 6826 4354 6860 4388
rect 1410 3251 1444 3285
rect 1410 3183 1444 3217
rect 1410 3115 1444 3149
rect 1568 3251 1602 3285
rect 1568 3183 1602 3217
rect 1568 3115 1602 3149
rect 1698 3251 1732 3285
rect 1698 3183 1732 3217
rect 1698 3115 1732 3149
rect 1856 3251 1890 3285
rect 1856 3183 1890 3217
rect 1856 3115 1890 3149
rect 2030 3251 2064 3285
rect 2030 3183 2064 3217
rect 2030 3115 2064 3149
rect 2188 3251 2222 3285
rect 2188 3183 2222 3217
rect 2188 3115 2222 3149
rect 2372 3251 2406 3285
rect 2372 3183 2406 3217
rect 2372 3115 2406 3149
rect 2530 3251 2564 3285
rect 2530 3183 2564 3217
rect 2530 3115 2564 3149
rect 2776 3251 2810 3285
rect 2776 3183 2810 3217
rect 2776 3115 2810 3149
rect 2934 3251 2968 3285
rect 2934 3183 2968 3217
rect 2934 3115 2968 3149
rect 3120 3251 3154 3285
rect 3120 3183 3154 3217
rect 3120 3115 3154 3149
rect 3278 3251 3312 3285
rect 3278 3183 3312 3217
rect 3278 3115 3312 3149
rect 3742 3261 3776 3295
rect 3742 3193 3776 3227
rect 3742 3125 3776 3159
rect 3900 3261 3934 3295
rect 3900 3193 3934 3227
rect 3900 3125 3934 3159
rect 4050 3261 4084 3295
rect 4050 3193 4084 3227
rect 4050 3125 4084 3159
rect 4208 3261 4242 3295
rect 4208 3193 4242 3227
rect 4208 3125 4242 3159
rect 4402 3261 4436 3295
rect 4402 3193 4436 3227
rect 4402 3125 4436 3159
rect 4560 3261 4594 3295
rect 4560 3193 4594 3227
rect 4560 3125 4594 3159
rect 4710 3261 4744 3295
rect 4710 3193 4744 3227
rect 4710 3125 4744 3159
rect 4868 3261 4902 3295
rect 4868 3193 4902 3227
rect 4868 3125 4902 3159
rect 5700 3262 5734 3296
rect 5700 3194 5734 3228
rect 5700 3126 5734 3160
rect 5858 3262 5892 3296
rect 5858 3194 5892 3228
rect 5858 3126 5892 3160
rect 6008 3262 6042 3296
rect 6008 3194 6042 3228
rect 6008 3126 6042 3160
rect 6166 3262 6200 3296
rect 6166 3194 6200 3228
rect 6166 3126 6200 3160
rect 6360 3262 6394 3296
rect 6360 3194 6394 3228
rect 6360 3126 6394 3160
rect 6518 3262 6552 3296
rect 6518 3194 6552 3228
rect 6518 3126 6552 3160
rect 6668 3262 6702 3296
rect 6668 3194 6702 3228
rect 6668 3126 6702 3160
rect 6826 3262 6860 3296
rect 6826 3194 6860 3228
rect 6826 3126 6860 3160
rect 1410 2023 1444 2057
rect 1410 1955 1444 1989
rect 1410 1887 1444 1921
rect 1568 2023 1602 2057
rect 1568 1955 1602 1989
rect 1568 1887 1602 1921
rect 1698 2023 1732 2057
rect 1698 1955 1732 1989
rect 1698 1887 1732 1921
rect 1856 2023 1890 2057
rect 1856 1955 1890 1989
rect 1856 1887 1890 1921
rect 2030 2023 2064 2057
rect 2030 1955 2064 1989
rect 2030 1887 2064 1921
rect 2188 2023 2222 2057
rect 2188 1955 2222 1989
rect 2188 1887 2222 1921
rect 2372 2023 2406 2057
rect 2372 1955 2406 1989
rect 2372 1887 2406 1921
rect 2530 2023 2564 2057
rect 2530 1955 2564 1989
rect 2530 1887 2564 1921
rect 2776 2023 2810 2057
rect 2776 1955 2810 1989
rect 2776 1887 2810 1921
rect 2934 2023 2968 2057
rect 2934 1955 2968 1989
rect 2934 1887 2968 1921
rect 3120 2023 3154 2057
rect 3120 1955 3154 1989
rect 3120 1887 3154 1921
rect 3278 2023 3312 2057
rect 3278 1955 3312 1989
rect 3278 1887 3312 1921
rect 3742 2033 3776 2067
rect 3742 1965 3776 1999
rect 3742 1897 3776 1931
rect 3900 2033 3934 2067
rect 3900 1965 3934 1999
rect 3900 1897 3934 1931
rect 4050 2033 4084 2067
rect 4050 1965 4084 1999
rect 4050 1897 4084 1931
rect 4208 2033 4242 2067
rect 4208 1965 4242 1999
rect 4208 1897 4242 1931
rect 4402 2033 4436 2067
rect 4402 1965 4436 1999
rect 4402 1897 4436 1931
rect 4560 2033 4594 2067
rect 4560 1965 4594 1999
rect 4560 1897 4594 1931
rect 4710 2033 4744 2067
rect 4710 1965 4744 1999
rect 4710 1897 4744 1931
rect 4868 2033 4902 2067
rect 4868 1965 4902 1999
rect 4868 1897 4902 1931
rect 5700 2034 5734 2068
rect 5700 1966 5734 2000
rect 5700 1898 5734 1932
rect 5858 2034 5892 2068
rect 5858 1966 5892 2000
rect 5858 1898 5892 1932
rect 6008 2034 6042 2068
rect 6008 1966 6042 2000
rect 6008 1898 6042 1932
rect 6166 2034 6200 2068
rect 6166 1966 6200 2000
rect 6166 1898 6200 1932
rect 6360 2034 6394 2068
rect 6360 1966 6394 2000
rect 6360 1898 6394 1932
rect 6518 2034 6552 2068
rect 6518 1966 6552 2000
rect 6518 1898 6552 1932
rect 6668 2034 6702 2068
rect 6668 1966 6702 2000
rect 6668 1898 6702 1932
rect 6826 2034 6860 2068
rect 6826 1966 6860 2000
rect 6826 1898 6860 1932
rect 1410 795 1444 829
rect 1410 727 1444 761
rect 1410 659 1444 693
rect 1568 795 1602 829
rect 1568 727 1602 761
rect 1568 659 1602 693
rect 1698 795 1732 829
rect 1698 727 1732 761
rect 1698 659 1732 693
rect 1856 795 1890 829
rect 1856 727 1890 761
rect 1856 659 1890 693
rect 2030 795 2064 829
rect 2030 727 2064 761
rect 2030 659 2064 693
rect 2188 795 2222 829
rect 2188 727 2222 761
rect 2188 659 2222 693
rect 2372 795 2406 829
rect 2372 727 2406 761
rect 2372 659 2406 693
rect 2530 795 2564 829
rect 2530 727 2564 761
rect 2530 659 2564 693
rect 2776 795 2810 829
rect 2776 727 2810 761
rect 2776 659 2810 693
rect 2934 795 2968 829
rect 2934 727 2968 761
rect 2934 659 2968 693
rect 3120 795 3154 829
rect 3120 727 3154 761
rect 3120 659 3154 693
rect 3278 795 3312 829
rect 3278 727 3312 761
rect 3278 659 3312 693
rect 3742 805 3776 839
rect 3742 737 3776 771
rect 3742 669 3776 703
rect 3900 805 3934 839
rect 3900 737 3934 771
rect 3900 669 3934 703
rect 4050 805 4084 839
rect 4050 737 4084 771
rect 4050 669 4084 703
rect 4208 805 4242 839
rect 4208 737 4242 771
rect 4208 669 4242 703
rect 4402 805 4436 839
rect 4402 737 4436 771
rect 4402 669 4436 703
rect 4560 805 4594 839
rect 4560 737 4594 771
rect 4560 669 4594 703
rect 4710 805 4744 839
rect 4710 737 4744 771
rect 4710 669 4744 703
rect 4868 805 4902 839
rect 4868 737 4902 771
rect 4868 669 4902 703
<< psubdiff >>
rect 1324 18716 1959 18768
rect 1324 18682 1353 18716
rect 1387 18682 1421 18716
rect 1455 18682 1489 18716
rect 1523 18682 1557 18716
rect 1591 18682 1625 18716
rect 1659 18682 1693 18716
rect 1727 18682 1761 18716
rect 1795 18682 1829 18716
rect 1863 18682 1897 18716
rect 1931 18682 1959 18716
rect 1324 18640 1959 18682
rect 3704 18727 4244 18780
rect 3704 18693 3753 18727
rect 3787 18693 3821 18727
rect 3855 18693 3889 18727
rect 3923 18693 3957 18727
rect 3991 18693 4025 18727
rect 4059 18693 4093 18727
rect 4127 18693 4161 18727
rect 4195 18693 4244 18727
rect 3704 18640 4244 18693
rect 5662 18728 6202 18780
rect 5662 18694 5712 18728
rect 5746 18694 5780 18728
rect 5814 18694 5848 18728
rect 5882 18694 5916 18728
rect 5950 18694 5984 18728
rect 6018 18694 6052 18728
rect 6086 18694 6120 18728
rect 6154 18694 6202 18728
rect 5662 18640 6202 18694
rect 1324 17488 1959 17540
rect 1324 17454 1353 17488
rect 1387 17454 1421 17488
rect 1455 17454 1489 17488
rect 1523 17454 1557 17488
rect 1591 17454 1625 17488
rect 1659 17454 1693 17488
rect 1727 17454 1761 17488
rect 1795 17454 1829 17488
rect 1863 17454 1897 17488
rect 1931 17454 1959 17488
rect 1324 17412 1959 17454
rect 3704 17499 4244 17552
rect 3704 17465 3753 17499
rect 3787 17465 3821 17499
rect 3855 17465 3889 17499
rect 3923 17465 3957 17499
rect 3991 17465 4025 17499
rect 4059 17465 4093 17499
rect 4127 17465 4161 17499
rect 4195 17465 4244 17499
rect 3704 17412 4244 17465
rect 5662 17500 6202 17552
rect 5662 17466 5712 17500
rect 5746 17466 5780 17500
rect 5814 17466 5848 17500
rect 5882 17466 5916 17500
rect 5950 17466 5984 17500
rect 6018 17466 6052 17500
rect 6086 17466 6120 17500
rect 6154 17466 6202 17500
rect 5662 17412 6202 17466
rect 1324 16260 1959 16312
rect 1324 16226 1353 16260
rect 1387 16226 1421 16260
rect 1455 16226 1489 16260
rect 1523 16226 1557 16260
rect 1591 16226 1625 16260
rect 1659 16226 1693 16260
rect 1727 16226 1761 16260
rect 1795 16226 1829 16260
rect 1863 16226 1897 16260
rect 1931 16226 1959 16260
rect 1324 16184 1959 16226
rect 3704 16271 4244 16324
rect 3704 16237 3753 16271
rect 3787 16237 3821 16271
rect 3855 16237 3889 16271
rect 3923 16237 3957 16271
rect 3991 16237 4025 16271
rect 4059 16237 4093 16271
rect 4127 16237 4161 16271
rect 4195 16237 4244 16271
rect 3704 16184 4244 16237
rect 5662 16272 6202 16324
rect 5662 16238 5712 16272
rect 5746 16238 5780 16272
rect 5814 16238 5848 16272
rect 5882 16238 5916 16272
rect 5950 16238 5984 16272
rect 6018 16238 6052 16272
rect 6086 16238 6120 16272
rect 6154 16238 6202 16272
rect 5662 16184 6202 16238
rect 1324 15032 1959 15084
rect 1324 14998 1353 15032
rect 1387 14998 1421 15032
rect 1455 14998 1489 15032
rect 1523 14998 1557 15032
rect 1591 14998 1625 15032
rect 1659 14998 1693 15032
rect 1727 14998 1761 15032
rect 1795 14998 1829 15032
rect 1863 14998 1897 15032
rect 1931 14998 1959 15032
rect 1324 14956 1959 14998
rect 3704 15043 4244 15096
rect 3704 15009 3753 15043
rect 3787 15009 3821 15043
rect 3855 15009 3889 15043
rect 3923 15009 3957 15043
rect 3991 15009 4025 15043
rect 4059 15009 4093 15043
rect 4127 15009 4161 15043
rect 4195 15009 4244 15043
rect 3704 14956 4244 15009
rect 5662 15044 6202 15096
rect 5662 15010 5712 15044
rect 5746 15010 5780 15044
rect 5814 15010 5848 15044
rect 5882 15010 5916 15044
rect 5950 15010 5984 15044
rect 6018 15010 6052 15044
rect 6086 15010 6120 15044
rect 6154 15010 6202 15044
rect 5662 14956 6202 15010
rect 1324 13804 1959 13856
rect 1324 13770 1353 13804
rect 1387 13770 1421 13804
rect 1455 13770 1489 13804
rect 1523 13770 1557 13804
rect 1591 13770 1625 13804
rect 1659 13770 1693 13804
rect 1727 13770 1761 13804
rect 1795 13770 1829 13804
rect 1863 13770 1897 13804
rect 1931 13770 1959 13804
rect 1324 13728 1959 13770
rect 3704 13815 4244 13868
rect 3704 13781 3753 13815
rect 3787 13781 3821 13815
rect 3855 13781 3889 13815
rect 3923 13781 3957 13815
rect 3991 13781 4025 13815
rect 4059 13781 4093 13815
rect 4127 13781 4161 13815
rect 4195 13781 4244 13815
rect 3704 13728 4244 13781
rect 5662 13816 6202 13868
rect 5662 13782 5712 13816
rect 5746 13782 5780 13816
rect 5814 13782 5848 13816
rect 5882 13782 5916 13816
rect 5950 13782 5984 13816
rect 6018 13782 6052 13816
rect 6086 13782 6120 13816
rect 6154 13782 6202 13816
rect 5662 13728 6202 13782
rect 1324 12576 1959 12628
rect 1324 12542 1353 12576
rect 1387 12542 1421 12576
rect 1455 12542 1489 12576
rect 1523 12542 1557 12576
rect 1591 12542 1625 12576
rect 1659 12542 1693 12576
rect 1727 12542 1761 12576
rect 1795 12542 1829 12576
rect 1863 12542 1897 12576
rect 1931 12542 1959 12576
rect 1324 12500 1959 12542
rect 3704 12587 4244 12640
rect 3704 12553 3753 12587
rect 3787 12553 3821 12587
rect 3855 12553 3889 12587
rect 3923 12553 3957 12587
rect 3991 12553 4025 12587
rect 4059 12553 4093 12587
rect 4127 12553 4161 12587
rect 4195 12553 4244 12587
rect 3704 12500 4244 12553
rect 5662 12588 6202 12640
rect 5662 12554 5712 12588
rect 5746 12554 5780 12588
rect 5814 12554 5848 12588
rect 5882 12554 5916 12588
rect 5950 12554 5984 12588
rect 6018 12554 6052 12588
rect 6086 12554 6120 12588
rect 6154 12554 6202 12588
rect 5662 12500 6202 12554
rect 1324 11348 1959 11400
rect 1324 11314 1353 11348
rect 1387 11314 1421 11348
rect 1455 11314 1489 11348
rect 1523 11314 1557 11348
rect 1591 11314 1625 11348
rect 1659 11314 1693 11348
rect 1727 11314 1761 11348
rect 1795 11314 1829 11348
rect 1863 11314 1897 11348
rect 1931 11314 1959 11348
rect 1324 11272 1959 11314
rect 3704 11359 4244 11412
rect 3704 11325 3753 11359
rect 3787 11325 3821 11359
rect 3855 11325 3889 11359
rect 3923 11325 3957 11359
rect 3991 11325 4025 11359
rect 4059 11325 4093 11359
rect 4127 11325 4161 11359
rect 4195 11325 4244 11359
rect 3704 11272 4244 11325
rect 5662 11360 6202 11412
rect 5662 11326 5712 11360
rect 5746 11326 5780 11360
rect 5814 11326 5848 11360
rect 5882 11326 5916 11360
rect 5950 11326 5984 11360
rect 6018 11326 6052 11360
rect 6086 11326 6120 11360
rect 6154 11326 6202 11360
rect 5662 11272 6202 11326
rect 1324 10120 1959 10172
rect 1324 10086 1353 10120
rect 1387 10086 1421 10120
rect 1455 10086 1489 10120
rect 1523 10086 1557 10120
rect 1591 10086 1625 10120
rect 1659 10086 1693 10120
rect 1727 10086 1761 10120
rect 1795 10086 1829 10120
rect 1863 10086 1897 10120
rect 1931 10086 1959 10120
rect 1324 10044 1959 10086
rect 3704 10131 4244 10184
rect 3704 10097 3753 10131
rect 3787 10097 3821 10131
rect 3855 10097 3889 10131
rect 3923 10097 3957 10131
rect 3991 10097 4025 10131
rect 4059 10097 4093 10131
rect 4127 10097 4161 10131
rect 4195 10097 4244 10131
rect 3704 10044 4244 10097
rect 5662 10132 6202 10184
rect 5662 10098 5712 10132
rect 5746 10098 5780 10132
rect 5814 10098 5848 10132
rect 5882 10098 5916 10132
rect 5950 10098 5984 10132
rect 6018 10098 6052 10132
rect 6086 10098 6120 10132
rect 6154 10098 6202 10132
rect 5662 10044 6202 10098
rect 1324 8892 1959 8944
rect 1324 8858 1353 8892
rect 1387 8858 1421 8892
rect 1455 8858 1489 8892
rect 1523 8858 1557 8892
rect 1591 8858 1625 8892
rect 1659 8858 1693 8892
rect 1727 8858 1761 8892
rect 1795 8858 1829 8892
rect 1863 8858 1897 8892
rect 1931 8858 1959 8892
rect 1324 8816 1959 8858
rect 3704 8903 4244 8956
rect 3704 8869 3753 8903
rect 3787 8869 3821 8903
rect 3855 8869 3889 8903
rect 3923 8869 3957 8903
rect 3991 8869 4025 8903
rect 4059 8869 4093 8903
rect 4127 8869 4161 8903
rect 4195 8869 4244 8903
rect 3704 8816 4244 8869
rect 5662 8904 6202 8956
rect 5662 8870 5712 8904
rect 5746 8870 5780 8904
rect 5814 8870 5848 8904
rect 5882 8870 5916 8904
rect 5950 8870 5984 8904
rect 6018 8870 6052 8904
rect 6086 8870 6120 8904
rect 6154 8870 6202 8904
rect 5662 8816 6202 8870
rect 1324 7664 1959 7716
rect 1324 7630 1353 7664
rect 1387 7630 1421 7664
rect 1455 7630 1489 7664
rect 1523 7630 1557 7664
rect 1591 7630 1625 7664
rect 1659 7630 1693 7664
rect 1727 7630 1761 7664
rect 1795 7630 1829 7664
rect 1863 7630 1897 7664
rect 1931 7630 1959 7664
rect 1324 7588 1959 7630
rect 3704 7675 4244 7728
rect 3704 7641 3753 7675
rect 3787 7641 3821 7675
rect 3855 7641 3889 7675
rect 3923 7641 3957 7675
rect 3991 7641 4025 7675
rect 4059 7641 4093 7675
rect 4127 7641 4161 7675
rect 4195 7641 4244 7675
rect 3704 7588 4244 7641
rect 5662 7676 6202 7728
rect 5662 7642 5712 7676
rect 5746 7642 5780 7676
rect 5814 7642 5848 7676
rect 5882 7642 5916 7676
rect 5950 7642 5984 7676
rect 6018 7642 6052 7676
rect 6086 7642 6120 7676
rect 6154 7642 6202 7676
rect 5662 7588 6202 7642
rect 1324 6436 1959 6488
rect 1324 6402 1353 6436
rect 1387 6402 1421 6436
rect 1455 6402 1489 6436
rect 1523 6402 1557 6436
rect 1591 6402 1625 6436
rect 1659 6402 1693 6436
rect 1727 6402 1761 6436
rect 1795 6402 1829 6436
rect 1863 6402 1897 6436
rect 1931 6402 1959 6436
rect 1324 6360 1959 6402
rect 3704 6447 4244 6500
rect 3704 6413 3753 6447
rect 3787 6413 3821 6447
rect 3855 6413 3889 6447
rect 3923 6413 3957 6447
rect 3991 6413 4025 6447
rect 4059 6413 4093 6447
rect 4127 6413 4161 6447
rect 4195 6413 4244 6447
rect 3704 6360 4244 6413
rect 5662 6448 6202 6500
rect 5662 6414 5712 6448
rect 5746 6414 5780 6448
rect 5814 6414 5848 6448
rect 5882 6414 5916 6448
rect 5950 6414 5984 6448
rect 6018 6414 6052 6448
rect 6086 6414 6120 6448
rect 6154 6414 6202 6448
rect 5662 6360 6202 6414
rect 1324 5208 1959 5260
rect 1324 5174 1353 5208
rect 1387 5174 1421 5208
rect 1455 5174 1489 5208
rect 1523 5174 1557 5208
rect 1591 5174 1625 5208
rect 1659 5174 1693 5208
rect 1727 5174 1761 5208
rect 1795 5174 1829 5208
rect 1863 5174 1897 5208
rect 1931 5174 1959 5208
rect 1324 5132 1959 5174
rect 3704 5219 4244 5272
rect 3704 5185 3753 5219
rect 3787 5185 3821 5219
rect 3855 5185 3889 5219
rect 3923 5185 3957 5219
rect 3991 5185 4025 5219
rect 4059 5185 4093 5219
rect 4127 5185 4161 5219
rect 4195 5185 4244 5219
rect 3704 5132 4244 5185
rect 5662 5220 6202 5272
rect 5662 5186 5712 5220
rect 5746 5186 5780 5220
rect 5814 5186 5848 5220
rect 5882 5186 5916 5220
rect 5950 5186 5984 5220
rect 6018 5186 6052 5220
rect 6086 5186 6120 5220
rect 6154 5186 6202 5220
rect 5662 5132 6202 5186
rect 1324 3980 1959 4032
rect 1324 3946 1353 3980
rect 1387 3946 1421 3980
rect 1455 3946 1489 3980
rect 1523 3946 1557 3980
rect 1591 3946 1625 3980
rect 1659 3946 1693 3980
rect 1727 3946 1761 3980
rect 1795 3946 1829 3980
rect 1863 3946 1897 3980
rect 1931 3946 1959 3980
rect 1324 3904 1959 3946
rect 3704 3991 4244 4044
rect 3704 3957 3753 3991
rect 3787 3957 3821 3991
rect 3855 3957 3889 3991
rect 3923 3957 3957 3991
rect 3991 3957 4025 3991
rect 4059 3957 4093 3991
rect 4127 3957 4161 3991
rect 4195 3957 4244 3991
rect 3704 3904 4244 3957
rect 5662 3992 6202 4044
rect 5662 3958 5712 3992
rect 5746 3958 5780 3992
rect 5814 3958 5848 3992
rect 5882 3958 5916 3992
rect 5950 3958 5984 3992
rect 6018 3958 6052 3992
rect 6086 3958 6120 3992
rect 6154 3958 6202 3992
rect 5662 3904 6202 3958
rect 1324 2752 1959 2804
rect 1324 2718 1353 2752
rect 1387 2718 1421 2752
rect 1455 2718 1489 2752
rect 1523 2718 1557 2752
rect 1591 2718 1625 2752
rect 1659 2718 1693 2752
rect 1727 2718 1761 2752
rect 1795 2718 1829 2752
rect 1863 2718 1897 2752
rect 1931 2718 1959 2752
rect 1324 2676 1959 2718
rect 3704 2763 4244 2816
rect 3704 2729 3753 2763
rect 3787 2729 3821 2763
rect 3855 2729 3889 2763
rect 3923 2729 3957 2763
rect 3991 2729 4025 2763
rect 4059 2729 4093 2763
rect 4127 2729 4161 2763
rect 4195 2729 4244 2763
rect 3704 2676 4244 2729
rect 5662 2764 6202 2816
rect 5662 2730 5712 2764
rect 5746 2730 5780 2764
rect 5814 2730 5848 2764
rect 5882 2730 5916 2764
rect 5950 2730 5984 2764
rect 6018 2730 6052 2764
rect 6086 2730 6120 2764
rect 6154 2730 6202 2764
rect 5662 2676 6202 2730
rect 1324 1524 1959 1576
rect 1324 1490 1353 1524
rect 1387 1490 1421 1524
rect 1455 1490 1489 1524
rect 1523 1490 1557 1524
rect 1591 1490 1625 1524
rect 1659 1490 1693 1524
rect 1727 1490 1761 1524
rect 1795 1490 1829 1524
rect 1863 1490 1897 1524
rect 1931 1490 1959 1524
rect 1324 1448 1959 1490
rect 3704 1535 4244 1588
rect 3704 1501 3753 1535
rect 3787 1501 3821 1535
rect 3855 1501 3889 1535
rect 3923 1501 3957 1535
rect 3991 1501 4025 1535
rect 4059 1501 4093 1535
rect 4127 1501 4161 1535
rect 4195 1501 4244 1535
rect 3704 1448 4244 1501
rect 5662 1536 6202 1588
rect 5662 1502 5712 1536
rect 5746 1502 5780 1536
rect 5814 1502 5848 1536
rect 5882 1502 5916 1536
rect 5950 1502 5984 1536
rect 6018 1502 6052 1536
rect 6086 1502 6120 1536
rect 6154 1502 6202 1536
rect 5662 1448 6202 1502
rect 1324 296 1959 348
rect 1324 262 1353 296
rect 1387 262 1421 296
rect 1455 262 1489 296
rect 1523 262 1557 296
rect 1591 262 1625 296
rect 1659 262 1693 296
rect 1727 262 1761 296
rect 1795 262 1829 296
rect 1863 262 1897 296
rect 1931 262 1959 296
rect 1324 220 1959 262
rect 3704 307 4244 360
rect 3704 273 3753 307
rect 3787 273 3821 307
rect 3855 273 3889 307
rect 3923 273 3957 307
rect 3991 273 4025 307
rect 4059 273 4093 307
rect 4127 273 4161 307
rect 4195 273 4244 307
rect 3704 220 4244 273
<< mvnsubdiff >>
rect 1348 19418 1880 19470
rect 1348 19384 1395 19418
rect 1429 19384 1463 19418
rect 1497 19384 1531 19418
rect 1565 19384 1599 19418
rect 1633 19384 1667 19418
rect 1701 19384 1735 19418
rect 1769 19384 1803 19418
rect 1837 19384 1880 19418
rect 1348 19330 1880 19384
rect 3734 19417 4254 19460
rect 3734 19383 3773 19417
rect 3807 19383 3841 19417
rect 3875 19383 3909 19417
rect 3943 19383 3977 19417
rect 4011 19383 4045 19417
rect 4079 19383 4113 19417
rect 4147 19383 4181 19417
rect 4215 19383 4254 19417
rect 3734 19340 4254 19383
rect 5692 19416 6212 19460
rect 5692 19382 5732 19416
rect 5766 19382 5800 19416
rect 5834 19382 5868 19416
rect 5902 19382 5936 19416
rect 5970 19382 6004 19416
rect 6038 19382 6072 19416
rect 6106 19382 6140 19416
rect 6174 19382 6212 19416
rect 5692 19340 6212 19382
rect 1348 18190 1880 18242
rect 1348 18156 1395 18190
rect 1429 18156 1463 18190
rect 1497 18156 1531 18190
rect 1565 18156 1599 18190
rect 1633 18156 1667 18190
rect 1701 18156 1735 18190
rect 1769 18156 1803 18190
rect 1837 18156 1880 18190
rect 1348 18102 1880 18156
rect 3734 18189 4254 18232
rect 3734 18155 3773 18189
rect 3807 18155 3841 18189
rect 3875 18155 3909 18189
rect 3943 18155 3977 18189
rect 4011 18155 4045 18189
rect 4079 18155 4113 18189
rect 4147 18155 4181 18189
rect 4215 18155 4254 18189
rect 3734 18112 4254 18155
rect 5692 18188 6212 18232
rect 5692 18154 5732 18188
rect 5766 18154 5800 18188
rect 5834 18154 5868 18188
rect 5902 18154 5936 18188
rect 5970 18154 6004 18188
rect 6038 18154 6072 18188
rect 6106 18154 6140 18188
rect 6174 18154 6212 18188
rect 5692 18112 6212 18154
rect 1348 16962 1880 17014
rect 1348 16928 1395 16962
rect 1429 16928 1463 16962
rect 1497 16928 1531 16962
rect 1565 16928 1599 16962
rect 1633 16928 1667 16962
rect 1701 16928 1735 16962
rect 1769 16928 1803 16962
rect 1837 16928 1880 16962
rect 1348 16874 1880 16928
rect 3734 16961 4254 17004
rect 3734 16927 3773 16961
rect 3807 16927 3841 16961
rect 3875 16927 3909 16961
rect 3943 16927 3977 16961
rect 4011 16927 4045 16961
rect 4079 16927 4113 16961
rect 4147 16927 4181 16961
rect 4215 16927 4254 16961
rect 3734 16884 4254 16927
rect 5692 16960 6212 17004
rect 5692 16926 5732 16960
rect 5766 16926 5800 16960
rect 5834 16926 5868 16960
rect 5902 16926 5936 16960
rect 5970 16926 6004 16960
rect 6038 16926 6072 16960
rect 6106 16926 6140 16960
rect 6174 16926 6212 16960
rect 5692 16884 6212 16926
rect 1348 15734 1880 15786
rect 1348 15700 1395 15734
rect 1429 15700 1463 15734
rect 1497 15700 1531 15734
rect 1565 15700 1599 15734
rect 1633 15700 1667 15734
rect 1701 15700 1735 15734
rect 1769 15700 1803 15734
rect 1837 15700 1880 15734
rect 1348 15646 1880 15700
rect 3734 15733 4254 15776
rect 3734 15699 3773 15733
rect 3807 15699 3841 15733
rect 3875 15699 3909 15733
rect 3943 15699 3977 15733
rect 4011 15699 4045 15733
rect 4079 15699 4113 15733
rect 4147 15699 4181 15733
rect 4215 15699 4254 15733
rect 3734 15656 4254 15699
rect 5692 15732 6212 15776
rect 5692 15698 5732 15732
rect 5766 15698 5800 15732
rect 5834 15698 5868 15732
rect 5902 15698 5936 15732
rect 5970 15698 6004 15732
rect 6038 15698 6072 15732
rect 6106 15698 6140 15732
rect 6174 15698 6212 15732
rect 5692 15656 6212 15698
rect 1348 14506 1880 14558
rect 1348 14472 1395 14506
rect 1429 14472 1463 14506
rect 1497 14472 1531 14506
rect 1565 14472 1599 14506
rect 1633 14472 1667 14506
rect 1701 14472 1735 14506
rect 1769 14472 1803 14506
rect 1837 14472 1880 14506
rect 1348 14418 1880 14472
rect 3734 14505 4254 14548
rect 3734 14471 3773 14505
rect 3807 14471 3841 14505
rect 3875 14471 3909 14505
rect 3943 14471 3977 14505
rect 4011 14471 4045 14505
rect 4079 14471 4113 14505
rect 4147 14471 4181 14505
rect 4215 14471 4254 14505
rect 3734 14428 4254 14471
rect 5692 14504 6212 14548
rect 5692 14470 5732 14504
rect 5766 14470 5800 14504
rect 5834 14470 5868 14504
rect 5902 14470 5936 14504
rect 5970 14470 6004 14504
rect 6038 14470 6072 14504
rect 6106 14470 6140 14504
rect 6174 14470 6212 14504
rect 5692 14428 6212 14470
rect 1348 13278 1880 13330
rect 1348 13244 1395 13278
rect 1429 13244 1463 13278
rect 1497 13244 1531 13278
rect 1565 13244 1599 13278
rect 1633 13244 1667 13278
rect 1701 13244 1735 13278
rect 1769 13244 1803 13278
rect 1837 13244 1880 13278
rect 1348 13190 1880 13244
rect 3734 13277 4254 13320
rect 3734 13243 3773 13277
rect 3807 13243 3841 13277
rect 3875 13243 3909 13277
rect 3943 13243 3977 13277
rect 4011 13243 4045 13277
rect 4079 13243 4113 13277
rect 4147 13243 4181 13277
rect 4215 13243 4254 13277
rect 3734 13200 4254 13243
rect 5692 13276 6212 13320
rect 5692 13242 5732 13276
rect 5766 13242 5800 13276
rect 5834 13242 5868 13276
rect 5902 13242 5936 13276
rect 5970 13242 6004 13276
rect 6038 13242 6072 13276
rect 6106 13242 6140 13276
rect 6174 13242 6212 13276
rect 5692 13200 6212 13242
rect 1348 12050 1880 12102
rect 1348 12016 1395 12050
rect 1429 12016 1463 12050
rect 1497 12016 1531 12050
rect 1565 12016 1599 12050
rect 1633 12016 1667 12050
rect 1701 12016 1735 12050
rect 1769 12016 1803 12050
rect 1837 12016 1880 12050
rect 1348 11962 1880 12016
rect 3734 12049 4254 12092
rect 3734 12015 3773 12049
rect 3807 12015 3841 12049
rect 3875 12015 3909 12049
rect 3943 12015 3977 12049
rect 4011 12015 4045 12049
rect 4079 12015 4113 12049
rect 4147 12015 4181 12049
rect 4215 12015 4254 12049
rect 3734 11972 4254 12015
rect 5692 12048 6212 12092
rect 5692 12014 5732 12048
rect 5766 12014 5800 12048
rect 5834 12014 5868 12048
rect 5902 12014 5936 12048
rect 5970 12014 6004 12048
rect 6038 12014 6072 12048
rect 6106 12014 6140 12048
rect 6174 12014 6212 12048
rect 5692 11972 6212 12014
rect 1348 10822 1880 10874
rect 1348 10788 1395 10822
rect 1429 10788 1463 10822
rect 1497 10788 1531 10822
rect 1565 10788 1599 10822
rect 1633 10788 1667 10822
rect 1701 10788 1735 10822
rect 1769 10788 1803 10822
rect 1837 10788 1880 10822
rect 1348 10734 1880 10788
rect 3734 10821 4254 10864
rect 3734 10787 3773 10821
rect 3807 10787 3841 10821
rect 3875 10787 3909 10821
rect 3943 10787 3977 10821
rect 4011 10787 4045 10821
rect 4079 10787 4113 10821
rect 4147 10787 4181 10821
rect 4215 10787 4254 10821
rect 3734 10744 4254 10787
rect 5692 10820 6212 10864
rect 5692 10786 5732 10820
rect 5766 10786 5800 10820
rect 5834 10786 5868 10820
rect 5902 10786 5936 10820
rect 5970 10786 6004 10820
rect 6038 10786 6072 10820
rect 6106 10786 6140 10820
rect 6174 10786 6212 10820
rect 5692 10744 6212 10786
rect 1348 9594 1880 9646
rect 1348 9560 1395 9594
rect 1429 9560 1463 9594
rect 1497 9560 1531 9594
rect 1565 9560 1599 9594
rect 1633 9560 1667 9594
rect 1701 9560 1735 9594
rect 1769 9560 1803 9594
rect 1837 9560 1880 9594
rect 1348 9506 1880 9560
rect 3734 9593 4254 9636
rect 3734 9559 3773 9593
rect 3807 9559 3841 9593
rect 3875 9559 3909 9593
rect 3943 9559 3977 9593
rect 4011 9559 4045 9593
rect 4079 9559 4113 9593
rect 4147 9559 4181 9593
rect 4215 9559 4254 9593
rect 3734 9516 4254 9559
rect 5692 9592 6212 9636
rect 5692 9558 5732 9592
rect 5766 9558 5800 9592
rect 5834 9558 5868 9592
rect 5902 9558 5936 9592
rect 5970 9558 6004 9592
rect 6038 9558 6072 9592
rect 6106 9558 6140 9592
rect 6174 9558 6212 9592
rect 5692 9516 6212 9558
rect 1348 8366 1880 8418
rect 1348 8332 1395 8366
rect 1429 8332 1463 8366
rect 1497 8332 1531 8366
rect 1565 8332 1599 8366
rect 1633 8332 1667 8366
rect 1701 8332 1735 8366
rect 1769 8332 1803 8366
rect 1837 8332 1880 8366
rect 1348 8278 1880 8332
rect 3734 8365 4254 8408
rect 3734 8331 3773 8365
rect 3807 8331 3841 8365
rect 3875 8331 3909 8365
rect 3943 8331 3977 8365
rect 4011 8331 4045 8365
rect 4079 8331 4113 8365
rect 4147 8331 4181 8365
rect 4215 8331 4254 8365
rect 3734 8288 4254 8331
rect 5692 8364 6212 8408
rect 5692 8330 5732 8364
rect 5766 8330 5800 8364
rect 5834 8330 5868 8364
rect 5902 8330 5936 8364
rect 5970 8330 6004 8364
rect 6038 8330 6072 8364
rect 6106 8330 6140 8364
rect 6174 8330 6212 8364
rect 5692 8288 6212 8330
rect 1348 7138 1880 7190
rect 1348 7104 1395 7138
rect 1429 7104 1463 7138
rect 1497 7104 1531 7138
rect 1565 7104 1599 7138
rect 1633 7104 1667 7138
rect 1701 7104 1735 7138
rect 1769 7104 1803 7138
rect 1837 7104 1880 7138
rect 1348 7050 1880 7104
rect 3734 7137 4254 7180
rect 3734 7103 3773 7137
rect 3807 7103 3841 7137
rect 3875 7103 3909 7137
rect 3943 7103 3977 7137
rect 4011 7103 4045 7137
rect 4079 7103 4113 7137
rect 4147 7103 4181 7137
rect 4215 7103 4254 7137
rect 3734 7060 4254 7103
rect 5692 7136 6212 7180
rect 5692 7102 5732 7136
rect 5766 7102 5800 7136
rect 5834 7102 5868 7136
rect 5902 7102 5936 7136
rect 5970 7102 6004 7136
rect 6038 7102 6072 7136
rect 6106 7102 6140 7136
rect 6174 7102 6212 7136
rect 5692 7060 6212 7102
rect 1348 5910 1880 5962
rect 1348 5876 1395 5910
rect 1429 5876 1463 5910
rect 1497 5876 1531 5910
rect 1565 5876 1599 5910
rect 1633 5876 1667 5910
rect 1701 5876 1735 5910
rect 1769 5876 1803 5910
rect 1837 5876 1880 5910
rect 1348 5822 1880 5876
rect 3734 5909 4254 5952
rect 3734 5875 3773 5909
rect 3807 5875 3841 5909
rect 3875 5875 3909 5909
rect 3943 5875 3977 5909
rect 4011 5875 4045 5909
rect 4079 5875 4113 5909
rect 4147 5875 4181 5909
rect 4215 5875 4254 5909
rect 3734 5832 4254 5875
rect 5692 5908 6212 5952
rect 5692 5874 5732 5908
rect 5766 5874 5800 5908
rect 5834 5874 5868 5908
rect 5902 5874 5936 5908
rect 5970 5874 6004 5908
rect 6038 5874 6072 5908
rect 6106 5874 6140 5908
rect 6174 5874 6212 5908
rect 5692 5832 6212 5874
rect 1348 4682 1880 4734
rect 1348 4648 1395 4682
rect 1429 4648 1463 4682
rect 1497 4648 1531 4682
rect 1565 4648 1599 4682
rect 1633 4648 1667 4682
rect 1701 4648 1735 4682
rect 1769 4648 1803 4682
rect 1837 4648 1880 4682
rect 1348 4594 1880 4648
rect 3734 4681 4254 4724
rect 3734 4647 3773 4681
rect 3807 4647 3841 4681
rect 3875 4647 3909 4681
rect 3943 4647 3977 4681
rect 4011 4647 4045 4681
rect 4079 4647 4113 4681
rect 4147 4647 4181 4681
rect 4215 4647 4254 4681
rect 3734 4604 4254 4647
rect 5692 4680 6212 4724
rect 5692 4646 5732 4680
rect 5766 4646 5800 4680
rect 5834 4646 5868 4680
rect 5902 4646 5936 4680
rect 5970 4646 6004 4680
rect 6038 4646 6072 4680
rect 6106 4646 6140 4680
rect 6174 4646 6212 4680
rect 5692 4604 6212 4646
rect 1348 3454 1880 3506
rect 1348 3420 1395 3454
rect 1429 3420 1463 3454
rect 1497 3420 1531 3454
rect 1565 3420 1599 3454
rect 1633 3420 1667 3454
rect 1701 3420 1735 3454
rect 1769 3420 1803 3454
rect 1837 3420 1880 3454
rect 1348 3366 1880 3420
rect 3734 3453 4254 3496
rect 3734 3419 3773 3453
rect 3807 3419 3841 3453
rect 3875 3419 3909 3453
rect 3943 3419 3977 3453
rect 4011 3419 4045 3453
rect 4079 3419 4113 3453
rect 4147 3419 4181 3453
rect 4215 3419 4254 3453
rect 3734 3376 4254 3419
rect 5692 3452 6212 3496
rect 5692 3418 5732 3452
rect 5766 3418 5800 3452
rect 5834 3418 5868 3452
rect 5902 3418 5936 3452
rect 5970 3418 6004 3452
rect 6038 3418 6072 3452
rect 6106 3418 6140 3452
rect 6174 3418 6212 3452
rect 5692 3376 6212 3418
rect 1348 2226 1880 2278
rect 1348 2192 1395 2226
rect 1429 2192 1463 2226
rect 1497 2192 1531 2226
rect 1565 2192 1599 2226
rect 1633 2192 1667 2226
rect 1701 2192 1735 2226
rect 1769 2192 1803 2226
rect 1837 2192 1880 2226
rect 1348 2138 1880 2192
rect 3734 2225 4254 2268
rect 3734 2191 3773 2225
rect 3807 2191 3841 2225
rect 3875 2191 3909 2225
rect 3943 2191 3977 2225
rect 4011 2191 4045 2225
rect 4079 2191 4113 2225
rect 4147 2191 4181 2225
rect 4215 2191 4254 2225
rect 3734 2148 4254 2191
rect 5692 2224 6212 2268
rect 5692 2190 5732 2224
rect 5766 2190 5800 2224
rect 5834 2190 5868 2224
rect 5902 2190 5936 2224
rect 5970 2190 6004 2224
rect 6038 2190 6072 2224
rect 6106 2190 6140 2224
rect 6174 2190 6212 2224
rect 5692 2148 6212 2190
rect 1348 998 1880 1050
rect 1348 964 1395 998
rect 1429 964 1463 998
rect 1497 964 1531 998
rect 1565 964 1599 998
rect 1633 964 1667 998
rect 1701 964 1735 998
rect 1769 964 1803 998
rect 1837 964 1880 998
rect 1348 910 1880 964
rect 3734 997 4254 1040
rect 3734 963 3773 997
rect 3807 963 3841 997
rect 3875 963 3909 997
rect 3943 963 3977 997
rect 4011 963 4045 997
rect 4079 963 4113 997
rect 4147 963 4181 997
rect 4215 963 4254 997
rect 3734 920 4254 963
<< psubdiffcont >>
rect 1353 18682 1387 18716
rect 1421 18682 1455 18716
rect 1489 18682 1523 18716
rect 1557 18682 1591 18716
rect 1625 18682 1659 18716
rect 1693 18682 1727 18716
rect 1761 18682 1795 18716
rect 1829 18682 1863 18716
rect 1897 18682 1931 18716
rect 3753 18693 3787 18727
rect 3821 18693 3855 18727
rect 3889 18693 3923 18727
rect 3957 18693 3991 18727
rect 4025 18693 4059 18727
rect 4093 18693 4127 18727
rect 4161 18693 4195 18727
rect 5712 18694 5746 18728
rect 5780 18694 5814 18728
rect 5848 18694 5882 18728
rect 5916 18694 5950 18728
rect 5984 18694 6018 18728
rect 6052 18694 6086 18728
rect 6120 18694 6154 18728
rect 1353 17454 1387 17488
rect 1421 17454 1455 17488
rect 1489 17454 1523 17488
rect 1557 17454 1591 17488
rect 1625 17454 1659 17488
rect 1693 17454 1727 17488
rect 1761 17454 1795 17488
rect 1829 17454 1863 17488
rect 1897 17454 1931 17488
rect 3753 17465 3787 17499
rect 3821 17465 3855 17499
rect 3889 17465 3923 17499
rect 3957 17465 3991 17499
rect 4025 17465 4059 17499
rect 4093 17465 4127 17499
rect 4161 17465 4195 17499
rect 5712 17466 5746 17500
rect 5780 17466 5814 17500
rect 5848 17466 5882 17500
rect 5916 17466 5950 17500
rect 5984 17466 6018 17500
rect 6052 17466 6086 17500
rect 6120 17466 6154 17500
rect 1353 16226 1387 16260
rect 1421 16226 1455 16260
rect 1489 16226 1523 16260
rect 1557 16226 1591 16260
rect 1625 16226 1659 16260
rect 1693 16226 1727 16260
rect 1761 16226 1795 16260
rect 1829 16226 1863 16260
rect 1897 16226 1931 16260
rect 3753 16237 3787 16271
rect 3821 16237 3855 16271
rect 3889 16237 3923 16271
rect 3957 16237 3991 16271
rect 4025 16237 4059 16271
rect 4093 16237 4127 16271
rect 4161 16237 4195 16271
rect 5712 16238 5746 16272
rect 5780 16238 5814 16272
rect 5848 16238 5882 16272
rect 5916 16238 5950 16272
rect 5984 16238 6018 16272
rect 6052 16238 6086 16272
rect 6120 16238 6154 16272
rect 1353 14998 1387 15032
rect 1421 14998 1455 15032
rect 1489 14998 1523 15032
rect 1557 14998 1591 15032
rect 1625 14998 1659 15032
rect 1693 14998 1727 15032
rect 1761 14998 1795 15032
rect 1829 14998 1863 15032
rect 1897 14998 1931 15032
rect 3753 15009 3787 15043
rect 3821 15009 3855 15043
rect 3889 15009 3923 15043
rect 3957 15009 3991 15043
rect 4025 15009 4059 15043
rect 4093 15009 4127 15043
rect 4161 15009 4195 15043
rect 5712 15010 5746 15044
rect 5780 15010 5814 15044
rect 5848 15010 5882 15044
rect 5916 15010 5950 15044
rect 5984 15010 6018 15044
rect 6052 15010 6086 15044
rect 6120 15010 6154 15044
rect 1353 13770 1387 13804
rect 1421 13770 1455 13804
rect 1489 13770 1523 13804
rect 1557 13770 1591 13804
rect 1625 13770 1659 13804
rect 1693 13770 1727 13804
rect 1761 13770 1795 13804
rect 1829 13770 1863 13804
rect 1897 13770 1931 13804
rect 3753 13781 3787 13815
rect 3821 13781 3855 13815
rect 3889 13781 3923 13815
rect 3957 13781 3991 13815
rect 4025 13781 4059 13815
rect 4093 13781 4127 13815
rect 4161 13781 4195 13815
rect 5712 13782 5746 13816
rect 5780 13782 5814 13816
rect 5848 13782 5882 13816
rect 5916 13782 5950 13816
rect 5984 13782 6018 13816
rect 6052 13782 6086 13816
rect 6120 13782 6154 13816
rect 1353 12542 1387 12576
rect 1421 12542 1455 12576
rect 1489 12542 1523 12576
rect 1557 12542 1591 12576
rect 1625 12542 1659 12576
rect 1693 12542 1727 12576
rect 1761 12542 1795 12576
rect 1829 12542 1863 12576
rect 1897 12542 1931 12576
rect 3753 12553 3787 12587
rect 3821 12553 3855 12587
rect 3889 12553 3923 12587
rect 3957 12553 3991 12587
rect 4025 12553 4059 12587
rect 4093 12553 4127 12587
rect 4161 12553 4195 12587
rect 5712 12554 5746 12588
rect 5780 12554 5814 12588
rect 5848 12554 5882 12588
rect 5916 12554 5950 12588
rect 5984 12554 6018 12588
rect 6052 12554 6086 12588
rect 6120 12554 6154 12588
rect 1353 11314 1387 11348
rect 1421 11314 1455 11348
rect 1489 11314 1523 11348
rect 1557 11314 1591 11348
rect 1625 11314 1659 11348
rect 1693 11314 1727 11348
rect 1761 11314 1795 11348
rect 1829 11314 1863 11348
rect 1897 11314 1931 11348
rect 3753 11325 3787 11359
rect 3821 11325 3855 11359
rect 3889 11325 3923 11359
rect 3957 11325 3991 11359
rect 4025 11325 4059 11359
rect 4093 11325 4127 11359
rect 4161 11325 4195 11359
rect 5712 11326 5746 11360
rect 5780 11326 5814 11360
rect 5848 11326 5882 11360
rect 5916 11326 5950 11360
rect 5984 11326 6018 11360
rect 6052 11326 6086 11360
rect 6120 11326 6154 11360
rect 1353 10086 1387 10120
rect 1421 10086 1455 10120
rect 1489 10086 1523 10120
rect 1557 10086 1591 10120
rect 1625 10086 1659 10120
rect 1693 10086 1727 10120
rect 1761 10086 1795 10120
rect 1829 10086 1863 10120
rect 1897 10086 1931 10120
rect 3753 10097 3787 10131
rect 3821 10097 3855 10131
rect 3889 10097 3923 10131
rect 3957 10097 3991 10131
rect 4025 10097 4059 10131
rect 4093 10097 4127 10131
rect 4161 10097 4195 10131
rect 5712 10098 5746 10132
rect 5780 10098 5814 10132
rect 5848 10098 5882 10132
rect 5916 10098 5950 10132
rect 5984 10098 6018 10132
rect 6052 10098 6086 10132
rect 6120 10098 6154 10132
rect 1353 8858 1387 8892
rect 1421 8858 1455 8892
rect 1489 8858 1523 8892
rect 1557 8858 1591 8892
rect 1625 8858 1659 8892
rect 1693 8858 1727 8892
rect 1761 8858 1795 8892
rect 1829 8858 1863 8892
rect 1897 8858 1931 8892
rect 3753 8869 3787 8903
rect 3821 8869 3855 8903
rect 3889 8869 3923 8903
rect 3957 8869 3991 8903
rect 4025 8869 4059 8903
rect 4093 8869 4127 8903
rect 4161 8869 4195 8903
rect 5712 8870 5746 8904
rect 5780 8870 5814 8904
rect 5848 8870 5882 8904
rect 5916 8870 5950 8904
rect 5984 8870 6018 8904
rect 6052 8870 6086 8904
rect 6120 8870 6154 8904
rect 1353 7630 1387 7664
rect 1421 7630 1455 7664
rect 1489 7630 1523 7664
rect 1557 7630 1591 7664
rect 1625 7630 1659 7664
rect 1693 7630 1727 7664
rect 1761 7630 1795 7664
rect 1829 7630 1863 7664
rect 1897 7630 1931 7664
rect 3753 7641 3787 7675
rect 3821 7641 3855 7675
rect 3889 7641 3923 7675
rect 3957 7641 3991 7675
rect 4025 7641 4059 7675
rect 4093 7641 4127 7675
rect 4161 7641 4195 7675
rect 5712 7642 5746 7676
rect 5780 7642 5814 7676
rect 5848 7642 5882 7676
rect 5916 7642 5950 7676
rect 5984 7642 6018 7676
rect 6052 7642 6086 7676
rect 6120 7642 6154 7676
rect 1353 6402 1387 6436
rect 1421 6402 1455 6436
rect 1489 6402 1523 6436
rect 1557 6402 1591 6436
rect 1625 6402 1659 6436
rect 1693 6402 1727 6436
rect 1761 6402 1795 6436
rect 1829 6402 1863 6436
rect 1897 6402 1931 6436
rect 3753 6413 3787 6447
rect 3821 6413 3855 6447
rect 3889 6413 3923 6447
rect 3957 6413 3991 6447
rect 4025 6413 4059 6447
rect 4093 6413 4127 6447
rect 4161 6413 4195 6447
rect 5712 6414 5746 6448
rect 5780 6414 5814 6448
rect 5848 6414 5882 6448
rect 5916 6414 5950 6448
rect 5984 6414 6018 6448
rect 6052 6414 6086 6448
rect 6120 6414 6154 6448
rect 1353 5174 1387 5208
rect 1421 5174 1455 5208
rect 1489 5174 1523 5208
rect 1557 5174 1591 5208
rect 1625 5174 1659 5208
rect 1693 5174 1727 5208
rect 1761 5174 1795 5208
rect 1829 5174 1863 5208
rect 1897 5174 1931 5208
rect 3753 5185 3787 5219
rect 3821 5185 3855 5219
rect 3889 5185 3923 5219
rect 3957 5185 3991 5219
rect 4025 5185 4059 5219
rect 4093 5185 4127 5219
rect 4161 5185 4195 5219
rect 5712 5186 5746 5220
rect 5780 5186 5814 5220
rect 5848 5186 5882 5220
rect 5916 5186 5950 5220
rect 5984 5186 6018 5220
rect 6052 5186 6086 5220
rect 6120 5186 6154 5220
rect 1353 3946 1387 3980
rect 1421 3946 1455 3980
rect 1489 3946 1523 3980
rect 1557 3946 1591 3980
rect 1625 3946 1659 3980
rect 1693 3946 1727 3980
rect 1761 3946 1795 3980
rect 1829 3946 1863 3980
rect 1897 3946 1931 3980
rect 3753 3957 3787 3991
rect 3821 3957 3855 3991
rect 3889 3957 3923 3991
rect 3957 3957 3991 3991
rect 4025 3957 4059 3991
rect 4093 3957 4127 3991
rect 4161 3957 4195 3991
rect 5712 3958 5746 3992
rect 5780 3958 5814 3992
rect 5848 3958 5882 3992
rect 5916 3958 5950 3992
rect 5984 3958 6018 3992
rect 6052 3958 6086 3992
rect 6120 3958 6154 3992
rect 1353 2718 1387 2752
rect 1421 2718 1455 2752
rect 1489 2718 1523 2752
rect 1557 2718 1591 2752
rect 1625 2718 1659 2752
rect 1693 2718 1727 2752
rect 1761 2718 1795 2752
rect 1829 2718 1863 2752
rect 1897 2718 1931 2752
rect 3753 2729 3787 2763
rect 3821 2729 3855 2763
rect 3889 2729 3923 2763
rect 3957 2729 3991 2763
rect 4025 2729 4059 2763
rect 4093 2729 4127 2763
rect 4161 2729 4195 2763
rect 5712 2730 5746 2764
rect 5780 2730 5814 2764
rect 5848 2730 5882 2764
rect 5916 2730 5950 2764
rect 5984 2730 6018 2764
rect 6052 2730 6086 2764
rect 6120 2730 6154 2764
rect 1353 1490 1387 1524
rect 1421 1490 1455 1524
rect 1489 1490 1523 1524
rect 1557 1490 1591 1524
rect 1625 1490 1659 1524
rect 1693 1490 1727 1524
rect 1761 1490 1795 1524
rect 1829 1490 1863 1524
rect 1897 1490 1931 1524
rect 3753 1501 3787 1535
rect 3821 1501 3855 1535
rect 3889 1501 3923 1535
rect 3957 1501 3991 1535
rect 4025 1501 4059 1535
rect 4093 1501 4127 1535
rect 4161 1501 4195 1535
rect 5712 1502 5746 1536
rect 5780 1502 5814 1536
rect 5848 1502 5882 1536
rect 5916 1502 5950 1536
rect 5984 1502 6018 1536
rect 6052 1502 6086 1536
rect 6120 1502 6154 1536
rect 1353 262 1387 296
rect 1421 262 1455 296
rect 1489 262 1523 296
rect 1557 262 1591 296
rect 1625 262 1659 296
rect 1693 262 1727 296
rect 1761 262 1795 296
rect 1829 262 1863 296
rect 1897 262 1931 296
rect 3753 273 3787 307
rect 3821 273 3855 307
rect 3889 273 3923 307
rect 3957 273 3991 307
rect 4025 273 4059 307
rect 4093 273 4127 307
rect 4161 273 4195 307
<< mvnsubdiffcont >>
rect 1395 19384 1429 19418
rect 1463 19384 1497 19418
rect 1531 19384 1565 19418
rect 1599 19384 1633 19418
rect 1667 19384 1701 19418
rect 1735 19384 1769 19418
rect 1803 19384 1837 19418
rect 3773 19383 3807 19417
rect 3841 19383 3875 19417
rect 3909 19383 3943 19417
rect 3977 19383 4011 19417
rect 4045 19383 4079 19417
rect 4113 19383 4147 19417
rect 4181 19383 4215 19417
rect 5732 19382 5766 19416
rect 5800 19382 5834 19416
rect 5868 19382 5902 19416
rect 5936 19382 5970 19416
rect 6004 19382 6038 19416
rect 6072 19382 6106 19416
rect 6140 19382 6174 19416
rect 1395 18156 1429 18190
rect 1463 18156 1497 18190
rect 1531 18156 1565 18190
rect 1599 18156 1633 18190
rect 1667 18156 1701 18190
rect 1735 18156 1769 18190
rect 1803 18156 1837 18190
rect 3773 18155 3807 18189
rect 3841 18155 3875 18189
rect 3909 18155 3943 18189
rect 3977 18155 4011 18189
rect 4045 18155 4079 18189
rect 4113 18155 4147 18189
rect 4181 18155 4215 18189
rect 5732 18154 5766 18188
rect 5800 18154 5834 18188
rect 5868 18154 5902 18188
rect 5936 18154 5970 18188
rect 6004 18154 6038 18188
rect 6072 18154 6106 18188
rect 6140 18154 6174 18188
rect 1395 16928 1429 16962
rect 1463 16928 1497 16962
rect 1531 16928 1565 16962
rect 1599 16928 1633 16962
rect 1667 16928 1701 16962
rect 1735 16928 1769 16962
rect 1803 16928 1837 16962
rect 3773 16927 3807 16961
rect 3841 16927 3875 16961
rect 3909 16927 3943 16961
rect 3977 16927 4011 16961
rect 4045 16927 4079 16961
rect 4113 16927 4147 16961
rect 4181 16927 4215 16961
rect 5732 16926 5766 16960
rect 5800 16926 5834 16960
rect 5868 16926 5902 16960
rect 5936 16926 5970 16960
rect 6004 16926 6038 16960
rect 6072 16926 6106 16960
rect 6140 16926 6174 16960
rect 1395 15700 1429 15734
rect 1463 15700 1497 15734
rect 1531 15700 1565 15734
rect 1599 15700 1633 15734
rect 1667 15700 1701 15734
rect 1735 15700 1769 15734
rect 1803 15700 1837 15734
rect 3773 15699 3807 15733
rect 3841 15699 3875 15733
rect 3909 15699 3943 15733
rect 3977 15699 4011 15733
rect 4045 15699 4079 15733
rect 4113 15699 4147 15733
rect 4181 15699 4215 15733
rect 5732 15698 5766 15732
rect 5800 15698 5834 15732
rect 5868 15698 5902 15732
rect 5936 15698 5970 15732
rect 6004 15698 6038 15732
rect 6072 15698 6106 15732
rect 6140 15698 6174 15732
rect 1395 14472 1429 14506
rect 1463 14472 1497 14506
rect 1531 14472 1565 14506
rect 1599 14472 1633 14506
rect 1667 14472 1701 14506
rect 1735 14472 1769 14506
rect 1803 14472 1837 14506
rect 3773 14471 3807 14505
rect 3841 14471 3875 14505
rect 3909 14471 3943 14505
rect 3977 14471 4011 14505
rect 4045 14471 4079 14505
rect 4113 14471 4147 14505
rect 4181 14471 4215 14505
rect 5732 14470 5766 14504
rect 5800 14470 5834 14504
rect 5868 14470 5902 14504
rect 5936 14470 5970 14504
rect 6004 14470 6038 14504
rect 6072 14470 6106 14504
rect 6140 14470 6174 14504
rect 1395 13244 1429 13278
rect 1463 13244 1497 13278
rect 1531 13244 1565 13278
rect 1599 13244 1633 13278
rect 1667 13244 1701 13278
rect 1735 13244 1769 13278
rect 1803 13244 1837 13278
rect 3773 13243 3807 13277
rect 3841 13243 3875 13277
rect 3909 13243 3943 13277
rect 3977 13243 4011 13277
rect 4045 13243 4079 13277
rect 4113 13243 4147 13277
rect 4181 13243 4215 13277
rect 5732 13242 5766 13276
rect 5800 13242 5834 13276
rect 5868 13242 5902 13276
rect 5936 13242 5970 13276
rect 6004 13242 6038 13276
rect 6072 13242 6106 13276
rect 6140 13242 6174 13276
rect 1395 12016 1429 12050
rect 1463 12016 1497 12050
rect 1531 12016 1565 12050
rect 1599 12016 1633 12050
rect 1667 12016 1701 12050
rect 1735 12016 1769 12050
rect 1803 12016 1837 12050
rect 3773 12015 3807 12049
rect 3841 12015 3875 12049
rect 3909 12015 3943 12049
rect 3977 12015 4011 12049
rect 4045 12015 4079 12049
rect 4113 12015 4147 12049
rect 4181 12015 4215 12049
rect 5732 12014 5766 12048
rect 5800 12014 5834 12048
rect 5868 12014 5902 12048
rect 5936 12014 5970 12048
rect 6004 12014 6038 12048
rect 6072 12014 6106 12048
rect 6140 12014 6174 12048
rect 1395 10788 1429 10822
rect 1463 10788 1497 10822
rect 1531 10788 1565 10822
rect 1599 10788 1633 10822
rect 1667 10788 1701 10822
rect 1735 10788 1769 10822
rect 1803 10788 1837 10822
rect 3773 10787 3807 10821
rect 3841 10787 3875 10821
rect 3909 10787 3943 10821
rect 3977 10787 4011 10821
rect 4045 10787 4079 10821
rect 4113 10787 4147 10821
rect 4181 10787 4215 10821
rect 5732 10786 5766 10820
rect 5800 10786 5834 10820
rect 5868 10786 5902 10820
rect 5936 10786 5970 10820
rect 6004 10786 6038 10820
rect 6072 10786 6106 10820
rect 6140 10786 6174 10820
rect 1395 9560 1429 9594
rect 1463 9560 1497 9594
rect 1531 9560 1565 9594
rect 1599 9560 1633 9594
rect 1667 9560 1701 9594
rect 1735 9560 1769 9594
rect 1803 9560 1837 9594
rect 3773 9559 3807 9593
rect 3841 9559 3875 9593
rect 3909 9559 3943 9593
rect 3977 9559 4011 9593
rect 4045 9559 4079 9593
rect 4113 9559 4147 9593
rect 4181 9559 4215 9593
rect 5732 9558 5766 9592
rect 5800 9558 5834 9592
rect 5868 9558 5902 9592
rect 5936 9558 5970 9592
rect 6004 9558 6038 9592
rect 6072 9558 6106 9592
rect 6140 9558 6174 9592
rect 1395 8332 1429 8366
rect 1463 8332 1497 8366
rect 1531 8332 1565 8366
rect 1599 8332 1633 8366
rect 1667 8332 1701 8366
rect 1735 8332 1769 8366
rect 1803 8332 1837 8366
rect 3773 8331 3807 8365
rect 3841 8331 3875 8365
rect 3909 8331 3943 8365
rect 3977 8331 4011 8365
rect 4045 8331 4079 8365
rect 4113 8331 4147 8365
rect 4181 8331 4215 8365
rect 5732 8330 5766 8364
rect 5800 8330 5834 8364
rect 5868 8330 5902 8364
rect 5936 8330 5970 8364
rect 6004 8330 6038 8364
rect 6072 8330 6106 8364
rect 6140 8330 6174 8364
rect 1395 7104 1429 7138
rect 1463 7104 1497 7138
rect 1531 7104 1565 7138
rect 1599 7104 1633 7138
rect 1667 7104 1701 7138
rect 1735 7104 1769 7138
rect 1803 7104 1837 7138
rect 3773 7103 3807 7137
rect 3841 7103 3875 7137
rect 3909 7103 3943 7137
rect 3977 7103 4011 7137
rect 4045 7103 4079 7137
rect 4113 7103 4147 7137
rect 4181 7103 4215 7137
rect 5732 7102 5766 7136
rect 5800 7102 5834 7136
rect 5868 7102 5902 7136
rect 5936 7102 5970 7136
rect 6004 7102 6038 7136
rect 6072 7102 6106 7136
rect 6140 7102 6174 7136
rect 1395 5876 1429 5910
rect 1463 5876 1497 5910
rect 1531 5876 1565 5910
rect 1599 5876 1633 5910
rect 1667 5876 1701 5910
rect 1735 5876 1769 5910
rect 1803 5876 1837 5910
rect 3773 5875 3807 5909
rect 3841 5875 3875 5909
rect 3909 5875 3943 5909
rect 3977 5875 4011 5909
rect 4045 5875 4079 5909
rect 4113 5875 4147 5909
rect 4181 5875 4215 5909
rect 5732 5874 5766 5908
rect 5800 5874 5834 5908
rect 5868 5874 5902 5908
rect 5936 5874 5970 5908
rect 6004 5874 6038 5908
rect 6072 5874 6106 5908
rect 6140 5874 6174 5908
rect 1395 4648 1429 4682
rect 1463 4648 1497 4682
rect 1531 4648 1565 4682
rect 1599 4648 1633 4682
rect 1667 4648 1701 4682
rect 1735 4648 1769 4682
rect 1803 4648 1837 4682
rect 3773 4647 3807 4681
rect 3841 4647 3875 4681
rect 3909 4647 3943 4681
rect 3977 4647 4011 4681
rect 4045 4647 4079 4681
rect 4113 4647 4147 4681
rect 4181 4647 4215 4681
rect 5732 4646 5766 4680
rect 5800 4646 5834 4680
rect 5868 4646 5902 4680
rect 5936 4646 5970 4680
rect 6004 4646 6038 4680
rect 6072 4646 6106 4680
rect 6140 4646 6174 4680
rect 1395 3420 1429 3454
rect 1463 3420 1497 3454
rect 1531 3420 1565 3454
rect 1599 3420 1633 3454
rect 1667 3420 1701 3454
rect 1735 3420 1769 3454
rect 1803 3420 1837 3454
rect 3773 3419 3807 3453
rect 3841 3419 3875 3453
rect 3909 3419 3943 3453
rect 3977 3419 4011 3453
rect 4045 3419 4079 3453
rect 4113 3419 4147 3453
rect 4181 3419 4215 3453
rect 5732 3418 5766 3452
rect 5800 3418 5834 3452
rect 5868 3418 5902 3452
rect 5936 3418 5970 3452
rect 6004 3418 6038 3452
rect 6072 3418 6106 3452
rect 6140 3418 6174 3452
rect 1395 2192 1429 2226
rect 1463 2192 1497 2226
rect 1531 2192 1565 2226
rect 1599 2192 1633 2226
rect 1667 2192 1701 2226
rect 1735 2192 1769 2226
rect 1803 2192 1837 2226
rect 3773 2191 3807 2225
rect 3841 2191 3875 2225
rect 3909 2191 3943 2225
rect 3977 2191 4011 2225
rect 4045 2191 4079 2225
rect 4113 2191 4147 2225
rect 4181 2191 4215 2225
rect 5732 2190 5766 2224
rect 5800 2190 5834 2224
rect 5868 2190 5902 2224
rect 5936 2190 5970 2224
rect 6004 2190 6038 2224
rect 6072 2190 6106 2224
rect 6140 2190 6174 2224
rect 1395 964 1429 998
rect 1463 964 1497 998
rect 1531 964 1565 998
rect 1599 964 1633 998
rect 1667 964 1701 998
rect 1735 964 1769 998
rect 1803 964 1837 998
rect 3773 963 3807 997
rect 3841 963 3875 997
rect 3909 963 3943 997
rect 3977 963 4011 997
rect 4045 963 4079 997
rect 4113 963 4147 997
rect 4181 963 4215 997
<< poly >>
rect 1456 19264 1556 19290
rect 1744 19264 1844 19290
rect 2076 19264 2176 19290
rect 2418 19264 2518 19290
rect 2822 19264 2922 19290
rect 3166 19264 3266 19290
rect 3788 19274 3888 19300
rect 4096 19274 4196 19300
rect 4448 19274 4548 19300
rect 4756 19274 4856 19300
rect 5746 19274 5846 19300
rect 6054 19274 6154 19300
rect 6406 19274 6506 19300
rect 6714 19274 6814 19300
rect 1456 19036 1556 19064
rect 1239 19011 1556 19036
rect 1239 18977 1269 19011
rect 1303 18977 1556 19011
rect 1239 18953 1556 18977
rect 1456 18926 1556 18953
rect 1744 19011 1844 19064
rect 1744 18977 1773 19011
rect 1807 18977 1844 19011
rect 1744 18926 1844 18977
rect 2076 19021 2176 19064
rect 2418 19042 2518 19064
rect 2621 19042 2707 19043
rect 2076 19009 2325 19021
rect 2076 18975 2273 19009
rect 2307 18975 2325 19009
rect 2076 18963 2325 18975
rect 2418 19019 2712 19042
rect 2418 18985 2647 19019
rect 2681 18985 2712 19019
rect 2076 18926 2176 18963
rect 2418 18951 2712 18985
rect 2822 19007 2922 19064
rect 2822 18973 2857 19007
rect 2891 18973 2922 19007
rect 2418 18926 2518 18951
rect 2822 18926 2922 18973
rect 3019 19017 3073 19023
rect 3166 19017 3266 19064
rect 3019 19007 3266 19017
rect 3019 18973 3029 19007
rect 3063 18973 3266 19007
rect 3654 19033 3720 19041
rect 3788 19033 3888 19074
rect 3654 19031 3888 19033
rect 3654 18997 3670 19031
rect 3704 18997 3888 19031
rect 3654 18994 3888 18997
rect 3654 18987 3720 18994
rect 3019 18963 3266 18973
rect 3019 18957 3073 18963
rect 3166 18926 3266 18963
rect 3788 18936 3888 18994
rect 3968 19024 4034 19032
rect 4096 19024 4196 19074
rect 3968 19022 4196 19024
rect 3968 18988 3984 19022
rect 4018 18988 4196 19022
rect 3968 18985 4196 18988
rect 3968 18978 4034 18985
rect 4096 18936 4196 18985
rect 4290 19016 4356 19026
rect 4448 19016 4548 19074
rect 4290 18982 4306 19016
rect 4340 18982 4548 19016
rect 4627 19034 4681 19050
rect 4627 19000 4637 19034
rect 4671 19032 4681 19034
rect 4756 19032 4856 19074
rect 4671 19001 4856 19032
rect 4671 19000 4681 19001
rect 4627 18984 4681 19000
rect 4290 18981 4548 18982
rect 4290 18972 4356 18981
rect 4448 18938 4548 18981
rect 4756 18938 4856 19001
rect 5612 19034 5678 19042
rect 5746 19034 5846 19074
rect 5612 19032 5846 19034
rect 5612 18998 5628 19032
rect 5662 18998 5846 19032
rect 5612 18994 5846 18998
rect 5612 18988 5678 18994
rect 5746 18936 5846 18994
rect 5926 19024 5992 19032
rect 6054 19024 6154 19074
rect 5926 19022 6154 19024
rect 5926 18988 5942 19022
rect 5976 18988 6154 19022
rect 5926 18986 6154 18988
rect 5926 18978 5992 18986
rect 6054 18936 6154 18986
rect 6248 19016 6314 19026
rect 6406 19016 6506 19074
rect 6248 18982 6264 19016
rect 6298 18982 6506 19016
rect 6586 19034 6640 19050
rect 6586 19000 6596 19034
rect 6630 19032 6640 19034
rect 6714 19032 6814 19074
rect 6630 19002 6814 19032
rect 6630 19000 6640 19002
rect 6586 18984 6640 19000
rect 6248 18972 6314 18982
rect 6406 18938 6506 18982
rect 6714 18938 6814 19002
rect 1456 18800 1556 18826
rect 1744 18800 1844 18826
rect 2076 18800 2176 18826
rect 2418 18800 2518 18826
rect 2822 18800 2922 18826
rect 3166 18800 3266 18826
rect 3788 18810 3888 18836
rect 4096 18810 4196 18836
rect 4448 18812 4548 18838
rect 4756 18812 4856 18838
rect 5746 18810 5846 18836
rect 6054 18810 6154 18836
rect 6406 18812 6506 18838
rect 6714 18812 6814 18838
rect 1456 18036 1556 18062
rect 1744 18036 1844 18062
rect 2076 18036 2176 18062
rect 2418 18036 2518 18062
rect 2822 18036 2922 18062
rect 3166 18036 3266 18062
rect 3788 18046 3888 18072
rect 4096 18046 4196 18072
rect 4448 18046 4548 18072
rect 4756 18046 4856 18072
rect 5746 18046 5846 18072
rect 6054 18046 6154 18072
rect 6406 18046 6506 18072
rect 6714 18046 6814 18072
rect 1456 17808 1556 17836
rect 1239 17783 1556 17808
rect 1239 17749 1269 17783
rect 1303 17749 1556 17783
rect 1239 17725 1556 17749
rect 1456 17698 1556 17725
rect 1744 17783 1844 17836
rect 1744 17749 1773 17783
rect 1807 17749 1844 17783
rect 1744 17698 1844 17749
rect 2076 17793 2176 17836
rect 2418 17814 2518 17836
rect 2621 17814 2707 17815
rect 2076 17781 2325 17793
rect 2076 17747 2273 17781
rect 2307 17747 2325 17781
rect 2076 17735 2325 17747
rect 2418 17791 2712 17814
rect 2418 17757 2647 17791
rect 2681 17757 2712 17791
rect 2076 17698 2176 17735
rect 2418 17723 2712 17757
rect 2822 17779 2922 17836
rect 2822 17745 2857 17779
rect 2891 17745 2922 17779
rect 2418 17698 2518 17723
rect 2822 17698 2922 17745
rect 3019 17789 3073 17795
rect 3166 17789 3266 17836
rect 3019 17779 3266 17789
rect 3019 17745 3029 17779
rect 3063 17745 3266 17779
rect 3654 17805 3720 17813
rect 3788 17805 3888 17846
rect 3654 17803 3888 17805
rect 3654 17769 3670 17803
rect 3704 17769 3888 17803
rect 3654 17766 3888 17769
rect 3654 17759 3720 17766
rect 3019 17735 3266 17745
rect 3019 17729 3073 17735
rect 3166 17698 3266 17735
rect 3788 17708 3888 17766
rect 3968 17796 4034 17804
rect 4096 17796 4196 17846
rect 3968 17794 4196 17796
rect 3968 17760 3984 17794
rect 4018 17760 4196 17794
rect 3968 17757 4196 17760
rect 3968 17750 4034 17757
rect 4096 17708 4196 17757
rect 4290 17788 4356 17798
rect 4448 17788 4548 17846
rect 4290 17754 4306 17788
rect 4340 17754 4548 17788
rect 4627 17806 4681 17822
rect 4627 17772 4637 17806
rect 4671 17804 4681 17806
rect 4756 17804 4856 17846
rect 4671 17773 4856 17804
rect 4671 17772 4681 17773
rect 4627 17756 4681 17772
rect 4290 17753 4548 17754
rect 4290 17744 4356 17753
rect 4448 17710 4548 17753
rect 4756 17710 4856 17773
rect 5612 17806 5678 17814
rect 5746 17806 5846 17846
rect 5612 17804 5846 17806
rect 5612 17770 5628 17804
rect 5662 17770 5846 17804
rect 5612 17766 5846 17770
rect 5612 17760 5678 17766
rect 5746 17708 5846 17766
rect 5926 17796 5992 17804
rect 6054 17796 6154 17846
rect 5926 17794 6154 17796
rect 5926 17760 5942 17794
rect 5976 17760 6154 17794
rect 5926 17758 6154 17760
rect 5926 17750 5992 17758
rect 6054 17708 6154 17758
rect 6248 17788 6314 17798
rect 6406 17788 6506 17846
rect 6248 17754 6264 17788
rect 6298 17754 6506 17788
rect 6586 17806 6640 17822
rect 6586 17772 6596 17806
rect 6630 17804 6640 17806
rect 6714 17804 6814 17846
rect 6630 17774 6814 17804
rect 6630 17772 6640 17774
rect 6586 17756 6640 17772
rect 6248 17744 6314 17754
rect 6406 17710 6506 17754
rect 6714 17710 6814 17774
rect 1456 17572 1556 17598
rect 1744 17572 1844 17598
rect 2076 17572 2176 17598
rect 2418 17572 2518 17598
rect 2822 17572 2922 17598
rect 3166 17572 3266 17598
rect 3788 17582 3888 17608
rect 4096 17582 4196 17608
rect 4448 17584 4548 17610
rect 4756 17584 4856 17610
rect 5746 17582 5846 17608
rect 6054 17582 6154 17608
rect 6406 17584 6506 17610
rect 6714 17584 6814 17610
rect 1456 16808 1556 16834
rect 1744 16808 1844 16834
rect 2076 16808 2176 16834
rect 2418 16808 2518 16834
rect 2822 16808 2922 16834
rect 3166 16808 3266 16834
rect 3788 16818 3888 16844
rect 4096 16818 4196 16844
rect 4448 16818 4548 16844
rect 4756 16818 4856 16844
rect 5746 16818 5846 16844
rect 6054 16818 6154 16844
rect 6406 16818 6506 16844
rect 6714 16818 6814 16844
rect 1456 16580 1556 16608
rect 1239 16555 1556 16580
rect 1239 16521 1269 16555
rect 1303 16521 1556 16555
rect 1239 16497 1556 16521
rect 1456 16470 1556 16497
rect 1744 16555 1844 16608
rect 1744 16521 1773 16555
rect 1807 16521 1844 16555
rect 1744 16470 1844 16521
rect 2076 16565 2176 16608
rect 2418 16586 2518 16608
rect 2621 16586 2707 16587
rect 2076 16553 2325 16565
rect 2076 16519 2273 16553
rect 2307 16519 2325 16553
rect 2076 16507 2325 16519
rect 2418 16563 2712 16586
rect 2418 16529 2647 16563
rect 2681 16529 2712 16563
rect 2076 16470 2176 16507
rect 2418 16495 2712 16529
rect 2822 16551 2922 16608
rect 2822 16517 2857 16551
rect 2891 16517 2922 16551
rect 2418 16470 2518 16495
rect 2822 16470 2922 16517
rect 3019 16561 3073 16567
rect 3166 16561 3266 16608
rect 3019 16551 3266 16561
rect 3019 16517 3029 16551
rect 3063 16517 3266 16551
rect 3654 16577 3720 16585
rect 3788 16577 3888 16618
rect 3654 16575 3888 16577
rect 3654 16541 3670 16575
rect 3704 16541 3888 16575
rect 3654 16538 3888 16541
rect 3654 16531 3720 16538
rect 3019 16507 3266 16517
rect 3019 16501 3073 16507
rect 3166 16470 3266 16507
rect 3788 16480 3888 16538
rect 3968 16568 4034 16576
rect 4096 16568 4196 16618
rect 3968 16566 4196 16568
rect 3968 16532 3984 16566
rect 4018 16532 4196 16566
rect 3968 16529 4196 16532
rect 3968 16522 4034 16529
rect 4096 16480 4196 16529
rect 4290 16560 4356 16570
rect 4448 16560 4548 16618
rect 4290 16526 4306 16560
rect 4340 16526 4548 16560
rect 4627 16578 4681 16594
rect 4627 16544 4637 16578
rect 4671 16576 4681 16578
rect 4756 16576 4856 16618
rect 4671 16545 4856 16576
rect 4671 16544 4681 16545
rect 4627 16528 4681 16544
rect 4290 16525 4548 16526
rect 4290 16516 4356 16525
rect 4448 16482 4548 16525
rect 4756 16482 4856 16545
rect 5612 16578 5678 16586
rect 5746 16578 5846 16618
rect 5612 16576 5846 16578
rect 5612 16542 5628 16576
rect 5662 16542 5846 16576
rect 5612 16538 5846 16542
rect 5612 16532 5678 16538
rect 5746 16480 5846 16538
rect 5926 16568 5992 16576
rect 6054 16568 6154 16618
rect 5926 16566 6154 16568
rect 5926 16532 5942 16566
rect 5976 16532 6154 16566
rect 5926 16530 6154 16532
rect 5926 16522 5992 16530
rect 6054 16480 6154 16530
rect 6248 16560 6314 16570
rect 6406 16560 6506 16618
rect 6248 16526 6264 16560
rect 6298 16526 6506 16560
rect 6586 16578 6640 16594
rect 6586 16544 6596 16578
rect 6630 16576 6640 16578
rect 6714 16576 6814 16618
rect 6630 16546 6814 16576
rect 6630 16544 6640 16546
rect 6586 16528 6640 16544
rect 6248 16516 6314 16526
rect 6406 16482 6506 16526
rect 6714 16482 6814 16546
rect 1456 16344 1556 16370
rect 1744 16344 1844 16370
rect 2076 16344 2176 16370
rect 2418 16344 2518 16370
rect 2822 16344 2922 16370
rect 3166 16344 3266 16370
rect 3788 16354 3888 16380
rect 4096 16354 4196 16380
rect 4448 16356 4548 16382
rect 4756 16356 4856 16382
rect 5746 16354 5846 16380
rect 6054 16354 6154 16380
rect 6406 16356 6506 16382
rect 6714 16356 6814 16382
rect 1456 15580 1556 15606
rect 1744 15580 1844 15606
rect 2076 15580 2176 15606
rect 2418 15580 2518 15606
rect 2822 15580 2922 15606
rect 3166 15580 3266 15606
rect 3788 15590 3888 15616
rect 4096 15590 4196 15616
rect 4448 15590 4548 15616
rect 4756 15590 4856 15616
rect 5746 15590 5846 15616
rect 6054 15590 6154 15616
rect 6406 15590 6506 15616
rect 6714 15590 6814 15616
rect 1456 15352 1556 15380
rect 1239 15327 1556 15352
rect 1239 15293 1269 15327
rect 1303 15293 1556 15327
rect 1239 15269 1556 15293
rect 1456 15242 1556 15269
rect 1744 15327 1844 15380
rect 1744 15293 1773 15327
rect 1807 15293 1844 15327
rect 1744 15242 1844 15293
rect 2076 15337 2176 15380
rect 2418 15358 2518 15380
rect 2621 15358 2707 15359
rect 2076 15325 2325 15337
rect 2076 15291 2273 15325
rect 2307 15291 2325 15325
rect 2076 15279 2325 15291
rect 2418 15335 2712 15358
rect 2418 15301 2647 15335
rect 2681 15301 2712 15335
rect 2076 15242 2176 15279
rect 2418 15267 2712 15301
rect 2822 15323 2922 15380
rect 2822 15289 2857 15323
rect 2891 15289 2922 15323
rect 2418 15242 2518 15267
rect 2822 15242 2922 15289
rect 3019 15333 3073 15339
rect 3166 15333 3266 15380
rect 3019 15323 3266 15333
rect 3019 15289 3029 15323
rect 3063 15289 3266 15323
rect 3654 15349 3720 15357
rect 3788 15349 3888 15390
rect 3654 15347 3888 15349
rect 3654 15313 3670 15347
rect 3704 15313 3888 15347
rect 3654 15310 3888 15313
rect 3654 15303 3720 15310
rect 3019 15279 3266 15289
rect 3019 15273 3073 15279
rect 3166 15242 3266 15279
rect 3788 15252 3888 15310
rect 3968 15340 4034 15348
rect 4096 15340 4196 15390
rect 3968 15338 4196 15340
rect 3968 15304 3984 15338
rect 4018 15304 4196 15338
rect 3968 15301 4196 15304
rect 3968 15294 4034 15301
rect 4096 15252 4196 15301
rect 4290 15332 4356 15342
rect 4448 15332 4548 15390
rect 4290 15298 4306 15332
rect 4340 15298 4548 15332
rect 4627 15350 4681 15366
rect 4627 15316 4637 15350
rect 4671 15348 4681 15350
rect 4756 15348 4856 15390
rect 4671 15317 4856 15348
rect 4671 15316 4681 15317
rect 4627 15300 4681 15316
rect 4290 15297 4548 15298
rect 4290 15288 4356 15297
rect 4448 15254 4548 15297
rect 4756 15254 4856 15317
rect 5612 15350 5678 15358
rect 5746 15350 5846 15390
rect 5612 15348 5846 15350
rect 5612 15314 5628 15348
rect 5662 15314 5846 15348
rect 5612 15310 5846 15314
rect 5612 15304 5678 15310
rect 5746 15252 5846 15310
rect 5926 15340 5992 15348
rect 6054 15340 6154 15390
rect 5926 15338 6154 15340
rect 5926 15304 5942 15338
rect 5976 15304 6154 15338
rect 5926 15302 6154 15304
rect 5926 15294 5992 15302
rect 6054 15252 6154 15302
rect 6248 15332 6314 15342
rect 6406 15332 6506 15390
rect 6248 15298 6264 15332
rect 6298 15298 6506 15332
rect 6586 15350 6640 15366
rect 6586 15316 6596 15350
rect 6630 15348 6640 15350
rect 6714 15348 6814 15390
rect 6630 15318 6814 15348
rect 6630 15316 6640 15318
rect 6586 15300 6640 15316
rect 6248 15288 6314 15298
rect 6406 15254 6506 15298
rect 6714 15254 6814 15318
rect 1456 15116 1556 15142
rect 1744 15116 1844 15142
rect 2076 15116 2176 15142
rect 2418 15116 2518 15142
rect 2822 15116 2922 15142
rect 3166 15116 3266 15142
rect 3788 15126 3888 15152
rect 4096 15126 4196 15152
rect 4448 15128 4548 15154
rect 4756 15128 4856 15154
rect 5746 15126 5846 15152
rect 6054 15126 6154 15152
rect 6406 15128 6506 15154
rect 6714 15128 6814 15154
rect 1456 14352 1556 14378
rect 1744 14352 1844 14378
rect 2076 14352 2176 14378
rect 2418 14352 2518 14378
rect 2822 14352 2922 14378
rect 3166 14352 3266 14378
rect 3788 14362 3888 14388
rect 4096 14362 4196 14388
rect 4448 14362 4548 14388
rect 4756 14362 4856 14388
rect 5746 14362 5846 14388
rect 6054 14362 6154 14388
rect 6406 14362 6506 14388
rect 6714 14362 6814 14388
rect 1456 14124 1556 14152
rect 1239 14099 1556 14124
rect 1239 14065 1269 14099
rect 1303 14065 1556 14099
rect 1239 14041 1556 14065
rect 1456 14014 1556 14041
rect 1744 14099 1844 14152
rect 1744 14065 1773 14099
rect 1807 14065 1844 14099
rect 1744 14014 1844 14065
rect 2076 14109 2176 14152
rect 2418 14130 2518 14152
rect 2621 14130 2707 14131
rect 2076 14097 2325 14109
rect 2076 14063 2273 14097
rect 2307 14063 2325 14097
rect 2076 14051 2325 14063
rect 2418 14107 2712 14130
rect 2418 14073 2647 14107
rect 2681 14073 2712 14107
rect 2076 14014 2176 14051
rect 2418 14039 2712 14073
rect 2822 14095 2922 14152
rect 2822 14061 2857 14095
rect 2891 14061 2922 14095
rect 2418 14014 2518 14039
rect 2822 14014 2922 14061
rect 3019 14105 3073 14111
rect 3166 14105 3266 14152
rect 3019 14095 3266 14105
rect 3019 14061 3029 14095
rect 3063 14061 3266 14095
rect 3654 14121 3720 14129
rect 3788 14121 3888 14162
rect 3654 14119 3888 14121
rect 3654 14085 3670 14119
rect 3704 14085 3888 14119
rect 3654 14082 3888 14085
rect 3654 14075 3720 14082
rect 3019 14051 3266 14061
rect 3019 14045 3073 14051
rect 3166 14014 3266 14051
rect 3788 14024 3888 14082
rect 3968 14112 4034 14120
rect 4096 14112 4196 14162
rect 3968 14110 4196 14112
rect 3968 14076 3984 14110
rect 4018 14076 4196 14110
rect 3968 14073 4196 14076
rect 3968 14066 4034 14073
rect 4096 14024 4196 14073
rect 4290 14104 4356 14114
rect 4448 14104 4548 14162
rect 4290 14070 4306 14104
rect 4340 14070 4548 14104
rect 4627 14122 4681 14138
rect 4627 14088 4637 14122
rect 4671 14120 4681 14122
rect 4756 14120 4856 14162
rect 4671 14089 4856 14120
rect 4671 14088 4681 14089
rect 4627 14072 4681 14088
rect 4290 14069 4548 14070
rect 4290 14060 4356 14069
rect 4448 14026 4548 14069
rect 4756 14026 4856 14089
rect 5612 14122 5678 14130
rect 5746 14122 5846 14162
rect 5612 14120 5846 14122
rect 5612 14086 5628 14120
rect 5662 14086 5846 14120
rect 5612 14082 5846 14086
rect 5612 14076 5678 14082
rect 5746 14024 5846 14082
rect 5926 14112 5992 14120
rect 6054 14112 6154 14162
rect 5926 14110 6154 14112
rect 5926 14076 5942 14110
rect 5976 14076 6154 14110
rect 5926 14074 6154 14076
rect 5926 14066 5992 14074
rect 6054 14024 6154 14074
rect 6248 14104 6314 14114
rect 6406 14104 6506 14162
rect 6248 14070 6264 14104
rect 6298 14070 6506 14104
rect 6586 14122 6640 14138
rect 6586 14088 6596 14122
rect 6630 14120 6640 14122
rect 6714 14120 6814 14162
rect 6630 14090 6814 14120
rect 6630 14088 6640 14090
rect 6586 14072 6640 14088
rect 6248 14060 6314 14070
rect 6406 14026 6506 14070
rect 6714 14026 6814 14090
rect 1456 13888 1556 13914
rect 1744 13888 1844 13914
rect 2076 13888 2176 13914
rect 2418 13888 2518 13914
rect 2822 13888 2922 13914
rect 3166 13888 3266 13914
rect 3788 13898 3888 13924
rect 4096 13898 4196 13924
rect 4448 13900 4548 13926
rect 4756 13900 4856 13926
rect 5746 13898 5846 13924
rect 6054 13898 6154 13924
rect 6406 13900 6506 13926
rect 6714 13900 6814 13926
rect 1456 13124 1556 13150
rect 1744 13124 1844 13150
rect 2076 13124 2176 13150
rect 2418 13124 2518 13150
rect 2822 13124 2922 13150
rect 3166 13124 3266 13150
rect 3788 13134 3888 13160
rect 4096 13134 4196 13160
rect 4448 13134 4548 13160
rect 4756 13134 4856 13160
rect 5746 13134 5846 13160
rect 6054 13134 6154 13160
rect 6406 13134 6506 13160
rect 6714 13134 6814 13160
rect 1456 12896 1556 12924
rect 1239 12871 1556 12896
rect 1239 12837 1269 12871
rect 1303 12837 1556 12871
rect 1239 12813 1556 12837
rect 1456 12786 1556 12813
rect 1744 12871 1844 12924
rect 1744 12837 1773 12871
rect 1807 12837 1844 12871
rect 1744 12786 1844 12837
rect 2076 12881 2176 12924
rect 2418 12902 2518 12924
rect 2621 12902 2707 12903
rect 2076 12869 2325 12881
rect 2076 12835 2273 12869
rect 2307 12835 2325 12869
rect 2076 12823 2325 12835
rect 2418 12879 2712 12902
rect 2418 12845 2647 12879
rect 2681 12845 2712 12879
rect 2076 12786 2176 12823
rect 2418 12811 2712 12845
rect 2822 12867 2922 12924
rect 2822 12833 2857 12867
rect 2891 12833 2922 12867
rect 2418 12786 2518 12811
rect 2822 12786 2922 12833
rect 3019 12877 3073 12883
rect 3166 12877 3266 12924
rect 3019 12867 3266 12877
rect 3019 12833 3029 12867
rect 3063 12833 3266 12867
rect 3654 12893 3720 12901
rect 3788 12893 3888 12934
rect 3654 12891 3888 12893
rect 3654 12857 3670 12891
rect 3704 12857 3888 12891
rect 3654 12854 3888 12857
rect 3654 12847 3720 12854
rect 3019 12823 3266 12833
rect 3019 12817 3073 12823
rect 3166 12786 3266 12823
rect 3788 12796 3888 12854
rect 3968 12884 4034 12892
rect 4096 12884 4196 12934
rect 3968 12882 4196 12884
rect 3968 12848 3984 12882
rect 4018 12848 4196 12882
rect 3968 12845 4196 12848
rect 3968 12838 4034 12845
rect 4096 12796 4196 12845
rect 4290 12876 4356 12886
rect 4448 12876 4548 12934
rect 4290 12842 4306 12876
rect 4340 12842 4548 12876
rect 4627 12894 4681 12910
rect 4627 12860 4637 12894
rect 4671 12892 4681 12894
rect 4756 12892 4856 12934
rect 4671 12861 4856 12892
rect 4671 12860 4681 12861
rect 4627 12844 4681 12860
rect 4290 12841 4548 12842
rect 4290 12832 4356 12841
rect 4448 12798 4548 12841
rect 4756 12798 4856 12861
rect 5612 12894 5678 12902
rect 5746 12894 5846 12934
rect 5612 12892 5846 12894
rect 5612 12858 5628 12892
rect 5662 12858 5846 12892
rect 5612 12854 5846 12858
rect 5612 12848 5678 12854
rect 5746 12796 5846 12854
rect 5926 12884 5992 12892
rect 6054 12884 6154 12934
rect 5926 12882 6154 12884
rect 5926 12848 5942 12882
rect 5976 12848 6154 12882
rect 5926 12846 6154 12848
rect 5926 12838 5992 12846
rect 6054 12796 6154 12846
rect 6248 12876 6314 12886
rect 6406 12876 6506 12934
rect 6248 12842 6264 12876
rect 6298 12842 6506 12876
rect 6586 12894 6640 12910
rect 6586 12860 6596 12894
rect 6630 12892 6640 12894
rect 6714 12892 6814 12934
rect 6630 12862 6814 12892
rect 6630 12860 6640 12862
rect 6586 12844 6640 12860
rect 6248 12832 6314 12842
rect 6406 12798 6506 12842
rect 6714 12798 6814 12862
rect 1456 12660 1556 12686
rect 1744 12660 1844 12686
rect 2076 12660 2176 12686
rect 2418 12660 2518 12686
rect 2822 12660 2922 12686
rect 3166 12660 3266 12686
rect 3788 12670 3888 12696
rect 4096 12670 4196 12696
rect 4448 12672 4548 12698
rect 4756 12672 4856 12698
rect 5746 12670 5846 12696
rect 6054 12670 6154 12696
rect 6406 12672 6506 12698
rect 6714 12672 6814 12698
rect 1456 11896 1556 11922
rect 1744 11896 1844 11922
rect 2076 11896 2176 11922
rect 2418 11896 2518 11922
rect 2822 11896 2922 11922
rect 3166 11896 3266 11922
rect 3788 11906 3888 11932
rect 4096 11906 4196 11932
rect 4448 11906 4548 11932
rect 4756 11906 4856 11932
rect 5746 11906 5846 11932
rect 6054 11906 6154 11932
rect 6406 11906 6506 11932
rect 6714 11906 6814 11932
rect 1456 11668 1556 11696
rect 1239 11643 1556 11668
rect 1239 11609 1269 11643
rect 1303 11609 1556 11643
rect 1239 11585 1556 11609
rect 1456 11558 1556 11585
rect 1744 11643 1844 11696
rect 1744 11609 1773 11643
rect 1807 11609 1844 11643
rect 1744 11558 1844 11609
rect 2076 11653 2176 11696
rect 2418 11674 2518 11696
rect 2621 11674 2707 11675
rect 2076 11641 2325 11653
rect 2076 11607 2273 11641
rect 2307 11607 2325 11641
rect 2076 11595 2325 11607
rect 2418 11651 2712 11674
rect 2418 11617 2647 11651
rect 2681 11617 2712 11651
rect 2076 11558 2176 11595
rect 2418 11583 2712 11617
rect 2822 11639 2922 11696
rect 2822 11605 2857 11639
rect 2891 11605 2922 11639
rect 2418 11558 2518 11583
rect 2822 11558 2922 11605
rect 3019 11649 3073 11655
rect 3166 11649 3266 11696
rect 3019 11639 3266 11649
rect 3019 11605 3029 11639
rect 3063 11605 3266 11639
rect 3654 11665 3720 11673
rect 3788 11665 3888 11706
rect 3654 11663 3888 11665
rect 3654 11629 3670 11663
rect 3704 11629 3888 11663
rect 3654 11626 3888 11629
rect 3654 11619 3720 11626
rect 3019 11595 3266 11605
rect 3019 11589 3073 11595
rect 3166 11558 3266 11595
rect 3788 11568 3888 11626
rect 3968 11656 4034 11664
rect 4096 11656 4196 11706
rect 3968 11654 4196 11656
rect 3968 11620 3984 11654
rect 4018 11620 4196 11654
rect 3968 11617 4196 11620
rect 3968 11610 4034 11617
rect 4096 11568 4196 11617
rect 4290 11648 4356 11658
rect 4448 11648 4548 11706
rect 4290 11614 4306 11648
rect 4340 11614 4548 11648
rect 4627 11666 4681 11682
rect 4627 11632 4637 11666
rect 4671 11664 4681 11666
rect 4756 11664 4856 11706
rect 4671 11633 4856 11664
rect 4671 11632 4681 11633
rect 4627 11616 4681 11632
rect 4290 11613 4548 11614
rect 4290 11604 4356 11613
rect 4448 11570 4548 11613
rect 4756 11570 4856 11633
rect 5612 11666 5678 11674
rect 5746 11666 5846 11706
rect 5612 11664 5846 11666
rect 5612 11630 5628 11664
rect 5662 11630 5846 11664
rect 5612 11626 5846 11630
rect 5612 11620 5678 11626
rect 5746 11568 5846 11626
rect 5926 11656 5992 11664
rect 6054 11656 6154 11706
rect 5926 11654 6154 11656
rect 5926 11620 5942 11654
rect 5976 11620 6154 11654
rect 5926 11618 6154 11620
rect 5926 11610 5992 11618
rect 6054 11568 6154 11618
rect 6248 11648 6314 11658
rect 6406 11648 6506 11706
rect 6248 11614 6264 11648
rect 6298 11614 6506 11648
rect 6586 11666 6640 11682
rect 6586 11632 6596 11666
rect 6630 11664 6640 11666
rect 6714 11664 6814 11706
rect 6630 11634 6814 11664
rect 6630 11632 6640 11634
rect 6586 11616 6640 11632
rect 6248 11604 6314 11614
rect 6406 11570 6506 11614
rect 6714 11570 6814 11634
rect 1456 11432 1556 11458
rect 1744 11432 1844 11458
rect 2076 11432 2176 11458
rect 2418 11432 2518 11458
rect 2822 11432 2922 11458
rect 3166 11432 3266 11458
rect 3788 11442 3888 11468
rect 4096 11442 4196 11468
rect 4448 11444 4548 11470
rect 4756 11444 4856 11470
rect 5746 11442 5846 11468
rect 6054 11442 6154 11468
rect 6406 11444 6506 11470
rect 6714 11444 6814 11470
rect 1456 10668 1556 10694
rect 1744 10668 1844 10694
rect 2076 10668 2176 10694
rect 2418 10668 2518 10694
rect 2822 10668 2922 10694
rect 3166 10668 3266 10694
rect 3788 10678 3888 10704
rect 4096 10678 4196 10704
rect 4448 10678 4548 10704
rect 4756 10678 4856 10704
rect 5746 10678 5846 10704
rect 6054 10678 6154 10704
rect 6406 10678 6506 10704
rect 6714 10678 6814 10704
rect 1456 10440 1556 10468
rect 1239 10415 1556 10440
rect 1239 10381 1269 10415
rect 1303 10381 1556 10415
rect 1239 10357 1556 10381
rect 1456 10330 1556 10357
rect 1744 10415 1844 10468
rect 1744 10381 1773 10415
rect 1807 10381 1844 10415
rect 1744 10330 1844 10381
rect 2076 10425 2176 10468
rect 2418 10446 2518 10468
rect 2621 10446 2707 10447
rect 2076 10413 2325 10425
rect 2076 10379 2273 10413
rect 2307 10379 2325 10413
rect 2076 10367 2325 10379
rect 2418 10423 2712 10446
rect 2418 10389 2647 10423
rect 2681 10389 2712 10423
rect 2076 10330 2176 10367
rect 2418 10355 2712 10389
rect 2822 10411 2922 10468
rect 2822 10377 2857 10411
rect 2891 10377 2922 10411
rect 2418 10330 2518 10355
rect 2822 10330 2922 10377
rect 3019 10421 3073 10427
rect 3166 10421 3266 10468
rect 3019 10411 3266 10421
rect 3019 10377 3029 10411
rect 3063 10377 3266 10411
rect 3654 10437 3720 10445
rect 3788 10437 3888 10478
rect 3654 10435 3888 10437
rect 3654 10401 3670 10435
rect 3704 10401 3888 10435
rect 3654 10398 3888 10401
rect 3654 10391 3720 10398
rect 3019 10367 3266 10377
rect 3019 10361 3073 10367
rect 3166 10330 3266 10367
rect 3788 10340 3888 10398
rect 3968 10428 4034 10436
rect 4096 10428 4196 10478
rect 3968 10426 4196 10428
rect 3968 10392 3984 10426
rect 4018 10392 4196 10426
rect 3968 10389 4196 10392
rect 3968 10382 4034 10389
rect 4096 10340 4196 10389
rect 4290 10420 4356 10430
rect 4448 10420 4548 10478
rect 4290 10386 4306 10420
rect 4340 10386 4548 10420
rect 4627 10438 4681 10454
rect 4627 10404 4637 10438
rect 4671 10436 4681 10438
rect 4756 10436 4856 10478
rect 4671 10405 4856 10436
rect 4671 10404 4681 10405
rect 4627 10388 4681 10404
rect 4290 10385 4548 10386
rect 4290 10376 4356 10385
rect 4448 10342 4548 10385
rect 4756 10342 4856 10405
rect 5612 10438 5678 10446
rect 5746 10438 5846 10478
rect 5612 10436 5846 10438
rect 5612 10402 5628 10436
rect 5662 10402 5846 10436
rect 5612 10398 5846 10402
rect 5612 10392 5678 10398
rect 5746 10340 5846 10398
rect 5926 10428 5992 10436
rect 6054 10428 6154 10478
rect 5926 10426 6154 10428
rect 5926 10392 5942 10426
rect 5976 10392 6154 10426
rect 5926 10390 6154 10392
rect 5926 10382 5992 10390
rect 6054 10340 6154 10390
rect 6248 10420 6314 10430
rect 6406 10420 6506 10478
rect 6248 10386 6264 10420
rect 6298 10386 6506 10420
rect 6586 10438 6640 10454
rect 6586 10404 6596 10438
rect 6630 10436 6640 10438
rect 6714 10436 6814 10478
rect 6630 10406 6814 10436
rect 6630 10404 6640 10406
rect 6586 10388 6640 10404
rect 6248 10376 6314 10386
rect 6406 10342 6506 10386
rect 6714 10342 6814 10406
rect 1456 10204 1556 10230
rect 1744 10204 1844 10230
rect 2076 10204 2176 10230
rect 2418 10204 2518 10230
rect 2822 10204 2922 10230
rect 3166 10204 3266 10230
rect 3788 10214 3888 10240
rect 4096 10214 4196 10240
rect 4448 10216 4548 10242
rect 4756 10216 4856 10242
rect 5746 10214 5846 10240
rect 6054 10214 6154 10240
rect 6406 10216 6506 10242
rect 6714 10216 6814 10242
rect 1456 9440 1556 9466
rect 1744 9440 1844 9466
rect 2076 9440 2176 9466
rect 2418 9440 2518 9466
rect 2822 9440 2922 9466
rect 3166 9440 3266 9466
rect 3788 9450 3888 9476
rect 4096 9450 4196 9476
rect 4448 9450 4548 9476
rect 4756 9450 4856 9476
rect 5746 9450 5846 9476
rect 6054 9450 6154 9476
rect 6406 9450 6506 9476
rect 6714 9450 6814 9476
rect 1456 9212 1556 9240
rect 1239 9187 1556 9212
rect 1239 9153 1269 9187
rect 1303 9153 1556 9187
rect 1239 9129 1556 9153
rect 1456 9102 1556 9129
rect 1744 9187 1844 9240
rect 1744 9153 1773 9187
rect 1807 9153 1844 9187
rect 1744 9102 1844 9153
rect 2076 9197 2176 9240
rect 2418 9218 2518 9240
rect 2621 9218 2707 9219
rect 2076 9185 2325 9197
rect 2076 9151 2273 9185
rect 2307 9151 2325 9185
rect 2076 9139 2325 9151
rect 2418 9195 2712 9218
rect 2418 9161 2647 9195
rect 2681 9161 2712 9195
rect 2076 9102 2176 9139
rect 2418 9127 2712 9161
rect 2822 9183 2922 9240
rect 2822 9149 2857 9183
rect 2891 9149 2922 9183
rect 2418 9102 2518 9127
rect 2822 9102 2922 9149
rect 3019 9193 3073 9199
rect 3166 9193 3266 9240
rect 3019 9183 3266 9193
rect 3019 9149 3029 9183
rect 3063 9149 3266 9183
rect 3654 9209 3720 9217
rect 3788 9209 3888 9250
rect 3654 9207 3888 9209
rect 3654 9173 3670 9207
rect 3704 9173 3888 9207
rect 3654 9170 3888 9173
rect 3654 9163 3720 9170
rect 3019 9139 3266 9149
rect 3019 9133 3073 9139
rect 3166 9102 3266 9139
rect 3788 9112 3888 9170
rect 3968 9200 4034 9208
rect 4096 9200 4196 9250
rect 3968 9198 4196 9200
rect 3968 9164 3984 9198
rect 4018 9164 4196 9198
rect 3968 9161 4196 9164
rect 3968 9154 4034 9161
rect 4096 9112 4196 9161
rect 4290 9192 4356 9202
rect 4448 9192 4548 9250
rect 4290 9158 4306 9192
rect 4340 9158 4548 9192
rect 4627 9210 4681 9226
rect 4627 9176 4637 9210
rect 4671 9208 4681 9210
rect 4756 9208 4856 9250
rect 4671 9177 4856 9208
rect 4671 9176 4681 9177
rect 4627 9160 4681 9176
rect 4290 9157 4548 9158
rect 4290 9148 4356 9157
rect 4448 9114 4548 9157
rect 4756 9114 4856 9177
rect 5612 9210 5678 9218
rect 5746 9210 5846 9250
rect 5612 9208 5846 9210
rect 5612 9174 5628 9208
rect 5662 9174 5846 9208
rect 5612 9170 5846 9174
rect 5612 9164 5678 9170
rect 5746 9112 5846 9170
rect 5926 9200 5992 9208
rect 6054 9200 6154 9250
rect 5926 9198 6154 9200
rect 5926 9164 5942 9198
rect 5976 9164 6154 9198
rect 5926 9162 6154 9164
rect 5926 9154 5992 9162
rect 6054 9112 6154 9162
rect 6248 9192 6314 9202
rect 6406 9192 6506 9250
rect 6248 9158 6264 9192
rect 6298 9158 6506 9192
rect 6586 9210 6640 9226
rect 6586 9176 6596 9210
rect 6630 9208 6640 9210
rect 6714 9208 6814 9250
rect 6630 9178 6814 9208
rect 6630 9176 6640 9178
rect 6586 9160 6640 9176
rect 6248 9148 6314 9158
rect 6406 9114 6506 9158
rect 6714 9114 6814 9178
rect 1456 8976 1556 9002
rect 1744 8976 1844 9002
rect 2076 8976 2176 9002
rect 2418 8976 2518 9002
rect 2822 8976 2922 9002
rect 3166 8976 3266 9002
rect 3788 8986 3888 9012
rect 4096 8986 4196 9012
rect 4448 8988 4548 9014
rect 4756 8988 4856 9014
rect 5746 8986 5846 9012
rect 6054 8986 6154 9012
rect 6406 8988 6506 9014
rect 6714 8988 6814 9014
rect 1456 8212 1556 8238
rect 1744 8212 1844 8238
rect 2076 8212 2176 8238
rect 2418 8212 2518 8238
rect 2822 8212 2922 8238
rect 3166 8212 3266 8238
rect 3788 8222 3888 8248
rect 4096 8222 4196 8248
rect 4448 8222 4548 8248
rect 4756 8222 4856 8248
rect 5746 8222 5846 8248
rect 6054 8222 6154 8248
rect 6406 8222 6506 8248
rect 6714 8222 6814 8248
rect 1456 7984 1556 8012
rect 1239 7959 1556 7984
rect 1239 7925 1269 7959
rect 1303 7925 1556 7959
rect 1239 7901 1556 7925
rect 1456 7874 1556 7901
rect 1744 7959 1844 8012
rect 1744 7925 1773 7959
rect 1807 7925 1844 7959
rect 1744 7874 1844 7925
rect 2076 7969 2176 8012
rect 2418 7990 2518 8012
rect 2621 7990 2707 7991
rect 2076 7957 2325 7969
rect 2076 7923 2273 7957
rect 2307 7923 2325 7957
rect 2076 7911 2325 7923
rect 2418 7967 2712 7990
rect 2418 7933 2647 7967
rect 2681 7933 2712 7967
rect 2076 7874 2176 7911
rect 2418 7899 2712 7933
rect 2822 7955 2922 8012
rect 2822 7921 2857 7955
rect 2891 7921 2922 7955
rect 2418 7874 2518 7899
rect 2822 7874 2922 7921
rect 3019 7965 3073 7971
rect 3166 7965 3266 8012
rect 3019 7955 3266 7965
rect 3019 7921 3029 7955
rect 3063 7921 3266 7955
rect 3654 7981 3720 7989
rect 3788 7981 3888 8022
rect 3654 7979 3888 7981
rect 3654 7945 3670 7979
rect 3704 7945 3888 7979
rect 3654 7942 3888 7945
rect 3654 7935 3720 7942
rect 3019 7911 3266 7921
rect 3019 7905 3073 7911
rect 3166 7874 3266 7911
rect 3788 7884 3888 7942
rect 3968 7972 4034 7980
rect 4096 7972 4196 8022
rect 3968 7970 4196 7972
rect 3968 7936 3984 7970
rect 4018 7936 4196 7970
rect 3968 7933 4196 7936
rect 3968 7926 4034 7933
rect 4096 7884 4196 7933
rect 4290 7964 4356 7974
rect 4448 7964 4548 8022
rect 4290 7930 4306 7964
rect 4340 7930 4548 7964
rect 4627 7982 4681 7998
rect 4627 7948 4637 7982
rect 4671 7980 4681 7982
rect 4756 7980 4856 8022
rect 4671 7949 4856 7980
rect 4671 7948 4681 7949
rect 4627 7932 4681 7948
rect 4290 7929 4548 7930
rect 4290 7920 4356 7929
rect 4448 7886 4548 7929
rect 4756 7886 4856 7949
rect 5612 7982 5678 7990
rect 5746 7982 5846 8022
rect 5612 7980 5846 7982
rect 5612 7946 5628 7980
rect 5662 7946 5846 7980
rect 5612 7942 5846 7946
rect 5612 7936 5678 7942
rect 5746 7884 5846 7942
rect 5926 7972 5992 7980
rect 6054 7972 6154 8022
rect 5926 7970 6154 7972
rect 5926 7936 5942 7970
rect 5976 7936 6154 7970
rect 5926 7934 6154 7936
rect 5926 7926 5992 7934
rect 6054 7884 6154 7934
rect 6248 7964 6314 7974
rect 6406 7964 6506 8022
rect 6248 7930 6264 7964
rect 6298 7930 6506 7964
rect 6586 7982 6640 7998
rect 6586 7948 6596 7982
rect 6630 7980 6640 7982
rect 6714 7980 6814 8022
rect 6630 7950 6814 7980
rect 6630 7948 6640 7950
rect 6586 7932 6640 7948
rect 6248 7920 6314 7930
rect 6406 7886 6506 7930
rect 6714 7886 6814 7950
rect 1456 7748 1556 7774
rect 1744 7748 1844 7774
rect 2076 7748 2176 7774
rect 2418 7748 2518 7774
rect 2822 7748 2922 7774
rect 3166 7748 3266 7774
rect 3788 7758 3888 7784
rect 4096 7758 4196 7784
rect 4448 7760 4548 7786
rect 4756 7760 4856 7786
rect 5746 7758 5846 7784
rect 6054 7758 6154 7784
rect 6406 7760 6506 7786
rect 6714 7760 6814 7786
rect 1456 6984 1556 7010
rect 1744 6984 1844 7010
rect 2076 6984 2176 7010
rect 2418 6984 2518 7010
rect 2822 6984 2922 7010
rect 3166 6984 3266 7010
rect 3788 6994 3888 7020
rect 4096 6994 4196 7020
rect 4448 6994 4548 7020
rect 4756 6994 4856 7020
rect 5746 6994 5846 7020
rect 6054 6994 6154 7020
rect 6406 6994 6506 7020
rect 6714 6994 6814 7020
rect 1456 6756 1556 6784
rect 1239 6731 1556 6756
rect 1239 6697 1269 6731
rect 1303 6697 1556 6731
rect 1239 6673 1556 6697
rect 1456 6646 1556 6673
rect 1744 6731 1844 6784
rect 1744 6697 1773 6731
rect 1807 6697 1844 6731
rect 1744 6646 1844 6697
rect 2076 6741 2176 6784
rect 2418 6762 2518 6784
rect 2621 6762 2707 6763
rect 2076 6729 2325 6741
rect 2076 6695 2273 6729
rect 2307 6695 2325 6729
rect 2076 6683 2325 6695
rect 2418 6739 2712 6762
rect 2418 6705 2647 6739
rect 2681 6705 2712 6739
rect 2076 6646 2176 6683
rect 2418 6671 2712 6705
rect 2822 6727 2922 6784
rect 2822 6693 2857 6727
rect 2891 6693 2922 6727
rect 2418 6646 2518 6671
rect 2822 6646 2922 6693
rect 3019 6737 3073 6743
rect 3166 6737 3266 6784
rect 3019 6727 3266 6737
rect 3019 6693 3029 6727
rect 3063 6693 3266 6727
rect 3654 6753 3720 6761
rect 3788 6753 3888 6794
rect 3654 6751 3888 6753
rect 3654 6717 3670 6751
rect 3704 6717 3888 6751
rect 3654 6714 3888 6717
rect 3654 6707 3720 6714
rect 3019 6683 3266 6693
rect 3019 6677 3073 6683
rect 3166 6646 3266 6683
rect 3788 6656 3888 6714
rect 3968 6744 4034 6752
rect 4096 6744 4196 6794
rect 3968 6742 4196 6744
rect 3968 6708 3984 6742
rect 4018 6708 4196 6742
rect 3968 6705 4196 6708
rect 3968 6698 4034 6705
rect 4096 6656 4196 6705
rect 4290 6736 4356 6746
rect 4448 6736 4548 6794
rect 4290 6702 4306 6736
rect 4340 6702 4548 6736
rect 4627 6754 4681 6770
rect 4627 6720 4637 6754
rect 4671 6752 4681 6754
rect 4756 6752 4856 6794
rect 4671 6721 4856 6752
rect 4671 6720 4681 6721
rect 4627 6704 4681 6720
rect 4290 6701 4548 6702
rect 4290 6692 4356 6701
rect 4448 6658 4548 6701
rect 4756 6658 4856 6721
rect 5612 6754 5678 6762
rect 5746 6754 5846 6794
rect 5612 6752 5846 6754
rect 5612 6718 5628 6752
rect 5662 6718 5846 6752
rect 5612 6714 5846 6718
rect 5612 6708 5678 6714
rect 5746 6656 5846 6714
rect 5926 6744 5992 6752
rect 6054 6744 6154 6794
rect 5926 6742 6154 6744
rect 5926 6708 5942 6742
rect 5976 6708 6154 6742
rect 5926 6706 6154 6708
rect 5926 6698 5992 6706
rect 6054 6656 6154 6706
rect 6248 6736 6314 6746
rect 6406 6736 6506 6794
rect 6248 6702 6264 6736
rect 6298 6702 6506 6736
rect 6586 6754 6640 6770
rect 6586 6720 6596 6754
rect 6630 6752 6640 6754
rect 6714 6752 6814 6794
rect 6630 6722 6814 6752
rect 6630 6720 6640 6722
rect 6586 6704 6640 6720
rect 6248 6692 6314 6702
rect 6406 6658 6506 6702
rect 6714 6658 6814 6722
rect 1456 6520 1556 6546
rect 1744 6520 1844 6546
rect 2076 6520 2176 6546
rect 2418 6520 2518 6546
rect 2822 6520 2922 6546
rect 3166 6520 3266 6546
rect 3788 6530 3888 6556
rect 4096 6530 4196 6556
rect 4448 6532 4548 6558
rect 4756 6532 4856 6558
rect 5746 6530 5846 6556
rect 6054 6530 6154 6556
rect 6406 6532 6506 6558
rect 6714 6532 6814 6558
rect 1456 5756 1556 5782
rect 1744 5756 1844 5782
rect 2076 5756 2176 5782
rect 2418 5756 2518 5782
rect 2822 5756 2922 5782
rect 3166 5756 3266 5782
rect 3788 5766 3888 5792
rect 4096 5766 4196 5792
rect 4448 5766 4548 5792
rect 4756 5766 4856 5792
rect 5746 5766 5846 5792
rect 6054 5766 6154 5792
rect 6406 5766 6506 5792
rect 6714 5766 6814 5792
rect 1456 5528 1556 5556
rect 1239 5503 1556 5528
rect 1239 5469 1269 5503
rect 1303 5469 1556 5503
rect 1239 5445 1556 5469
rect 1456 5418 1556 5445
rect 1744 5503 1844 5556
rect 1744 5469 1773 5503
rect 1807 5469 1844 5503
rect 1744 5418 1844 5469
rect 2076 5513 2176 5556
rect 2418 5534 2518 5556
rect 2621 5534 2707 5535
rect 2076 5501 2325 5513
rect 2076 5467 2273 5501
rect 2307 5467 2325 5501
rect 2076 5455 2325 5467
rect 2418 5511 2712 5534
rect 2418 5477 2647 5511
rect 2681 5477 2712 5511
rect 2076 5418 2176 5455
rect 2418 5443 2712 5477
rect 2822 5499 2922 5556
rect 2822 5465 2857 5499
rect 2891 5465 2922 5499
rect 2418 5418 2518 5443
rect 2822 5418 2922 5465
rect 3019 5509 3073 5515
rect 3166 5509 3266 5556
rect 3019 5499 3266 5509
rect 3019 5465 3029 5499
rect 3063 5465 3266 5499
rect 3654 5525 3720 5533
rect 3788 5525 3888 5566
rect 3654 5523 3888 5525
rect 3654 5489 3670 5523
rect 3704 5489 3888 5523
rect 3654 5486 3888 5489
rect 3654 5479 3720 5486
rect 3019 5455 3266 5465
rect 3019 5449 3073 5455
rect 3166 5418 3266 5455
rect 3788 5428 3888 5486
rect 3968 5516 4034 5524
rect 4096 5516 4196 5566
rect 3968 5514 4196 5516
rect 3968 5480 3984 5514
rect 4018 5480 4196 5514
rect 3968 5477 4196 5480
rect 3968 5470 4034 5477
rect 4096 5428 4196 5477
rect 4290 5508 4356 5518
rect 4448 5508 4548 5566
rect 4290 5474 4306 5508
rect 4340 5474 4548 5508
rect 4627 5526 4681 5542
rect 4627 5492 4637 5526
rect 4671 5524 4681 5526
rect 4756 5524 4856 5566
rect 4671 5493 4856 5524
rect 4671 5492 4681 5493
rect 4627 5476 4681 5492
rect 4290 5473 4548 5474
rect 4290 5464 4356 5473
rect 4448 5430 4548 5473
rect 4756 5430 4856 5493
rect 5612 5526 5678 5534
rect 5746 5526 5846 5566
rect 5612 5524 5846 5526
rect 5612 5490 5628 5524
rect 5662 5490 5846 5524
rect 5612 5486 5846 5490
rect 5612 5480 5678 5486
rect 5746 5428 5846 5486
rect 5926 5516 5992 5524
rect 6054 5516 6154 5566
rect 5926 5514 6154 5516
rect 5926 5480 5942 5514
rect 5976 5480 6154 5514
rect 5926 5478 6154 5480
rect 5926 5470 5992 5478
rect 6054 5428 6154 5478
rect 6248 5508 6314 5518
rect 6406 5508 6506 5566
rect 6248 5474 6264 5508
rect 6298 5474 6506 5508
rect 6586 5526 6640 5542
rect 6586 5492 6596 5526
rect 6630 5524 6640 5526
rect 6714 5524 6814 5566
rect 6630 5494 6814 5524
rect 6630 5492 6640 5494
rect 6586 5476 6640 5492
rect 6248 5464 6314 5474
rect 6406 5430 6506 5474
rect 6714 5430 6814 5494
rect 1456 5292 1556 5318
rect 1744 5292 1844 5318
rect 2076 5292 2176 5318
rect 2418 5292 2518 5318
rect 2822 5292 2922 5318
rect 3166 5292 3266 5318
rect 3788 5302 3888 5328
rect 4096 5302 4196 5328
rect 4448 5304 4548 5330
rect 4756 5304 4856 5330
rect 5746 5302 5846 5328
rect 6054 5302 6154 5328
rect 6406 5304 6506 5330
rect 6714 5304 6814 5330
rect 1456 4528 1556 4554
rect 1744 4528 1844 4554
rect 2076 4528 2176 4554
rect 2418 4528 2518 4554
rect 2822 4528 2922 4554
rect 3166 4528 3266 4554
rect 3788 4538 3888 4564
rect 4096 4538 4196 4564
rect 4448 4538 4548 4564
rect 4756 4538 4856 4564
rect 5746 4538 5846 4564
rect 6054 4538 6154 4564
rect 6406 4538 6506 4564
rect 6714 4538 6814 4564
rect 1456 4300 1556 4328
rect 1239 4275 1556 4300
rect 1239 4241 1269 4275
rect 1303 4241 1556 4275
rect 1239 4217 1556 4241
rect 1456 4190 1556 4217
rect 1744 4275 1844 4328
rect 1744 4241 1773 4275
rect 1807 4241 1844 4275
rect 1744 4190 1844 4241
rect 2076 4285 2176 4328
rect 2418 4306 2518 4328
rect 2621 4306 2707 4307
rect 2076 4273 2325 4285
rect 2076 4239 2273 4273
rect 2307 4239 2325 4273
rect 2076 4227 2325 4239
rect 2418 4283 2712 4306
rect 2418 4249 2647 4283
rect 2681 4249 2712 4283
rect 2076 4190 2176 4227
rect 2418 4215 2712 4249
rect 2822 4271 2922 4328
rect 2822 4237 2857 4271
rect 2891 4237 2922 4271
rect 2418 4190 2518 4215
rect 2822 4190 2922 4237
rect 3019 4281 3073 4287
rect 3166 4281 3266 4328
rect 3019 4271 3266 4281
rect 3019 4237 3029 4271
rect 3063 4237 3266 4271
rect 3654 4297 3720 4305
rect 3788 4297 3888 4338
rect 3654 4295 3888 4297
rect 3654 4261 3670 4295
rect 3704 4261 3888 4295
rect 3654 4258 3888 4261
rect 3654 4251 3720 4258
rect 3019 4227 3266 4237
rect 3019 4221 3073 4227
rect 3166 4190 3266 4227
rect 3788 4200 3888 4258
rect 3968 4288 4034 4296
rect 4096 4288 4196 4338
rect 3968 4286 4196 4288
rect 3968 4252 3984 4286
rect 4018 4252 4196 4286
rect 3968 4249 4196 4252
rect 3968 4242 4034 4249
rect 4096 4200 4196 4249
rect 4290 4280 4356 4290
rect 4448 4280 4548 4338
rect 4290 4246 4306 4280
rect 4340 4246 4548 4280
rect 4627 4298 4681 4314
rect 4627 4264 4637 4298
rect 4671 4296 4681 4298
rect 4756 4296 4856 4338
rect 4671 4265 4856 4296
rect 4671 4264 4681 4265
rect 4627 4248 4681 4264
rect 4290 4245 4548 4246
rect 4290 4236 4356 4245
rect 4448 4202 4548 4245
rect 4756 4202 4856 4265
rect 5612 4298 5678 4306
rect 5746 4298 5846 4338
rect 5612 4296 5846 4298
rect 5612 4262 5628 4296
rect 5662 4262 5846 4296
rect 5612 4258 5846 4262
rect 5612 4252 5678 4258
rect 5746 4200 5846 4258
rect 5926 4288 5992 4296
rect 6054 4288 6154 4338
rect 5926 4286 6154 4288
rect 5926 4252 5942 4286
rect 5976 4252 6154 4286
rect 5926 4250 6154 4252
rect 5926 4242 5992 4250
rect 6054 4200 6154 4250
rect 6248 4280 6314 4290
rect 6406 4280 6506 4338
rect 6248 4246 6264 4280
rect 6298 4246 6506 4280
rect 6586 4298 6640 4314
rect 6586 4264 6596 4298
rect 6630 4296 6640 4298
rect 6714 4296 6814 4338
rect 6630 4266 6814 4296
rect 6630 4264 6640 4266
rect 6586 4248 6640 4264
rect 6248 4236 6314 4246
rect 6406 4202 6506 4246
rect 6714 4202 6814 4266
rect 1456 4064 1556 4090
rect 1744 4064 1844 4090
rect 2076 4064 2176 4090
rect 2418 4064 2518 4090
rect 2822 4064 2922 4090
rect 3166 4064 3266 4090
rect 3788 4074 3888 4100
rect 4096 4074 4196 4100
rect 4448 4076 4548 4102
rect 4756 4076 4856 4102
rect 5746 4074 5846 4100
rect 6054 4074 6154 4100
rect 6406 4076 6506 4102
rect 6714 4076 6814 4102
rect 1456 3300 1556 3326
rect 1744 3300 1844 3326
rect 2076 3300 2176 3326
rect 2418 3300 2518 3326
rect 2822 3300 2922 3326
rect 3166 3300 3266 3326
rect 3788 3310 3888 3336
rect 4096 3310 4196 3336
rect 4448 3310 4548 3336
rect 4756 3310 4856 3336
rect 5746 3310 5846 3336
rect 6054 3310 6154 3336
rect 6406 3310 6506 3336
rect 6714 3310 6814 3336
rect 1456 3072 1556 3100
rect 1239 3047 1556 3072
rect 1239 3013 1269 3047
rect 1303 3013 1556 3047
rect 1239 2989 1556 3013
rect 1456 2962 1556 2989
rect 1744 3047 1844 3100
rect 1744 3013 1773 3047
rect 1807 3013 1844 3047
rect 1744 2962 1844 3013
rect 2076 3057 2176 3100
rect 2418 3078 2518 3100
rect 2621 3078 2707 3079
rect 2076 3045 2325 3057
rect 2076 3011 2273 3045
rect 2307 3011 2325 3045
rect 2076 2999 2325 3011
rect 2418 3055 2712 3078
rect 2418 3021 2647 3055
rect 2681 3021 2712 3055
rect 2076 2962 2176 2999
rect 2418 2987 2712 3021
rect 2822 3043 2922 3100
rect 2822 3009 2857 3043
rect 2891 3009 2922 3043
rect 2418 2962 2518 2987
rect 2822 2962 2922 3009
rect 3019 3053 3073 3059
rect 3166 3053 3266 3100
rect 3019 3043 3266 3053
rect 3019 3009 3029 3043
rect 3063 3009 3266 3043
rect 3654 3069 3720 3077
rect 3788 3069 3888 3110
rect 3654 3067 3888 3069
rect 3654 3033 3670 3067
rect 3704 3033 3888 3067
rect 3654 3030 3888 3033
rect 3654 3023 3720 3030
rect 3019 2999 3266 3009
rect 3019 2993 3073 2999
rect 3166 2962 3266 2999
rect 3788 2972 3888 3030
rect 3968 3060 4034 3068
rect 4096 3060 4196 3110
rect 3968 3058 4196 3060
rect 3968 3024 3984 3058
rect 4018 3024 4196 3058
rect 3968 3021 4196 3024
rect 3968 3014 4034 3021
rect 4096 2972 4196 3021
rect 4290 3052 4356 3062
rect 4448 3052 4548 3110
rect 4290 3018 4306 3052
rect 4340 3018 4548 3052
rect 4627 3070 4681 3086
rect 4627 3036 4637 3070
rect 4671 3068 4681 3070
rect 4756 3068 4856 3110
rect 4671 3037 4856 3068
rect 4671 3036 4681 3037
rect 4627 3020 4681 3036
rect 4290 3017 4548 3018
rect 4290 3008 4356 3017
rect 4448 2974 4548 3017
rect 4756 2974 4856 3037
rect 5612 3070 5678 3078
rect 5746 3070 5846 3110
rect 5612 3068 5846 3070
rect 5612 3034 5628 3068
rect 5662 3034 5846 3068
rect 5612 3030 5846 3034
rect 5612 3024 5678 3030
rect 5746 2972 5846 3030
rect 5926 3060 5992 3068
rect 6054 3060 6154 3110
rect 5926 3058 6154 3060
rect 5926 3024 5942 3058
rect 5976 3024 6154 3058
rect 5926 3022 6154 3024
rect 5926 3014 5992 3022
rect 6054 2972 6154 3022
rect 6248 3052 6314 3062
rect 6406 3052 6506 3110
rect 6248 3018 6264 3052
rect 6298 3018 6506 3052
rect 6586 3070 6640 3086
rect 6586 3036 6596 3070
rect 6630 3068 6640 3070
rect 6714 3068 6814 3110
rect 6630 3038 6814 3068
rect 6630 3036 6640 3038
rect 6586 3020 6640 3036
rect 6248 3008 6314 3018
rect 6406 2974 6506 3018
rect 6714 2974 6814 3038
rect 1456 2836 1556 2862
rect 1744 2836 1844 2862
rect 2076 2836 2176 2862
rect 2418 2836 2518 2862
rect 2822 2836 2922 2862
rect 3166 2836 3266 2862
rect 3788 2846 3888 2872
rect 4096 2846 4196 2872
rect 4448 2848 4548 2874
rect 4756 2848 4856 2874
rect 5746 2846 5846 2872
rect 6054 2846 6154 2872
rect 6406 2848 6506 2874
rect 6714 2848 6814 2874
rect 1456 2072 1556 2098
rect 1744 2072 1844 2098
rect 2076 2072 2176 2098
rect 2418 2072 2518 2098
rect 2822 2072 2922 2098
rect 3166 2072 3266 2098
rect 3788 2082 3888 2108
rect 4096 2082 4196 2108
rect 4448 2082 4548 2108
rect 4756 2082 4856 2108
rect 5746 2082 5846 2108
rect 6054 2082 6154 2108
rect 6406 2082 6506 2108
rect 6714 2082 6814 2108
rect 1456 1844 1556 1872
rect 1239 1819 1556 1844
rect 1239 1785 1269 1819
rect 1303 1785 1556 1819
rect 1239 1761 1556 1785
rect 1456 1734 1556 1761
rect 1744 1819 1844 1872
rect 1744 1785 1773 1819
rect 1807 1785 1844 1819
rect 1744 1734 1844 1785
rect 2076 1829 2176 1872
rect 2418 1850 2518 1872
rect 2621 1850 2707 1851
rect 2076 1817 2325 1829
rect 2076 1783 2273 1817
rect 2307 1783 2325 1817
rect 2076 1771 2325 1783
rect 2418 1827 2712 1850
rect 2418 1793 2647 1827
rect 2681 1793 2712 1827
rect 2076 1734 2176 1771
rect 2418 1759 2712 1793
rect 2822 1815 2922 1872
rect 2822 1781 2857 1815
rect 2891 1781 2922 1815
rect 2418 1734 2518 1759
rect 2822 1734 2922 1781
rect 3019 1825 3073 1831
rect 3166 1825 3266 1872
rect 3019 1815 3266 1825
rect 3019 1781 3029 1815
rect 3063 1781 3266 1815
rect 3654 1841 3720 1849
rect 3788 1841 3888 1882
rect 3654 1839 3888 1841
rect 3654 1805 3670 1839
rect 3704 1805 3888 1839
rect 3654 1802 3888 1805
rect 3654 1795 3720 1802
rect 3019 1771 3266 1781
rect 3019 1765 3073 1771
rect 3166 1734 3266 1771
rect 3788 1744 3888 1802
rect 3968 1832 4034 1840
rect 4096 1832 4196 1882
rect 3968 1830 4196 1832
rect 3968 1796 3984 1830
rect 4018 1796 4196 1830
rect 3968 1793 4196 1796
rect 3968 1786 4034 1793
rect 4096 1744 4196 1793
rect 4290 1824 4356 1834
rect 4448 1824 4548 1882
rect 4290 1790 4306 1824
rect 4340 1790 4548 1824
rect 4627 1842 4681 1858
rect 4627 1808 4637 1842
rect 4671 1840 4681 1842
rect 4756 1840 4856 1882
rect 4671 1809 4856 1840
rect 4671 1808 4681 1809
rect 4627 1792 4681 1808
rect 4290 1789 4548 1790
rect 4290 1780 4356 1789
rect 4448 1746 4548 1789
rect 4756 1746 4856 1809
rect 5612 1842 5678 1850
rect 5746 1842 5846 1882
rect 5612 1840 5846 1842
rect 5612 1806 5628 1840
rect 5662 1806 5846 1840
rect 5612 1802 5846 1806
rect 5612 1796 5678 1802
rect 5746 1744 5846 1802
rect 5926 1832 5992 1840
rect 6054 1832 6154 1882
rect 5926 1830 6154 1832
rect 5926 1796 5942 1830
rect 5976 1796 6154 1830
rect 5926 1794 6154 1796
rect 5926 1786 5992 1794
rect 6054 1744 6154 1794
rect 6248 1824 6314 1834
rect 6406 1824 6506 1882
rect 6248 1790 6264 1824
rect 6298 1790 6506 1824
rect 6586 1842 6640 1858
rect 6586 1808 6596 1842
rect 6630 1840 6640 1842
rect 6714 1840 6814 1882
rect 6630 1810 6814 1840
rect 6630 1808 6640 1810
rect 6586 1792 6640 1808
rect 6248 1780 6314 1790
rect 6406 1746 6506 1790
rect 6714 1746 6814 1810
rect 1456 1608 1556 1634
rect 1744 1608 1844 1634
rect 2076 1608 2176 1634
rect 2418 1608 2518 1634
rect 2822 1608 2922 1634
rect 3166 1608 3266 1634
rect 3788 1618 3888 1644
rect 4096 1618 4196 1644
rect 4448 1620 4548 1646
rect 4756 1620 4856 1646
rect 5746 1618 5846 1644
rect 6054 1618 6154 1644
rect 6406 1620 6506 1646
rect 6714 1620 6814 1646
rect 1456 844 1556 870
rect 1744 844 1844 870
rect 2076 844 2176 870
rect 2418 844 2518 870
rect 2822 844 2922 870
rect 3166 844 3266 870
rect 3788 854 3888 880
rect 4096 854 4196 880
rect 4448 854 4548 880
rect 4756 854 4856 880
rect 1456 616 1556 644
rect 1239 591 1556 616
rect 1239 557 1269 591
rect 1303 557 1556 591
rect 1239 533 1556 557
rect 1456 506 1556 533
rect 1744 591 1844 644
rect 1744 557 1773 591
rect 1807 557 1844 591
rect 1744 506 1844 557
rect 2076 601 2176 644
rect 2418 622 2518 644
rect 2621 622 2707 623
rect 2076 589 2325 601
rect 2076 555 2273 589
rect 2307 555 2325 589
rect 2076 543 2325 555
rect 2418 599 2712 622
rect 2418 565 2647 599
rect 2681 565 2712 599
rect 2076 506 2176 543
rect 2418 531 2712 565
rect 2822 587 2922 644
rect 2822 553 2857 587
rect 2891 553 2922 587
rect 2418 506 2518 531
rect 2822 506 2922 553
rect 3019 597 3073 603
rect 3166 597 3266 644
rect 3019 587 3266 597
rect 3019 553 3029 587
rect 3063 553 3266 587
rect 3654 613 3720 621
rect 3788 613 3888 654
rect 3654 611 3888 613
rect 3654 577 3670 611
rect 3704 577 3888 611
rect 3654 574 3888 577
rect 3654 567 3720 574
rect 3019 543 3266 553
rect 3019 537 3073 543
rect 3166 506 3266 543
rect 3788 516 3888 574
rect 3968 604 4034 612
rect 4096 604 4196 654
rect 3968 602 4196 604
rect 3968 568 3984 602
rect 4018 568 4196 602
rect 3968 565 4196 568
rect 3968 558 4034 565
rect 4096 516 4196 565
rect 4290 596 4356 606
rect 4448 596 4548 654
rect 4290 562 4306 596
rect 4340 562 4548 596
rect 4627 614 4681 630
rect 4627 580 4637 614
rect 4671 612 4681 614
rect 4756 612 4856 654
rect 4671 581 4856 612
rect 4671 580 4681 581
rect 4627 564 4681 580
rect 4290 561 4548 562
rect 4290 552 4356 561
rect 4448 518 4548 561
rect 4756 518 4856 581
rect 1456 380 1556 406
rect 1744 380 1844 406
rect 2076 380 2176 406
rect 2418 380 2518 406
rect 2822 380 2922 406
rect 3166 380 3266 406
rect 3788 390 3888 416
rect 4096 390 4196 416
rect 4448 392 4548 418
rect 4756 392 4856 418
<< polycont >>
rect 1269 18977 1303 19011
rect 1773 18977 1807 19011
rect 2273 18975 2307 19009
rect 2647 18985 2681 19019
rect 2857 18973 2891 19007
rect 3029 18973 3063 19007
rect 3670 18997 3704 19031
rect 3984 18988 4018 19022
rect 4306 18982 4340 19016
rect 4637 19000 4671 19034
rect 5628 18998 5662 19032
rect 5942 18988 5976 19022
rect 6264 18982 6298 19016
rect 6596 19000 6630 19034
rect 1269 17749 1303 17783
rect 1773 17749 1807 17783
rect 2273 17747 2307 17781
rect 2647 17757 2681 17791
rect 2857 17745 2891 17779
rect 3029 17745 3063 17779
rect 3670 17769 3704 17803
rect 3984 17760 4018 17794
rect 4306 17754 4340 17788
rect 4637 17772 4671 17806
rect 5628 17770 5662 17804
rect 5942 17760 5976 17794
rect 6264 17754 6298 17788
rect 6596 17772 6630 17806
rect 1269 16521 1303 16555
rect 1773 16521 1807 16555
rect 2273 16519 2307 16553
rect 2647 16529 2681 16563
rect 2857 16517 2891 16551
rect 3029 16517 3063 16551
rect 3670 16541 3704 16575
rect 3984 16532 4018 16566
rect 4306 16526 4340 16560
rect 4637 16544 4671 16578
rect 5628 16542 5662 16576
rect 5942 16532 5976 16566
rect 6264 16526 6298 16560
rect 6596 16544 6630 16578
rect 1269 15293 1303 15327
rect 1773 15293 1807 15327
rect 2273 15291 2307 15325
rect 2647 15301 2681 15335
rect 2857 15289 2891 15323
rect 3029 15289 3063 15323
rect 3670 15313 3704 15347
rect 3984 15304 4018 15338
rect 4306 15298 4340 15332
rect 4637 15316 4671 15350
rect 5628 15314 5662 15348
rect 5942 15304 5976 15338
rect 6264 15298 6298 15332
rect 6596 15316 6630 15350
rect 1269 14065 1303 14099
rect 1773 14065 1807 14099
rect 2273 14063 2307 14097
rect 2647 14073 2681 14107
rect 2857 14061 2891 14095
rect 3029 14061 3063 14095
rect 3670 14085 3704 14119
rect 3984 14076 4018 14110
rect 4306 14070 4340 14104
rect 4637 14088 4671 14122
rect 5628 14086 5662 14120
rect 5942 14076 5976 14110
rect 6264 14070 6298 14104
rect 6596 14088 6630 14122
rect 1269 12837 1303 12871
rect 1773 12837 1807 12871
rect 2273 12835 2307 12869
rect 2647 12845 2681 12879
rect 2857 12833 2891 12867
rect 3029 12833 3063 12867
rect 3670 12857 3704 12891
rect 3984 12848 4018 12882
rect 4306 12842 4340 12876
rect 4637 12860 4671 12894
rect 5628 12858 5662 12892
rect 5942 12848 5976 12882
rect 6264 12842 6298 12876
rect 6596 12860 6630 12894
rect 1269 11609 1303 11643
rect 1773 11609 1807 11643
rect 2273 11607 2307 11641
rect 2647 11617 2681 11651
rect 2857 11605 2891 11639
rect 3029 11605 3063 11639
rect 3670 11629 3704 11663
rect 3984 11620 4018 11654
rect 4306 11614 4340 11648
rect 4637 11632 4671 11666
rect 5628 11630 5662 11664
rect 5942 11620 5976 11654
rect 6264 11614 6298 11648
rect 6596 11632 6630 11666
rect 1269 10381 1303 10415
rect 1773 10381 1807 10415
rect 2273 10379 2307 10413
rect 2647 10389 2681 10423
rect 2857 10377 2891 10411
rect 3029 10377 3063 10411
rect 3670 10401 3704 10435
rect 3984 10392 4018 10426
rect 4306 10386 4340 10420
rect 4637 10404 4671 10438
rect 5628 10402 5662 10436
rect 5942 10392 5976 10426
rect 6264 10386 6298 10420
rect 6596 10404 6630 10438
rect 1269 9153 1303 9187
rect 1773 9153 1807 9187
rect 2273 9151 2307 9185
rect 2647 9161 2681 9195
rect 2857 9149 2891 9183
rect 3029 9149 3063 9183
rect 3670 9173 3704 9207
rect 3984 9164 4018 9198
rect 4306 9158 4340 9192
rect 4637 9176 4671 9210
rect 5628 9174 5662 9208
rect 5942 9164 5976 9198
rect 6264 9158 6298 9192
rect 6596 9176 6630 9210
rect 1269 7925 1303 7959
rect 1773 7925 1807 7959
rect 2273 7923 2307 7957
rect 2647 7933 2681 7967
rect 2857 7921 2891 7955
rect 3029 7921 3063 7955
rect 3670 7945 3704 7979
rect 3984 7936 4018 7970
rect 4306 7930 4340 7964
rect 4637 7948 4671 7982
rect 5628 7946 5662 7980
rect 5942 7936 5976 7970
rect 6264 7930 6298 7964
rect 6596 7948 6630 7982
rect 1269 6697 1303 6731
rect 1773 6697 1807 6731
rect 2273 6695 2307 6729
rect 2647 6705 2681 6739
rect 2857 6693 2891 6727
rect 3029 6693 3063 6727
rect 3670 6717 3704 6751
rect 3984 6708 4018 6742
rect 4306 6702 4340 6736
rect 4637 6720 4671 6754
rect 5628 6718 5662 6752
rect 5942 6708 5976 6742
rect 6264 6702 6298 6736
rect 6596 6720 6630 6754
rect 1269 5469 1303 5503
rect 1773 5469 1807 5503
rect 2273 5467 2307 5501
rect 2647 5477 2681 5511
rect 2857 5465 2891 5499
rect 3029 5465 3063 5499
rect 3670 5489 3704 5523
rect 3984 5480 4018 5514
rect 4306 5474 4340 5508
rect 4637 5492 4671 5526
rect 5628 5490 5662 5524
rect 5942 5480 5976 5514
rect 6264 5474 6298 5508
rect 6596 5492 6630 5526
rect 1269 4241 1303 4275
rect 1773 4241 1807 4275
rect 2273 4239 2307 4273
rect 2647 4249 2681 4283
rect 2857 4237 2891 4271
rect 3029 4237 3063 4271
rect 3670 4261 3704 4295
rect 3984 4252 4018 4286
rect 4306 4246 4340 4280
rect 4637 4264 4671 4298
rect 5628 4262 5662 4296
rect 5942 4252 5976 4286
rect 6264 4246 6298 4280
rect 6596 4264 6630 4298
rect 1269 3013 1303 3047
rect 1773 3013 1807 3047
rect 2273 3011 2307 3045
rect 2647 3021 2681 3055
rect 2857 3009 2891 3043
rect 3029 3009 3063 3043
rect 3670 3033 3704 3067
rect 3984 3024 4018 3058
rect 4306 3018 4340 3052
rect 4637 3036 4671 3070
rect 5628 3034 5662 3068
rect 5942 3024 5976 3058
rect 6264 3018 6298 3052
rect 6596 3036 6630 3070
rect 1269 1785 1303 1819
rect 1773 1785 1807 1819
rect 2273 1783 2307 1817
rect 2647 1793 2681 1827
rect 2857 1781 2891 1815
rect 3029 1781 3063 1815
rect 3670 1805 3704 1839
rect 3984 1796 4018 1830
rect 4306 1790 4340 1824
rect 4637 1808 4671 1842
rect 5628 1806 5662 1840
rect 5942 1796 5976 1830
rect 6264 1790 6298 1824
rect 6596 1808 6630 1842
rect 1269 557 1303 591
rect 1773 557 1807 591
rect 2273 555 2307 589
rect 2647 565 2681 599
rect 2857 553 2891 587
rect 3029 553 3063 587
rect 3670 577 3704 611
rect 3984 568 4018 602
rect 4306 562 4340 596
rect 4637 580 4671 614
<< mvndiffres >>
rect 544 18837 628 19257
rect 690 18837 774 19257
rect 834 18843 918 19263
rect 988 18843 1072 19263
rect 544 17609 628 18029
rect 690 17609 774 18029
rect 834 17615 918 18035
rect 988 17615 1072 18035
rect 544 16381 628 16801
rect 690 16381 774 16801
rect 834 16387 918 16807
rect 988 16387 1072 16807
rect 544 15153 628 15573
rect 690 15153 774 15573
rect 834 15159 918 15579
rect 988 15159 1072 15579
rect 544 13925 628 14345
rect 690 13925 774 14345
rect 834 13931 918 14351
rect 988 13931 1072 14351
rect 544 12697 628 13117
rect 690 12697 774 13117
rect 834 12703 918 13123
rect 988 12703 1072 13123
rect 544 11469 628 11889
rect 690 11469 774 11889
rect 834 11475 918 11895
rect 988 11475 1072 11895
rect 544 10241 628 10661
rect 690 10241 774 10661
rect 834 10247 918 10667
rect 988 10247 1072 10667
rect 544 9013 628 9433
rect 690 9013 774 9433
rect 834 9019 918 9439
rect 988 9019 1072 9439
rect 544 7785 628 8205
rect 690 7785 774 8205
rect 834 7791 918 8211
rect 988 7791 1072 8211
rect 544 6557 628 6977
rect 690 6557 774 6977
rect 834 6563 918 6983
rect 988 6563 1072 6983
rect 544 5329 628 5749
rect 690 5329 774 5749
rect 834 5335 918 5755
rect 988 5335 1072 5755
rect 544 4101 628 4521
rect 690 4101 774 4521
rect 834 4107 918 4527
rect 988 4107 1072 4527
rect 544 2873 628 3293
rect 690 2873 774 3293
rect 834 2879 918 3299
rect 988 2879 1072 3299
rect 544 1645 628 2065
rect 690 1645 774 2065
rect 834 1651 918 2071
rect 988 1651 1072 2071
rect 544 417 628 837
rect 690 417 774 837
rect 834 423 918 843
rect 988 423 1072 843
<< locali >>
rect 1348 19418 1880 19470
rect 1348 19384 1383 19418
rect 1429 19384 1455 19418
rect 1497 19384 1527 19418
rect 1565 19384 1599 19418
rect 1633 19384 1667 19418
rect 1705 19384 1735 19418
rect 1777 19384 1803 19418
rect 1849 19384 1880 19418
rect 3724 19417 4264 19470
rect 540 19332 569 19348
rect 603 19332 632 19348
rect 540 19314 566 19332
rect 607 19314 632 19332
rect 686 19332 715 19348
rect 749 19332 778 19348
rect 686 19314 710 19332
rect 751 19314 778 19332
rect 830 19337 859 19354
rect 893 19337 922 19354
rect 830 19320 856 19337
rect 897 19320 922 19337
rect 984 19337 1013 19354
rect 1047 19337 1076 19354
rect 984 19320 1009 19337
rect 1050 19320 1076 19337
rect 1348 19330 1880 19384
rect 2627 19337 3073 19391
rect 556 19292 566 19314
rect 607 19292 616 19314
rect 556 19274 616 19292
rect 702 19292 710 19314
rect 751 19292 762 19314
rect 702 19274 762 19292
rect 846 19297 856 19320
rect 897 19297 906 19320
rect 846 19280 906 19297
rect 1000 19297 1009 19320
rect 1050 19297 1060 19320
rect 1000 19280 1060 19297
rect 1410 19249 1444 19268
rect 1410 19181 1444 19183
rect 1410 19145 1444 19147
rect 1410 19060 1444 19079
rect 1568 19249 1602 19268
rect 1568 19181 1602 19183
rect 1568 19145 1602 19147
rect 1568 19060 1602 19079
rect 1698 19249 1732 19268
rect 1698 19181 1732 19183
rect 1698 19145 1732 19147
rect 1698 19060 1732 19079
rect 1856 19249 1890 19268
rect 1856 19181 1890 19183
rect 1856 19145 1890 19147
rect 1856 19060 1890 19079
rect 2030 19249 2064 19268
rect 2030 19181 2064 19183
rect 2030 19145 2064 19147
rect 2030 19060 2064 19079
rect 2188 19249 2222 19268
rect 2188 19181 2222 19183
rect 2188 19145 2222 19147
rect 2188 19060 2222 19079
rect 2372 19249 2406 19268
rect 2372 19181 2406 19183
rect 2372 19145 2406 19147
rect 2372 19060 2406 19079
rect 2530 19249 2564 19268
rect 2627 19187 2681 19337
rect 2776 19249 2810 19268
rect 2530 19181 2564 19183
rect 2530 19145 2564 19147
rect 2530 19060 2564 19079
rect 2625 19165 2703 19187
rect 2625 19131 2647 19165
rect 2681 19131 2703 19165
rect 1255 19030 1318 19042
rect 1251 19011 1322 19030
rect 2625 19027 2703 19131
rect 2776 19181 2810 19183
rect 2776 19145 2810 19147
rect 2776 19060 2810 19079
rect 2934 19249 2968 19268
rect 2934 19181 2968 19183
rect 2934 19145 2968 19147
rect 2934 19060 2968 19079
rect 1773 19018 1807 19027
rect 2271 19021 2309 19027
rect 1251 18977 1269 19011
rect 1303 18977 1322 19011
rect 1251 18959 1322 18977
rect 1766 19011 1814 19018
rect 1766 18977 1773 19011
rect 1807 18977 1814 19011
rect 1766 18970 1814 18977
rect 2261 19009 2319 19021
rect 2261 18975 2273 19009
rect 2307 18975 2319 19009
rect 2615 19019 2713 19027
rect 2615 18985 2647 19019
rect 2681 18985 2713 19019
rect 2857 19014 2891 19023
rect 2615 18978 2713 18985
rect 2850 19007 2898 19014
rect 3019 19007 3073 19337
rect 3724 19383 3773 19417
rect 3831 19383 3841 19417
rect 3903 19383 3909 19417
rect 3975 19383 3977 19417
rect 4011 19383 4013 19417
rect 4079 19383 4085 19417
rect 4147 19383 4157 19417
rect 4215 19383 4264 19417
rect 3724 19330 4264 19383
rect 5682 19416 6222 19470
rect 5682 19382 5732 19416
rect 5790 19382 5800 19416
rect 5862 19382 5868 19416
rect 5934 19382 5936 19416
rect 5970 19382 5972 19416
rect 6038 19382 6044 19416
rect 6106 19382 6116 19416
rect 6174 19382 6222 19416
rect 5682 19330 6222 19382
rect 3120 19249 3154 19268
rect 3120 19181 3154 19183
rect 3120 19145 3154 19147
rect 3120 19060 3154 19079
rect 3278 19249 3312 19268
rect 3278 19181 3312 19183
rect 3278 19145 3312 19147
rect 3278 19060 3312 19079
rect 3742 19259 3776 19278
rect 3742 19191 3776 19193
rect 3742 19155 3776 19157
rect 3742 19070 3776 19089
rect 3900 19259 3934 19278
rect 3900 19191 3934 19193
rect 3900 19155 3934 19157
rect 3900 19070 3934 19089
rect 4050 19259 4084 19278
rect 4050 19191 4084 19193
rect 4050 19155 4084 19157
rect 4050 19070 4084 19089
rect 4208 19259 4242 19278
rect 4208 19191 4242 19193
rect 4208 19155 4242 19157
rect 4208 19070 4242 19089
rect 4402 19259 4436 19278
rect 4402 19191 4436 19193
rect 4402 19155 4436 19157
rect 4402 19070 4436 19089
rect 4560 19259 4594 19278
rect 4560 19191 4594 19193
rect 4560 19155 4594 19157
rect 4560 19070 4594 19089
rect 4710 19259 4744 19278
rect 4710 19191 4744 19193
rect 4710 19155 4744 19157
rect 4710 19070 4744 19089
rect 4868 19259 4902 19278
rect 4868 19191 4902 19193
rect 4868 19155 4902 19157
rect 4868 19070 4902 19089
rect 5700 19260 5734 19278
rect 5700 19192 5734 19194
rect 5700 19156 5734 19158
rect 5700 19070 5734 19090
rect 5858 19260 5892 19278
rect 5858 19192 5892 19194
rect 5858 19156 5892 19158
rect 5858 19070 5892 19090
rect 6008 19260 6042 19278
rect 6008 19192 6042 19194
rect 6008 19156 6042 19158
rect 6008 19070 6042 19090
rect 6166 19260 6200 19278
rect 6166 19192 6200 19194
rect 6166 19156 6200 19158
rect 6166 19070 6200 19090
rect 6360 19260 6394 19278
rect 6360 19192 6394 19194
rect 6360 19156 6394 19158
rect 6360 19070 6394 19090
rect 6518 19260 6552 19278
rect 6518 19192 6552 19194
rect 6518 19156 6552 19158
rect 6518 19070 6552 19090
rect 6668 19260 6702 19278
rect 6668 19192 6702 19194
rect 6668 19156 6702 19158
rect 6668 19070 6702 19090
rect 6826 19260 6860 19278
rect 6826 19192 6860 19194
rect 6826 19156 6860 19158
rect 6826 19070 6860 19090
rect 3670 19034 3704 19047
rect 3668 19031 3707 19034
rect 1773 18961 1807 18970
rect 2261 18963 2319 18975
rect 2625 18964 2703 18978
rect 2850 18973 2857 19007
rect 2891 18973 2898 19007
rect 3013 18973 3029 19007
rect 3063 18973 3079 19007
rect 3668 18997 3670 19031
rect 3704 18997 3707 19031
rect 3984 19025 4018 19038
rect 5628 19034 5662 19048
rect 3668 18995 3707 18997
rect 3982 19022 4021 19025
rect 3670 18981 3704 18995
rect 3982 18988 3984 19022
rect 4018 18988 4021 19022
rect 3982 18986 4021 18988
rect 4306 19017 4340 19032
rect 4306 19016 4341 19017
rect 2850 18966 2898 18973
rect 1255 18947 1318 18959
rect 2271 18957 2309 18963
rect 1410 18893 1444 18930
rect 556 18804 616 18820
rect 556 18780 565 18804
rect 606 18780 616 18804
rect 702 18804 762 18820
rect 702 18780 712 18804
rect 753 18780 762 18804
rect 846 18809 906 18826
rect 846 18786 856 18809
rect 897 18786 906 18809
rect 1000 18810 1060 18826
rect 1410 18822 1444 18859
rect 1568 18893 1602 18930
rect 1568 18822 1602 18859
rect 1698 18893 1732 18930
rect 1698 18822 1732 18859
rect 1856 18893 1890 18930
rect 1856 18822 1890 18859
rect 2030 18893 2064 18930
rect 2030 18822 2064 18859
rect 2188 18893 2222 18930
rect 2188 18822 2222 18859
rect 2352 18893 2420 18936
rect 2352 18859 2372 18893
rect 2406 18859 2420 18893
rect 1000 18786 1010 18810
rect 1051 18786 1060 18810
rect 540 18764 565 18780
rect 606 18764 632 18780
rect 540 18746 569 18764
rect 603 18746 632 18764
rect 686 18764 712 18780
rect 753 18764 778 18780
rect 686 18746 715 18764
rect 749 18746 778 18764
rect 830 18769 856 18786
rect 897 18769 922 18786
rect 830 18752 859 18769
rect 893 18752 922 18769
rect 984 18770 1010 18786
rect 1051 18770 1076 18786
rect 984 18752 1013 18770
rect 1047 18752 1076 18770
rect 1324 18716 1960 18780
rect 1324 18682 1353 18716
rect 1407 18682 1421 18716
rect 1479 18682 1489 18716
rect 1551 18682 1557 18716
rect 1623 18682 1625 18716
rect 1659 18682 1661 18716
rect 1727 18682 1733 18716
rect 1795 18682 1805 18716
rect 1863 18682 1877 18716
rect 1931 18682 1960 18716
rect 1324 18640 1960 18682
rect 2352 18691 2420 18859
rect 2530 18893 2564 18930
rect 2530 18822 2564 18859
rect 2352 18657 2369 18691
rect 2403 18657 2420 18691
rect 2352 18640 2420 18657
rect 2642 18595 2696 18964
rect 2857 18957 2891 18966
rect 3019 18963 3073 18973
rect 3984 18972 4018 18986
rect 4340 18982 4341 19016
rect 4621 19000 4637 19034
rect 4671 19000 4687 19034
rect 5626 19032 5666 19034
rect 5626 18998 5628 19032
rect 5662 18998 5666 19032
rect 5942 19026 5976 19038
rect 5626 18996 5666 18998
rect 5940 19022 5980 19026
rect 5628 18982 5662 18996
rect 5940 18988 5942 19022
rect 5976 18988 5980 19022
rect 5940 18986 5980 18988
rect 6264 19018 6298 19032
rect 6264 19016 6300 19018
rect 4306 18966 4340 18982
rect 5942 18972 5976 18986
rect 6298 18982 6300 19016
rect 6580 19000 6596 19034
rect 6630 19000 6646 19034
rect 6264 18966 6298 18982
rect 2776 18893 2810 18930
rect 2776 18822 2810 18859
rect 2934 18893 2968 18930
rect 2934 18822 2968 18859
rect 3120 18893 3154 18930
rect 3120 18822 3154 18859
rect 3278 18893 3312 18930
rect 3278 18822 3312 18859
rect 3742 18903 3776 18940
rect 3742 18832 3776 18869
rect 3900 18903 3934 18940
rect 3900 18832 3934 18869
rect 4050 18903 4084 18940
rect 4050 18832 4084 18869
rect 4208 18903 4242 18940
rect 4208 18832 4242 18869
rect 4402 18905 4436 18942
rect 4402 18834 4436 18871
rect 4560 18905 4594 18942
rect 4560 18834 4594 18871
rect 4710 18905 4744 18942
rect 4710 18834 4744 18871
rect 4868 18905 4902 18942
rect 4868 18834 4902 18871
rect 5700 18904 5734 18940
rect 5700 18832 5734 18870
rect 5858 18904 5892 18940
rect 5858 18832 5892 18870
rect 6008 18904 6042 18940
rect 6008 18832 6042 18870
rect 6166 18904 6200 18940
rect 6166 18832 6200 18870
rect 6360 18906 6394 18942
rect 6360 18834 6394 18872
rect 6518 18906 6552 18942
rect 6518 18834 6552 18872
rect 6668 18906 6702 18942
rect 6668 18834 6702 18872
rect 6826 18906 6860 18942
rect 6826 18834 6860 18872
rect 3704 18727 4244 18780
rect 3704 18693 3741 18727
rect 3787 18693 3813 18727
rect 3855 18693 3885 18727
rect 3923 18693 3957 18727
rect 3991 18693 4025 18727
rect 4063 18693 4093 18727
rect 4135 18693 4161 18727
rect 4207 18693 4244 18727
rect 3704 18640 4244 18693
rect 5662 18728 6202 18780
rect 5662 18694 5700 18728
rect 5746 18694 5772 18728
rect 5814 18694 5844 18728
rect 5882 18694 5916 18728
rect 5950 18694 5984 18728
rect 6022 18694 6052 18728
rect 6094 18694 6120 18728
rect 6166 18694 6202 18728
rect 5662 18640 6202 18694
rect 1348 18190 1880 18242
rect 1348 18156 1383 18190
rect 1429 18156 1455 18190
rect 1497 18156 1527 18190
rect 1565 18156 1599 18190
rect 1633 18156 1667 18190
rect 1705 18156 1735 18190
rect 1777 18156 1803 18190
rect 1849 18156 1880 18190
rect 3724 18189 4264 18242
rect 540 18104 569 18120
rect 603 18104 632 18120
rect 540 18086 566 18104
rect 607 18086 632 18104
rect 686 18104 715 18120
rect 749 18104 778 18120
rect 686 18086 710 18104
rect 751 18086 778 18104
rect 830 18109 859 18126
rect 893 18109 922 18126
rect 830 18092 856 18109
rect 897 18092 922 18109
rect 984 18109 1013 18126
rect 1047 18109 1076 18126
rect 984 18092 1009 18109
rect 1050 18092 1076 18109
rect 1348 18102 1880 18156
rect 2627 18109 3073 18163
rect 556 18064 566 18086
rect 607 18064 616 18086
rect 556 18046 616 18064
rect 702 18064 710 18086
rect 751 18064 762 18086
rect 702 18046 762 18064
rect 846 18069 856 18092
rect 897 18069 906 18092
rect 846 18052 906 18069
rect 1000 18069 1009 18092
rect 1050 18069 1060 18092
rect 1000 18052 1060 18069
rect 1410 18021 1444 18040
rect 1410 17953 1444 17955
rect 1410 17917 1444 17919
rect 1410 17832 1444 17851
rect 1568 18021 1602 18040
rect 1568 17953 1602 17955
rect 1568 17917 1602 17919
rect 1568 17832 1602 17851
rect 1698 18021 1732 18040
rect 1698 17953 1732 17955
rect 1698 17917 1732 17919
rect 1698 17832 1732 17851
rect 1856 18021 1890 18040
rect 1856 17953 1890 17955
rect 1856 17917 1890 17919
rect 1856 17832 1890 17851
rect 2030 18021 2064 18040
rect 2030 17953 2064 17955
rect 2030 17917 2064 17919
rect 2030 17832 2064 17851
rect 2188 18021 2222 18040
rect 2188 17953 2222 17955
rect 2188 17917 2222 17919
rect 2188 17832 2222 17851
rect 2372 18021 2406 18040
rect 2372 17953 2406 17955
rect 2372 17917 2406 17919
rect 2372 17832 2406 17851
rect 2530 18021 2564 18040
rect 2627 17959 2681 18109
rect 2776 18021 2810 18040
rect 2530 17953 2564 17955
rect 2530 17917 2564 17919
rect 2530 17832 2564 17851
rect 2625 17937 2703 17959
rect 2625 17903 2647 17937
rect 2681 17903 2703 17937
rect 1255 17802 1318 17814
rect 1251 17783 1322 17802
rect 2625 17799 2703 17903
rect 2776 17953 2810 17955
rect 2776 17917 2810 17919
rect 2776 17832 2810 17851
rect 2934 18021 2968 18040
rect 2934 17953 2968 17955
rect 2934 17917 2968 17919
rect 2934 17832 2968 17851
rect 1773 17790 1807 17799
rect 2271 17793 2309 17799
rect 1251 17749 1269 17783
rect 1303 17749 1322 17783
rect 1251 17731 1322 17749
rect 1766 17783 1814 17790
rect 1766 17749 1773 17783
rect 1807 17749 1814 17783
rect 1766 17742 1814 17749
rect 2261 17781 2319 17793
rect 2261 17747 2273 17781
rect 2307 17747 2319 17781
rect 2615 17791 2713 17799
rect 2615 17757 2647 17791
rect 2681 17757 2713 17791
rect 2857 17786 2891 17795
rect 2615 17750 2713 17757
rect 2850 17779 2898 17786
rect 3019 17779 3073 18109
rect 3724 18155 3773 18189
rect 3831 18155 3841 18189
rect 3903 18155 3909 18189
rect 3975 18155 3977 18189
rect 4011 18155 4013 18189
rect 4079 18155 4085 18189
rect 4147 18155 4157 18189
rect 4215 18155 4264 18189
rect 3724 18102 4264 18155
rect 5682 18188 6222 18242
rect 5682 18154 5732 18188
rect 5790 18154 5800 18188
rect 5862 18154 5868 18188
rect 5934 18154 5936 18188
rect 5970 18154 5972 18188
rect 6038 18154 6044 18188
rect 6106 18154 6116 18188
rect 6174 18154 6222 18188
rect 5682 18102 6222 18154
rect 3120 18021 3154 18040
rect 3120 17953 3154 17955
rect 3120 17917 3154 17919
rect 3120 17832 3154 17851
rect 3278 18021 3312 18040
rect 3278 17953 3312 17955
rect 3278 17917 3312 17919
rect 3278 17832 3312 17851
rect 3742 18031 3776 18050
rect 3742 17963 3776 17965
rect 3742 17927 3776 17929
rect 3742 17842 3776 17861
rect 3900 18031 3934 18050
rect 3900 17963 3934 17965
rect 3900 17927 3934 17929
rect 3900 17842 3934 17861
rect 4050 18031 4084 18050
rect 4050 17963 4084 17965
rect 4050 17927 4084 17929
rect 4050 17842 4084 17861
rect 4208 18031 4242 18050
rect 4208 17963 4242 17965
rect 4208 17927 4242 17929
rect 4208 17842 4242 17861
rect 4402 18031 4436 18050
rect 4402 17963 4436 17965
rect 4402 17927 4436 17929
rect 4402 17842 4436 17861
rect 4560 18031 4594 18050
rect 4560 17963 4594 17965
rect 4560 17927 4594 17929
rect 4560 17842 4594 17861
rect 4710 18031 4744 18050
rect 4710 17963 4744 17965
rect 4710 17927 4744 17929
rect 4710 17842 4744 17861
rect 4868 18031 4902 18050
rect 4868 17963 4902 17965
rect 4868 17927 4902 17929
rect 4868 17842 4902 17861
rect 5700 18032 5734 18050
rect 5700 17964 5734 17966
rect 5700 17928 5734 17930
rect 5700 17842 5734 17862
rect 5858 18032 5892 18050
rect 5858 17964 5892 17966
rect 5858 17928 5892 17930
rect 5858 17842 5892 17862
rect 6008 18032 6042 18050
rect 6008 17964 6042 17966
rect 6008 17928 6042 17930
rect 6008 17842 6042 17862
rect 6166 18032 6200 18050
rect 6166 17964 6200 17966
rect 6166 17928 6200 17930
rect 6166 17842 6200 17862
rect 6360 18032 6394 18050
rect 6360 17964 6394 17966
rect 6360 17928 6394 17930
rect 6360 17842 6394 17862
rect 6518 18032 6552 18050
rect 6518 17964 6552 17966
rect 6518 17928 6552 17930
rect 6518 17842 6552 17862
rect 6668 18032 6702 18050
rect 6668 17964 6702 17966
rect 6668 17928 6702 17930
rect 6668 17842 6702 17862
rect 6826 18032 6860 18050
rect 6826 17964 6860 17966
rect 6826 17928 6860 17930
rect 6826 17842 6860 17862
rect 3670 17806 3704 17819
rect 3668 17803 3707 17806
rect 1773 17733 1807 17742
rect 2261 17735 2319 17747
rect 2625 17736 2703 17750
rect 2850 17745 2857 17779
rect 2891 17745 2898 17779
rect 3013 17745 3029 17779
rect 3063 17745 3079 17779
rect 3668 17769 3670 17803
rect 3704 17769 3707 17803
rect 3984 17797 4018 17810
rect 5628 17806 5662 17820
rect 3668 17767 3707 17769
rect 3982 17794 4021 17797
rect 3670 17753 3704 17767
rect 3982 17760 3984 17794
rect 4018 17760 4021 17794
rect 3982 17758 4021 17760
rect 4306 17789 4340 17804
rect 4306 17788 4341 17789
rect 2850 17738 2898 17745
rect 1255 17719 1318 17731
rect 2271 17729 2309 17735
rect 1410 17665 1444 17702
rect 556 17576 616 17592
rect 556 17552 565 17576
rect 606 17552 616 17576
rect 702 17576 762 17592
rect 702 17552 712 17576
rect 753 17552 762 17576
rect 846 17581 906 17598
rect 846 17558 856 17581
rect 897 17558 906 17581
rect 1000 17582 1060 17598
rect 1410 17594 1444 17631
rect 1568 17665 1602 17702
rect 1568 17594 1602 17631
rect 1698 17665 1732 17702
rect 1698 17594 1732 17631
rect 1856 17665 1890 17702
rect 1856 17594 1890 17631
rect 2030 17665 2064 17702
rect 2030 17594 2064 17631
rect 2188 17665 2222 17702
rect 2188 17594 2222 17631
rect 2352 17665 2420 17708
rect 2352 17631 2372 17665
rect 2406 17631 2420 17665
rect 1000 17558 1010 17582
rect 1051 17558 1060 17582
rect 540 17536 565 17552
rect 606 17536 632 17552
rect 540 17518 569 17536
rect 603 17518 632 17536
rect 686 17536 712 17552
rect 753 17536 778 17552
rect 686 17518 715 17536
rect 749 17518 778 17536
rect 830 17541 856 17558
rect 897 17541 922 17558
rect 830 17524 859 17541
rect 893 17524 922 17541
rect 984 17542 1010 17558
rect 1051 17542 1076 17558
rect 984 17524 1013 17542
rect 1047 17524 1076 17542
rect 1324 17488 1960 17552
rect 1324 17454 1353 17488
rect 1407 17454 1421 17488
rect 1479 17454 1489 17488
rect 1551 17454 1557 17488
rect 1623 17454 1625 17488
rect 1659 17454 1661 17488
rect 1727 17454 1733 17488
rect 1795 17454 1805 17488
rect 1863 17454 1877 17488
rect 1931 17454 1960 17488
rect 1324 17412 1960 17454
rect 2352 17463 2420 17631
rect 2530 17665 2564 17702
rect 2530 17594 2564 17631
rect 2352 17429 2369 17463
rect 2403 17429 2420 17463
rect 2352 17412 2420 17429
rect 2642 17367 2696 17736
rect 2857 17729 2891 17738
rect 3019 17735 3073 17745
rect 3984 17744 4018 17758
rect 4340 17754 4341 17788
rect 4621 17772 4637 17806
rect 4671 17772 4687 17806
rect 5626 17804 5666 17806
rect 5626 17770 5628 17804
rect 5662 17770 5666 17804
rect 5942 17798 5976 17810
rect 5626 17768 5666 17770
rect 5940 17794 5980 17798
rect 5628 17754 5662 17768
rect 5940 17760 5942 17794
rect 5976 17760 5980 17794
rect 5940 17758 5980 17760
rect 6264 17790 6298 17804
rect 6264 17788 6300 17790
rect 4306 17738 4340 17754
rect 5942 17744 5976 17758
rect 6298 17754 6300 17788
rect 6580 17772 6596 17806
rect 6630 17772 6646 17806
rect 6264 17738 6298 17754
rect 2776 17665 2810 17702
rect 2776 17594 2810 17631
rect 2934 17665 2968 17702
rect 2934 17594 2968 17631
rect 3120 17665 3154 17702
rect 3120 17594 3154 17631
rect 3278 17665 3312 17702
rect 3278 17594 3312 17631
rect 3742 17675 3776 17712
rect 3742 17604 3776 17641
rect 3900 17675 3934 17712
rect 3900 17604 3934 17641
rect 4050 17675 4084 17712
rect 4050 17604 4084 17641
rect 4208 17675 4242 17712
rect 4208 17604 4242 17641
rect 4402 17677 4436 17714
rect 4402 17606 4436 17643
rect 4560 17677 4594 17714
rect 4560 17606 4594 17643
rect 4710 17677 4744 17714
rect 4710 17606 4744 17643
rect 4868 17677 4902 17714
rect 4868 17606 4902 17643
rect 5700 17676 5734 17712
rect 5700 17604 5734 17642
rect 5858 17676 5892 17712
rect 5858 17604 5892 17642
rect 6008 17676 6042 17712
rect 6008 17604 6042 17642
rect 6166 17676 6200 17712
rect 6166 17604 6200 17642
rect 6360 17678 6394 17714
rect 6360 17606 6394 17644
rect 6518 17678 6552 17714
rect 6518 17606 6552 17644
rect 6668 17678 6702 17714
rect 6668 17606 6702 17644
rect 6826 17678 6860 17714
rect 6826 17606 6860 17644
rect 3704 17499 4244 17552
rect 3704 17465 3741 17499
rect 3787 17465 3813 17499
rect 3855 17465 3885 17499
rect 3923 17465 3957 17499
rect 3991 17465 4025 17499
rect 4063 17465 4093 17499
rect 4135 17465 4161 17499
rect 4207 17465 4244 17499
rect 3704 17412 4244 17465
rect 5662 17500 6202 17552
rect 5662 17466 5700 17500
rect 5746 17466 5772 17500
rect 5814 17466 5844 17500
rect 5882 17466 5916 17500
rect 5950 17466 5984 17500
rect 6022 17466 6052 17500
rect 6094 17466 6120 17500
rect 6166 17466 6202 17500
rect 5662 17412 6202 17466
rect 1348 16962 1880 17014
rect 1348 16928 1383 16962
rect 1429 16928 1455 16962
rect 1497 16928 1527 16962
rect 1565 16928 1599 16962
rect 1633 16928 1667 16962
rect 1705 16928 1735 16962
rect 1777 16928 1803 16962
rect 1849 16928 1880 16962
rect 3724 16961 4264 17014
rect 540 16876 569 16892
rect 603 16876 632 16892
rect 540 16858 566 16876
rect 607 16858 632 16876
rect 686 16876 715 16892
rect 749 16876 778 16892
rect 686 16858 710 16876
rect 751 16858 778 16876
rect 830 16881 859 16898
rect 893 16881 922 16898
rect 830 16864 856 16881
rect 897 16864 922 16881
rect 984 16881 1013 16898
rect 1047 16881 1076 16898
rect 984 16864 1009 16881
rect 1050 16864 1076 16881
rect 1348 16874 1880 16928
rect 2627 16881 3073 16935
rect 556 16836 566 16858
rect 607 16836 616 16858
rect 556 16818 616 16836
rect 702 16836 710 16858
rect 751 16836 762 16858
rect 702 16818 762 16836
rect 846 16841 856 16864
rect 897 16841 906 16864
rect 846 16824 906 16841
rect 1000 16841 1009 16864
rect 1050 16841 1060 16864
rect 1000 16824 1060 16841
rect 1410 16793 1444 16812
rect 1410 16725 1444 16727
rect 1410 16689 1444 16691
rect 1410 16604 1444 16623
rect 1568 16793 1602 16812
rect 1568 16725 1602 16727
rect 1568 16689 1602 16691
rect 1568 16604 1602 16623
rect 1698 16793 1732 16812
rect 1698 16725 1732 16727
rect 1698 16689 1732 16691
rect 1698 16604 1732 16623
rect 1856 16793 1890 16812
rect 1856 16725 1890 16727
rect 1856 16689 1890 16691
rect 1856 16604 1890 16623
rect 2030 16793 2064 16812
rect 2030 16725 2064 16727
rect 2030 16689 2064 16691
rect 2030 16604 2064 16623
rect 2188 16793 2222 16812
rect 2188 16725 2222 16727
rect 2188 16689 2222 16691
rect 2188 16604 2222 16623
rect 2372 16793 2406 16812
rect 2372 16725 2406 16727
rect 2372 16689 2406 16691
rect 2372 16604 2406 16623
rect 2530 16793 2564 16812
rect 2627 16731 2681 16881
rect 2776 16793 2810 16812
rect 2530 16725 2564 16727
rect 2530 16689 2564 16691
rect 2530 16604 2564 16623
rect 2625 16709 2703 16731
rect 2625 16675 2647 16709
rect 2681 16675 2703 16709
rect 1255 16574 1318 16586
rect 1251 16555 1322 16574
rect 2625 16571 2703 16675
rect 2776 16725 2810 16727
rect 2776 16689 2810 16691
rect 2776 16604 2810 16623
rect 2934 16793 2968 16812
rect 2934 16725 2968 16727
rect 2934 16689 2968 16691
rect 2934 16604 2968 16623
rect 1773 16562 1807 16571
rect 2271 16565 2309 16571
rect 1251 16521 1269 16555
rect 1303 16521 1322 16555
rect 1251 16503 1322 16521
rect 1766 16555 1814 16562
rect 1766 16521 1773 16555
rect 1807 16521 1814 16555
rect 1766 16514 1814 16521
rect 2261 16553 2319 16565
rect 2261 16519 2273 16553
rect 2307 16519 2319 16553
rect 2615 16563 2713 16571
rect 2615 16529 2647 16563
rect 2681 16529 2713 16563
rect 2857 16558 2891 16567
rect 2615 16522 2713 16529
rect 2850 16551 2898 16558
rect 3019 16551 3073 16881
rect 3724 16927 3773 16961
rect 3831 16927 3841 16961
rect 3903 16927 3909 16961
rect 3975 16927 3977 16961
rect 4011 16927 4013 16961
rect 4079 16927 4085 16961
rect 4147 16927 4157 16961
rect 4215 16927 4264 16961
rect 3724 16874 4264 16927
rect 5682 16960 6222 17014
rect 5682 16926 5732 16960
rect 5790 16926 5800 16960
rect 5862 16926 5868 16960
rect 5934 16926 5936 16960
rect 5970 16926 5972 16960
rect 6038 16926 6044 16960
rect 6106 16926 6116 16960
rect 6174 16926 6222 16960
rect 5682 16874 6222 16926
rect 3120 16793 3154 16812
rect 3120 16725 3154 16727
rect 3120 16689 3154 16691
rect 3120 16604 3154 16623
rect 3278 16793 3312 16812
rect 3278 16725 3312 16727
rect 3278 16689 3312 16691
rect 3278 16604 3312 16623
rect 3742 16803 3776 16822
rect 3742 16735 3776 16737
rect 3742 16699 3776 16701
rect 3742 16614 3776 16633
rect 3900 16803 3934 16822
rect 3900 16735 3934 16737
rect 3900 16699 3934 16701
rect 3900 16614 3934 16633
rect 4050 16803 4084 16822
rect 4050 16735 4084 16737
rect 4050 16699 4084 16701
rect 4050 16614 4084 16633
rect 4208 16803 4242 16822
rect 4208 16735 4242 16737
rect 4208 16699 4242 16701
rect 4208 16614 4242 16633
rect 4402 16803 4436 16822
rect 4402 16735 4436 16737
rect 4402 16699 4436 16701
rect 4402 16614 4436 16633
rect 4560 16803 4594 16822
rect 4560 16735 4594 16737
rect 4560 16699 4594 16701
rect 4560 16614 4594 16633
rect 4710 16803 4744 16822
rect 4710 16735 4744 16737
rect 4710 16699 4744 16701
rect 4710 16614 4744 16633
rect 4868 16803 4902 16822
rect 4868 16735 4902 16737
rect 4868 16699 4902 16701
rect 4868 16614 4902 16633
rect 5700 16804 5734 16822
rect 5700 16736 5734 16738
rect 5700 16700 5734 16702
rect 5700 16614 5734 16634
rect 5858 16804 5892 16822
rect 5858 16736 5892 16738
rect 5858 16700 5892 16702
rect 5858 16614 5892 16634
rect 6008 16804 6042 16822
rect 6008 16736 6042 16738
rect 6008 16700 6042 16702
rect 6008 16614 6042 16634
rect 6166 16804 6200 16822
rect 6166 16736 6200 16738
rect 6166 16700 6200 16702
rect 6166 16614 6200 16634
rect 6360 16804 6394 16822
rect 6360 16736 6394 16738
rect 6360 16700 6394 16702
rect 6360 16614 6394 16634
rect 6518 16804 6552 16822
rect 6518 16736 6552 16738
rect 6518 16700 6552 16702
rect 6518 16614 6552 16634
rect 6668 16804 6702 16822
rect 6668 16736 6702 16738
rect 6668 16700 6702 16702
rect 6668 16614 6702 16634
rect 6826 16804 6860 16822
rect 6826 16736 6860 16738
rect 6826 16700 6860 16702
rect 6826 16614 6860 16634
rect 3670 16578 3704 16591
rect 3668 16575 3707 16578
rect 1773 16505 1807 16514
rect 2261 16507 2319 16519
rect 2625 16508 2703 16522
rect 2850 16517 2857 16551
rect 2891 16517 2898 16551
rect 3013 16517 3029 16551
rect 3063 16517 3079 16551
rect 3668 16541 3670 16575
rect 3704 16541 3707 16575
rect 3984 16569 4018 16582
rect 5628 16578 5662 16592
rect 3668 16539 3707 16541
rect 3982 16566 4021 16569
rect 3670 16525 3704 16539
rect 3982 16532 3984 16566
rect 4018 16532 4021 16566
rect 3982 16530 4021 16532
rect 4306 16561 4340 16576
rect 4306 16560 4341 16561
rect 2850 16510 2898 16517
rect 1255 16491 1318 16503
rect 2271 16501 2309 16507
rect 1410 16437 1444 16474
rect 556 16348 616 16364
rect 556 16324 565 16348
rect 606 16324 616 16348
rect 702 16348 762 16364
rect 702 16324 712 16348
rect 753 16324 762 16348
rect 846 16353 906 16370
rect 846 16330 856 16353
rect 897 16330 906 16353
rect 1000 16354 1060 16370
rect 1410 16366 1444 16403
rect 1568 16437 1602 16474
rect 1568 16366 1602 16403
rect 1698 16437 1732 16474
rect 1698 16366 1732 16403
rect 1856 16437 1890 16474
rect 1856 16366 1890 16403
rect 2030 16437 2064 16474
rect 2030 16366 2064 16403
rect 2188 16437 2222 16474
rect 2188 16366 2222 16403
rect 2352 16437 2420 16480
rect 2352 16403 2372 16437
rect 2406 16403 2420 16437
rect 1000 16330 1010 16354
rect 1051 16330 1060 16354
rect 540 16308 565 16324
rect 606 16308 632 16324
rect 540 16290 569 16308
rect 603 16290 632 16308
rect 686 16308 712 16324
rect 753 16308 778 16324
rect 686 16290 715 16308
rect 749 16290 778 16308
rect 830 16313 856 16330
rect 897 16313 922 16330
rect 830 16296 859 16313
rect 893 16296 922 16313
rect 984 16314 1010 16330
rect 1051 16314 1076 16330
rect 984 16296 1013 16314
rect 1047 16296 1076 16314
rect 1324 16260 1960 16324
rect 1324 16226 1353 16260
rect 1407 16226 1421 16260
rect 1479 16226 1489 16260
rect 1551 16226 1557 16260
rect 1623 16226 1625 16260
rect 1659 16226 1661 16260
rect 1727 16226 1733 16260
rect 1795 16226 1805 16260
rect 1863 16226 1877 16260
rect 1931 16226 1960 16260
rect 1324 16184 1960 16226
rect 2352 16235 2420 16403
rect 2530 16437 2564 16474
rect 2530 16366 2564 16403
rect 2352 16201 2369 16235
rect 2403 16201 2420 16235
rect 2352 16184 2420 16201
rect 2642 16139 2696 16508
rect 2857 16501 2891 16510
rect 3019 16507 3073 16517
rect 3984 16516 4018 16530
rect 4340 16526 4341 16560
rect 4621 16544 4637 16578
rect 4671 16544 4687 16578
rect 5626 16576 5666 16578
rect 5626 16542 5628 16576
rect 5662 16542 5666 16576
rect 5942 16570 5976 16582
rect 5626 16540 5666 16542
rect 5940 16566 5980 16570
rect 5628 16526 5662 16540
rect 5940 16532 5942 16566
rect 5976 16532 5980 16566
rect 5940 16530 5980 16532
rect 6264 16562 6298 16576
rect 6264 16560 6300 16562
rect 4306 16510 4340 16526
rect 5942 16516 5976 16530
rect 6298 16526 6300 16560
rect 6580 16544 6596 16578
rect 6630 16544 6646 16578
rect 6264 16510 6298 16526
rect 2776 16437 2810 16474
rect 2776 16366 2810 16403
rect 2934 16437 2968 16474
rect 2934 16366 2968 16403
rect 3120 16437 3154 16474
rect 3120 16366 3154 16403
rect 3278 16437 3312 16474
rect 3278 16366 3312 16403
rect 3742 16447 3776 16484
rect 3742 16376 3776 16413
rect 3900 16447 3934 16484
rect 3900 16376 3934 16413
rect 4050 16447 4084 16484
rect 4050 16376 4084 16413
rect 4208 16447 4242 16484
rect 4208 16376 4242 16413
rect 4402 16449 4436 16486
rect 4402 16378 4436 16415
rect 4560 16449 4594 16486
rect 4560 16378 4594 16415
rect 4710 16449 4744 16486
rect 4710 16378 4744 16415
rect 4868 16449 4902 16486
rect 4868 16378 4902 16415
rect 5700 16448 5734 16484
rect 5700 16376 5734 16414
rect 5858 16448 5892 16484
rect 5858 16376 5892 16414
rect 6008 16448 6042 16484
rect 6008 16376 6042 16414
rect 6166 16448 6200 16484
rect 6166 16376 6200 16414
rect 6360 16450 6394 16486
rect 6360 16378 6394 16416
rect 6518 16450 6552 16486
rect 6518 16378 6552 16416
rect 6668 16450 6702 16486
rect 6668 16378 6702 16416
rect 6826 16450 6860 16486
rect 6826 16378 6860 16416
rect 3704 16271 4244 16324
rect 3704 16237 3741 16271
rect 3787 16237 3813 16271
rect 3855 16237 3885 16271
rect 3923 16237 3957 16271
rect 3991 16237 4025 16271
rect 4063 16237 4093 16271
rect 4135 16237 4161 16271
rect 4207 16237 4244 16271
rect 3704 16184 4244 16237
rect 5662 16272 6202 16324
rect 5662 16238 5700 16272
rect 5746 16238 5772 16272
rect 5814 16238 5844 16272
rect 5882 16238 5916 16272
rect 5950 16238 5984 16272
rect 6022 16238 6052 16272
rect 6094 16238 6120 16272
rect 6166 16238 6202 16272
rect 5662 16184 6202 16238
rect 1348 15734 1880 15786
rect 1348 15700 1383 15734
rect 1429 15700 1455 15734
rect 1497 15700 1527 15734
rect 1565 15700 1599 15734
rect 1633 15700 1667 15734
rect 1705 15700 1735 15734
rect 1777 15700 1803 15734
rect 1849 15700 1880 15734
rect 3724 15733 4264 15786
rect 540 15648 569 15664
rect 603 15648 632 15664
rect 540 15630 566 15648
rect 607 15630 632 15648
rect 686 15648 715 15664
rect 749 15648 778 15664
rect 686 15630 710 15648
rect 751 15630 778 15648
rect 830 15653 859 15670
rect 893 15653 922 15670
rect 830 15636 856 15653
rect 897 15636 922 15653
rect 984 15653 1013 15670
rect 1047 15653 1076 15670
rect 984 15636 1009 15653
rect 1050 15636 1076 15653
rect 1348 15646 1880 15700
rect 2627 15653 3073 15707
rect 556 15608 566 15630
rect 607 15608 616 15630
rect 556 15590 616 15608
rect 702 15608 710 15630
rect 751 15608 762 15630
rect 702 15590 762 15608
rect 846 15613 856 15636
rect 897 15613 906 15636
rect 846 15596 906 15613
rect 1000 15613 1009 15636
rect 1050 15613 1060 15636
rect 1000 15596 1060 15613
rect 1410 15565 1444 15584
rect 1410 15497 1444 15499
rect 1410 15461 1444 15463
rect 1410 15376 1444 15395
rect 1568 15565 1602 15584
rect 1568 15497 1602 15499
rect 1568 15461 1602 15463
rect 1568 15376 1602 15395
rect 1698 15565 1732 15584
rect 1698 15497 1732 15499
rect 1698 15461 1732 15463
rect 1698 15376 1732 15395
rect 1856 15565 1890 15584
rect 1856 15497 1890 15499
rect 1856 15461 1890 15463
rect 1856 15376 1890 15395
rect 2030 15565 2064 15584
rect 2030 15497 2064 15499
rect 2030 15461 2064 15463
rect 2030 15376 2064 15395
rect 2188 15565 2222 15584
rect 2188 15497 2222 15499
rect 2188 15461 2222 15463
rect 2188 15376 2222 15395
rect 2372 15565 2406 15584
rect 2372 15497 2406 15499
rect 2372 15461 2406 15463
rect 2372 15376 2406 15395
rect 2530 15565 2564 15584
rect 2627 15503 2681 15653
rect 2776 15565 2810 15584
rect 2530 15497 2564 15499
rect 2530 15461 2564 15463
rect 2530 15376 2564 15395
rect 2625 15481 2703 15503
rect 2625 15447 2647 15481
rect 2681 15447 2703 15481
rect 1255 15346 1318 15358
rect 1251 15327 1322 15346
rect 2625 15343 2703 15447
rect 2776 15497 2810 15499
rect 2776 15461 2810 15463
rect 2776 15376 2810 15395
rect 2934 15565 2968 15584
rect 2934 15497 2968 15499
rect 2934 15461 2968 15463
rect 2934 15376 2968 15395
rect 1773 15334 1807 15343
rect 2271 15337 2309 15343
rect 1251 15293 1269 15327
rect 1303 15293 1322 15327
rect 1251 15275 1322 15293
rect 1766 15327 1814 15334
rect 1766 15293 1773 15327
rect 1807 15293 1814 15327
rect 1766 15286 1814 15293
rect 2261 15325 2319 15337
rect 2261 15291 2273 15325
rect 2307 15291 2319 15325
rect 2615 15335 2713 15343
rect 2615 15301 2647 15335
rect 2681 15301 2713 15335
rect 2857 15330 2891 15339
rect 2615 15294 2713 15301
rect 2850 15323 2898 15330
rect 3019 15323 3073 15653
rect 3724 15699 3773 15733
rect 3831 15699 3841 15733
rect 3903 15699 3909 15733
rect 3975 15699 3977 15733
rect 4011 15699 4013 15733
rect 4079 15699 4085 15733
rect 4147 15699 4157 15733
rect 4215 15699 4264 15733
rect 3724 15646 4264 15699
rect 5682 15732 6222 15786
rect 5682 15698 5732 15732
rect 5790 15698 5800 15732
rect 5862 15698 5868 15732
rect 5934 15698 5936 15732
rect 5970 15698 5972 15732
rect 6038 15698 6044 15732
rect 6106 15698 6116 15732
rect 6174 15698 6222 15732
rect 5682 15646 6222 15698
rect 3120 15565 3154 15584
rect 3120 15497 3154 15499
rect 3120 15461 3154 15463
rect 3120 15376 3154 15395
rect 3278 15565 3312 15584
rect 3278 15497 3312 15499
rect 3278 15461 3312 15463
rect 3278 15376 3312 15395
rect 3742 15575 3776 15594
rect 3742 15507 3776 15509
rect 3742 15471 3776 15473
rect 3742 15386 3776 15405
rect 3900 15575 3934 15594
rect 3900 15507 3934 15509
rect 3900 15471 3934 15473
rect 3900 15386 3934 15405
rect 4050 15575 4084 15594
rect 4050 15507 4084 15509
rect 4050 15471 4084 15473
rect 4050 15386 4084 15405
rect 4208 15575 4242 15594
rect 4208 15507 4242 15509
rect 4208 15471 4242 15473
rect 4208 15386 4242 15405
rect 4402 15575 4436 15594
rect 4402 15507 4436 15509
rect 4402 15471 4436 15473
rect 4402 15386 4436 15405
rect 4560 15575 4594 15594
rect 4560 15507 4594 15509
rect 4560 15471 4594 15473
rect 4560 15386 4594 15405
rect 4710 15575 4744 15594
rect 4710 15507 4744 15509
rect 4710 15471 4744 15473
rect 4710 15386 4744 15405
rect 4868 15575 4902 15594
rect 4868 15507 4902 15509
rect 4868 15471 4902 15473
rect 4868 15386 4902 15405
rect 5700 15576 5734 15594
rect 5700 15508 5734 15510
rect 5700 15472 5734 15474
rect 5700 15386 5734 15406
rect 5858 15576 5892 15594
rect 5858 15508 5892 15510
rect 5858 15472 5892 15474
rect 5858 15386 5892 15406
rect 6008 15576 6042 15594
rect 6008 15508 6042 15510
rect 6008 15472 6042 15474
rect 6008 15386 6042 15406
rect 6166 15576 6200 15594
rect 6166 15508 6200 15510
rect 6166 15472 6200 15474
rect 6166 15386 6200 15406
rect 6360 15576 6394 15594
rect 6360 15508 6394 15510
rect 6360 15472 6394 15474
rect 6360 15386 6394 15406
rect 6518 15576 6552 15594
rect 6518 15508 6552 15510
rect 6518 15472 6552 15474
rect 6518 15386 6552 15406
rect 6668 15576 6702 15594
rect 6668 15508 6702 15510
rect 6668 15472 6702 15474
rect 6668 15386 6702 15406
rect 6826 15576 6860 15594
rect 6826 15508 6860 15510
rect 6826 15472 6860 15474
rect 6826 15386 6860 15406
rect 3670 15350 3704 15363
rect 3668 15347 3707 15350
rect 1773 15277 1807 15286
rect 2261 15279 2319 15291
rect 2625 15280 2703 15294
rect 2850 15289 2857 15323
rect 2891 15289 2898 15323
rect 3013 15289 3029 15323
rect 3063 15289 3079 15323
rect 3668 15313 3670 15347
rect 3704 15313 3707 15347
rect 3984 15341 4018 15354
rect 5628 15350 5662 15364
rect 3668 15311 3707 15313
rect 3982 15338 4021 15341
rect 3670 15297 3704 15311
rect 3982 15304 3984 15338
rect 4018 15304 4021 15338
rect 3982 15302 4021 15304
rect 4306 15333 4340 15348
rect 4306 15332 4341 15333
rect 2850 15282 2898 15289
rect 1255 15263 1318 15275
rect 2271 15273 2309 15279
rect 1410 15209 1444 15246
rect 556 15120 616 15136
rect 556 15096 565 15120
rect 606 15096 616 15120
rect 702 15120 762 15136
rect 702 15096 712 15120
rect 753 15096 762 15120
rect 846 15125 906 15142
rect 846 15102 856 15125
rect 897 15102 906 15125
rect 1000 15126 1060 15142
rect 1410 15138 1444 15175
rect 1568 15209 1602 15246
rect 1568 15138 1602 15175
rect 1698 15209 1732 15246
rect 1698 15138 1732 15175
rect 1856 15209 1890 15246
rect 1856 15138 1890 15175
rect 2030 15209 2064 15246
rect 2030 15138 2064 15175
rect 2188 15209 2222 15246
rect 2188 15138 2222 15175
rect 2352 15209 2420 15252
rect 2352 15175 2372 15209
rect 2406 15175 2420 15209
rect 1000 15102 1010 15126
rect 1051 15102 1060 15126
rect 540 15080 565 15096
rect 606 15080 632 15096
rect 540 15062 569 15080
rect 603 15062 632 15080
rect 686 15080 712 15096
rect 753 15080 778 15096
rect 686 15062 715 15080
rect 749 15062 778 15080
rect 830 15085 856 15102
rect 897 15085 922 15102
rect 830 15068 859 15085
rect 893 15068 922 15085
rect 984 15086 1010 15102
rect 1051 15086 1076 15102
rect 984 15068 1013 15086
rect 1047 15068 1076 15086
rect 1324 15032 1960 15096
rect 1324 14998 1353 15032
rect 1407 14998 1421 15032
rect 1479 14998 1489 15032
rect 1551 14998 1557 15032
rect 1623 14998 1625 15032
rect 1659 14998 1661 15032
rect 1727 14998 1733 15032
rect 1795 14998 1805 15032
rect 1863 14998 1877 15032
rect 1931 14998 1960 15032
rect 1324 14956 1960 14998
rect 2352 15007 2420 15175
rect 2530 15209 2564 15246
rect 2530 15138 2564 15175
rect 2352 14973 2369 15007
rect 2403 14973 2420 15007
rect 2352 14956 2420 14973
rect 2642 14911 2696 15280
rect 2857 15273 2891 15282
rect 3019 15279 3073 15289
rect 3984 15288 4018 15302
rect 4340 15298 4341 15332
rect 4621 15316 4637 15350
rect 4671 15316 4687 15350
rect 5626 15348 5666 15350
rect 5626 15314 5628 15348
rect 5662 15314 5666 15348
rect 5942 15342 5976 15354
rect 5626 15312 5666 15314
rect 5940 15338 5980 15342
rect 5628 15298 5662 15312
rect 5940 15304 5942 15338
rect 5976 15304 5980 15338
rect 5940 15302 5980 15304
rect 6264 15334 6298 15348
rect 6264 15332 6300 15334
rect 4306 15282 4340 15298
rect 5942 15288 5976 15302
rect 6298 15298 6300 15332
rect 6580 15316 6596 15350
rect 6630 15316 6646 15350
rect 6264 15282 6298 15298
rect 2776 15209 2810 15246
rect 2776 15138 2810 15175
rect 2934 15209 2968 15246
rect 2934 15138 2968 15175
rect 3120 15209 3154 15246
rect 3120 15138 3154 15175
rect 3278 15209 3312 15246
rect 3278 15138 3312 15175
rect 3742 15219 3776 15256
rect 3742 15148 3776 15185
rect 3900 15219 3934 15256
rect 3900 15148 3934 15185
rect 4050 15219 4084 15256
rect 4050 15148 4084 15185
rect 4208 15219 4242 15256
rect 4208 15148 4242 15185
rect 4402 15221 4436 15258
rect 4402 15150 4436 15187
rect 4560 15221 4594 15258
rect 4560 15150 4594 15187
rect 4710 15221 4744 15258
rect 4710 15150 4744 15187
rect 4868 15221 4902 15258
rect 4868 15150 4902 15187
rect 5700 15220 5734 15256
rect 5700 15148 5734 15186
rect 5858 15220 5892 15256
rect 5858 15148 5892 15186
rect 6008 15220 6042 15256
rect 6008 15148 6042 15186
rect 6166 15220 6200 15256
rect 6166 15148 6200 15186
rect 6360 15222 6394 15258
rect 6360 15150 6394 15188
rect 6518 15222 6552 15258
rect 6518 15150 6552 15188
rect 6668 15222 6702 15258
rect 6668 15150 6702 15188
rect 6826 15222 6860 15258
rect 6826 15150 6860 15188
rect 3704 15043 4244 15096
rect 3704 15009 3741 15043
rect 3787 15009 3813 15043
rect 3855 15009 3885 15043
rect 3923 15009 3957 15043
rect 3991 15009 4025 15043
rect 4063 15009 4093 15043
rect 4135 15009 4161 15043
rect 4207 15009 4244 15043
rect 3704 14956 4244 15009
rect 5662 15044 6202 15096
rect 5662 15010 5700 15044
rect 5746 15010 5772 15044
rect 5814 15010 5844 15044
rect 5882 15010 5916 15044
rect 5950 15010 5984 15044
rect 6022 15010 6052 15044
rect 6094 15010 6120 15044
rect 6166 15010 6202 15044
rect 5662 14956 6202 15010
rect 1348 14506 1880 14558
rect 1348 14472 1383 14506
rect 1429 14472 1455 14506
rect 1497 14472 1527 14506
rect 1565 14472 1599 14506
rect 1633 14472 1667 14506
rect 1705 14472 1735 14506
rect 1777 14472 1803 14506
rect 1849 14472 1880 14506
rect 3724 14505 4264 14558
rect 540 14420 569 14436
rect 603 14420 632 14436
rect 540 14402 566 14420
rect 607 14402 632 14420
rect 686 14420 715 14436
rect 749 14420 778 14436
rect 686 14402 710 14420
rect 751 14402 778 14420
rect 830 14425 859 14442
rect 893 14425 922 14442
rect 830 14408 856 14425
rect 897 14408 922 14425
rect 984 14425 1013 14442
rect 1047 14425 1076 14442
rect 984 14408 1009 14425
rect 1050 14408 1076 14425
rect 1348 14418 1880 14472
rect 2627 14425 3073 14479
rect 556 14380 566 14402
rect 607 14380 616 14402
rect 556 14362 616 14380
rect 702 14380 710 14402
rect 751 14380 762 14402
rect 702 14362 762 14380
rect 846 14385 856 14408
rect 897 14385 906 14408
rect 846 14368 906 14385
rect 1000 14385 1009 14408
rect 1050 14385 1060 14408
rect 1000 14368 1060 14385
rect 1410 14337 1444 14356
rect 1410 14269 1444 14271
rect 1410 14233 1444 14235
rect 1410 14148 1444 14167
rect 1568 14337 1602 14356
rect 1568 14269 1602 14271
rect 1568 14233 1602 14235
rect 1568 14148 1602 14167
rect 1698 14337 1732 14356
rect 1698 14269 1732 14271
rect 1698 14233 1732 14235
rect 1698 14148 1732 14167
rect 1856 14337 1890 14356
rect 1856 14269 1890 14271
rect 1856 14233 1890 14235
rect 1856 14148 1890 14167
rect 2030 14337 2064 14356
rect 2030 14269 2064 14271
rect 2030 14233 2064 14235
rect 2030 14148 2064 14167
rect 2188 14337 2222 14356
rect 2188 14269 2222 14271
rect 2188 14233 2222 14235
rect 2188 14148 2222 14167
rect 2372 14337 2406 14356
rect 2372 14269 2406 14271
rect 2372 14233 2406 14235
rect 2372 14148 2406 14167
rect 2530 14337 2564 14356
rect 2627 14275 2681 14425
rect 2776 14337 2810 14356
rect 2530 14269 2564 14271
rect 2530 14233 2564 14235
rect 2530 14148 2564 14167
rect 2625 14253 2703 14275
rect 2625 14219 2647 14253
rect 2681 14219 2703 14253
rect 1255 14118 1318 14130
rect 1251 14099 1322 14118
rect 2625 14115 2703 14219
rect 2776 14269 2810 14271
rect 2776 14233 2810 14235
rect 2776 14148 2810 14167
rect 2934 14337 2968 14356
rect 2934 14269 2968 14271
rect 2934 14233 2968 14235
rect 2934 14148 2968 14167
rect 1773 14106 1807 14115
rect 2271 14109 2309 14115
rect 1251 14065 1269 14099
rect 1303 14065 1322 14099
rect 1251 14047 1322 14065
rect 1766 14099 1814 14106
rect 1766 14065 1773 14099
rect 1807 14065 1814 14099
rect 1766 14058 1814 14065
rect 2261 14097 2319 14109
rect 2261 14063 2273 14097
rect 2307 14063 2319 14097
rect 2615 14107 2713 14115
rect 2615 14073 2647 14107
rect 2681 14073 2713 14107
rect 2857 14102 2891 14111
rect 2615 14066 2713 14073
rect 2850 14095 2898 14102
rect 3019 14095 3073 14425
rect 3724 14471 3773 14505
rect 3831 14471 3841 14505
rect 3903 14471 3909 14505
rect 3975 14471 3977 14505
rect 4011 14471 4013 14505
rect 4079 14471 4085 14505
rect 4147 14471 4157 14505
rect 4215 14471 4264 14505
rect 3724 14418 4264 14471
rect 5682 14504 6222 14558
rect 5682 14470 5732 14504
rect 5790 14470 5800 14504
rect 5862 14470 5868 14504
rect 5934 14470 5936 14504
rect 5970 14470 5972 14504
rect 6038 14470 6044 14504
rect 6106 14470 6116 14504
rect 6174 14470 6222 14504
rect 5682 14418 6222 14470
rect 3120 14337 3154 14356
rect 3120 14269 3154 14271
rect 3120 14233 3154 14235
rect 3120 14148 3154 14167
rect 3278 14337 3312 14356
rect 3278 14269 3312 14271
rect 3278 14233 3312 14235
rect 3278 14148 3312 14167
rect 3742 14347 3776 14366
rect 3742 14279 3776 14281
rect 3742 14243 3776 14245
rect 3742 14158 3776 14177
rect 3900 14347 3934 14366
rect 3900 14279 3934 14281
rect 3900 14243 3934 14245
rect 3900 14158 3934 14177
rect 4050 14347 4084 14366
rect 4050 14279 4084 14281
rect 4050 14243 4084 14245
rect 4050 14158 4084 14177
rect 4208 14347 4242 14366
rect 4208 14279 4242 14281
rect 4208 14243 4242 14245
rect 4208 14158 4242 14177
rect 4402 14347 4436 14366
rect 4402 14279 4436 14281
rect 4402 14243 4436 14245
rect 4402 14158 4436 14177
rect 4560 14347 4594 14366
rect 4560 14279 4594 14281
rect 4560 14243 4594 14245
rect 4560 14158 4594 14177
rect 4710 14347 4744 14366
rect 4710 14279 4744 14281
rect 4710 14243 4744 14245
rect 4710 14158 4744 14177
rect 4868 14347 4902 14366
rect 4868 14279 4902 14281
rect 4868 14243 4902 14245
rect 4868 14158 4902 14177
rect 5700 14348 5734 14366
rect 5700 14280 5734 14282
rect 5700 14244 5734 14246
rect 5700 14158 5734 14178
rect 5858 14348 5892 14366
rect 5858 14280 5892 14282
rect 5858 14244 5892 14246
rect 5858 14158 5892 14178
rect 6008 14348 6042 14366
rect 6008 14280 6042 14282
rect 6008 14244 6042 14246
rect 6008 14158 6042 14178
rect 6166 14348 6200 14366
rect 6166 14280 6200 14282
rect 6166 14244 6200 14246
rect 6166 14158 6200 14178
rect 6360 14348 6394 14366
rect 6360 14280 6394 14282
rect 6360 14244 6394 14246
rect 6360 14158 6394 14178
rect 6518 14348 6552 14366
rect 6518 14280 6552 14282
rect 6518 14244 6552 14246
rect 6518 14158 6552 14178
rect 6668 14348 6702 14366
rect 6668 14280 6702 14282
rect 6668 14244 6702 14246
rect 6668 14158 6702 14178
rect 6826 14348 6860 14366
rect 6826 14280 6860 14282
rect 6826 14244 6860 14246
rect 6826 14158 6860 14178
rect 3670 14122 3704 14135
rect 3668 14119 3707 14122
rect 1773 14049 1807 14058
rect 2261 14051 2319 14063
rect 2625 14052 2703 14066
rect 2850 14061 2857 14095
rect 2891 14061 2898 14095
rect 3013 14061 3029 14095
rect 3063 14061 3079 14095
rect 3668 14085 3670 14119
rect 3704 14085 3707 14119
rect 3984 14113 4018 14126
rect 5628 14122 5662 14136
rect 3668 14083 3707 14085
rect 3982 14110 4021 14113
rect 3670 14069 3704 14083
rect 3982 14076 3984 14110
rect 4018 14076 4021 14110
rect 3982 14074 4021 14076
rect 4306 14105 4340 14120
rect 4306 14104 4341 14105
rect 2850 14054 2898 14061
rect 1255 14035 1318 14047
rect 2271 14045 2309 14051
rect 1410 13981 1444 14018
rect 556 13892 616 13908
rect 556 13868 565 13892
rect 606 13868 616 13892
rect 702 13892 762 13908
rect 702 13868 712 13892
rect 753 13868 762 13892
rect 846 13897 906 13914
rect 846 13874 856 13897
rect 897 13874 906 13897
rect 1000 13898 1060 13914
rect 1410 13910 1444 13947
rect 1568 13981 1602 14018
rect 1568 13910 1602 13947
rect 1698 13981 1732 14018
rect 1698 13910 1732 13947
rect 1856 13981 1890 14018
rect 1856 13910 1890 13947
rect 2030 13981 2064 14018
rect 2030 13910 2064 13947
rect 2188 13981 2222 14018
rect 2188 13910 2222 13947
rect 2352 13981 2420 14024
rect 2352 13947 2372 13981
rect 2406 13947 2420 13981
rect 1000 13874 1010 13898
rect 1051 13874 1060 13898
rect 540 13852 565 13868
rect 606 13852 632 13868
rect 540 13834 569 13852
rect 603 13834 632 13852
rect 686 13852 712 13868
rect 753 13852 778 13868
rect 686 13834 715 13852
rect 749 13834 778 13852
rect 830 13857 856 13874
rect 897 13857 922 13874
rect 830 13840 859 13857
rect 893 13840 922 13857
rect 984 13858 1010 13874
rect 1051 13858 1076 13874
rect 984 13840 1013 13858
rect 1047 13840 1076 13858
rect 1324 13804 1960 13868
rect 1324 13770 1353 13804
rect 1407 13770 1421 13804
rect 1479 13770 1489 13804
rect 1551 13770 1557 13804
rect 1623 13770 1625 13804
rect 1659 13770 1661 13804
rect 1727 13770 1733 13804
rect 1795 13770 1805 13804
rect 1863 13770 1877 13804
rect 1931 13770 1960 13804
rect 1324 13728 1960 13770
rect 2352 13779 2420 13947
rect 2530 13981 2564 14018
rect 2530 13910 2564 13947
rect 2352 13745 2369 13779
rect 2403 13745 2420 13779
rect 2352 13728 2420 13745
rect 2642 13683 2696 14052
rect 2857 14045 2891 14054
rect 3019 14051 3073 14061
rect 3984 14060 4018 14074
rect 4340 14070 4341 14104
rect 4621 14088 4637 14122
rect 4671 14088 4687 14122
rect 5626 14120 5666 14122
rect 5626 14086 5628 14120
rect 5662 14086 5666 14120
rect 5942 14114 5976 14126
rect 5626 14084 5666 14086
rect 5940 14110 5980 14114
rect 5628 14070 5662 14084
rect 5940 14076 5942 14110
rect 5976 14076 5980 14110
rect 5940 14074 5980 14076
rect 6264 14106 6298 14120
rect 6264 14104 6300 14106
rect 4306 14054 4340 14070
rect 5942 14060 5976 14074
rect 6298 14070 6300 14104
rect 6580 14088 6596 14122
rect 6630 14088 6646 14122
rect 6264 14054 6298 14070
rect 2776 13981 2810 14018
rect 2776 13910 2810 13947
rect 2934 13981 2968 14018
rect 2934 13910 2968 13947
rect 3120 13981 3154 14018
rect 3120 13910 3154 13947
rect 3278 13981 3312 14018
rect 3278 13910 3312 13947
rect 3742 13991 3776 14028
rect 3742 13920 3776 13957
rect 3900 13991 3934 14028
rect 3900 13920 3934 13957
rect 4050 13991 4084 14028
rect 4050 13920 4084 13957
rect 4208 13991 4242 14028
rect 4208 13920 4242 13957
rect 4402 13993 4436 14030
rect 4402 13922 4436 13959
rect 4560 13993 4594 14030
rect 4560 13922 4594 13959
rect 4710 13993 4744 14030
rect 4710 13922 4744 13959
rect 4868 13993 4902 14030
rect 4868 13922 4902 13959
rect 5700 13992 5734 14028
rect 5700 13920 5734 13958
rect 5858 13992 5892 14028
rect 5858 13920 5892 13958
rect 6008 13992 6042 14028
rect 6008 13920 6042 13958
rect 6166 13992 6200 14028
rect 6166 13920 6200 13958
rect 6360 13994 6394 14030
rect 6360 13922 6394 13960
rect 6518 13994 6552 14030
rect 6518 13922 6552 13960
rect 6668 13994 6702 14030
rect 6668 13922 6702 13960
rect 6826 13994 6860 14030
rect 6826 13922 6860 13960
rect 3704 13815 4244 13868
rect 3704 13781 3741 13815
rect 3787 13781 3813 13815
rect 3855 13781 3885 13815
rect 3923 13781 3957 13815
rect 3991 13781 4025 13815
rect 4063 13781 4093 13815
rect 4135 13781 4161 13815
rect 4207 13781 4244 13815
rect 3704 13728 4244 13781
rect 5662 13816 6202 13868
rect 5662 13782 5700 13816
rect 5746 13782 5772 13816
rect 5814 13782 5844 13816
rect 5882 13782 5916 13816
rect 5950 13782 5984 13816
rect 6022 13782 6052 13816
rect 6094 13782 6120 13816
rect 6166 13782 6202 13816
rect 5662 13728 6202 13782
rect 1348 13278 1880 13330
rect 1348 13244 1383 13278
rect 1429 13244 1455 13278
rect 1497 13244 1527 13278
rect 1565 13244 1599 13278
rect 1633 13244 1667 13278
rect 1705 13244 1735 13278
rect 1777 13244 1803 13278
rect 1849 13244 1880 13278
rect 3724 13277 4264 13330
rect 540 13192 569 13208
rect 603 13192 632 13208
rect 540 13174 566 13192
rect 607 13174 632 13192
rect 686 13192 715 13208
rect 749 13192 778 13208
rect 686 13174 710 13192
rect 751 13174 778 13192
rect 830 13197 859 13214
rect 893 13197 922 13214
rect 830 13180 856 13197
rect 897 13180 922 13197
rect 984 13197 1013 13214
rect 1047 13197 1076 13214
rect 984 13180 1009 13197
rect 1050 13180 1076 13197
rect 1348 13190 1880 13244
rect 2627 13197 3073 13251
rect 556 13152 566 13174
rect 607 13152 616 13174
rect 556 13134 616 13152
rect 702 13152 710 13174
rect 751 13152 762 13174
rect 702 13134 762 13152
rect 846 13157 856 13180
rect 897 13157 906 13180
rect 846 13140 906 13157
rect 1000 13157 1009 13180
rect 1050 13157 1060 13180
rect 1000 13140 1060 13157
rect 1410 13109 1444 13128
rect 1410 13041 1444 13043
rect 1410 13005 1444 13007
rect 1410 12920 1444 12939
rect 1568 13109 1602 13128
rect 1568 13041 1602 13043
rect 1568 13005 1602 13007
rect 1568 12920 1602 12939
rect 1698 13109 1732 13128
rect 1698 13041 1732 13043
rect 1698 13005 1732 13007
rect 1698 12920 1732 12939
rect 1856 13109 1890 13128
rect 1856 13041 1890 13043
rect 1856 13005 1890 13007
rect 1856 12920 1890 12939
rect 2030 13109 2064 13128
rect 2030 13041 2064 13043
rect 2030 13005 2064 13007
rect 2030 12920 2064 12939
rect 2188 13109 2222 13128
rect 2188 13041 2222 13043
rect 2188 13005 2222 13007
rect 2188 12920 2222 12939
rect 2372 13109 2406 13128
rect 2372 13041 2406 13043
rect 2372 13005 2406 13007
rect 2372 12920 2406 12939
rect 2530 13109 2564 13128
rect 2627 13047 2681 13197
rect 2776 13109 2810 13128
rect 2530 13041 2564 13043
rect 2530 13005 2564 13007
rect 2530 12920 2564 12939
rect 2625 13025 2703 13047
rect 2625 12991 2647 13025
rect 2681 12991 2703 13025
rect 1255 12890 1318 12902
rect 1251 12871 1322 12890
rect 2625 12887 2703 12991
rect 2776 13041 2810 13043
rect 2776 13005 2810 13007
rect 2776 12920 2810 12939
rect 2934 13109 2968 13128
rect 2934 13041 2968 13043
rect 2934 13005 2968 13007
rect 2934 12920 2968 12939
rect 1773 12878 1807 12887
rect 2271 12881 2309 12887
rect 1251 12837 1269 12871
rect 1303 12837 1322 12871
rect 1251 12819 1322 12837
rect 1766 12871 1814 12878
rect 1766 12837 1773 12871
rect 1807 12837 1814 12871
rect 1766 12830 1814 12837
rect 2261 12869 2319 12881
rect 2261 12835 2273 12869
rect 2307 12835 2319 12869
rect 2615 12879 2713 12887
rect 2615 12845 2647 12879
rect 2681 12845 2713 12879
rect 2857 12874 2891 12883
rect 2615 12838 2713 12845
rect 2850 12867 2898 12874
rect 3019 12867 3073 13197
rect 3724 13243 3773 13277
rect 3831 13243 3841 13277
rect 3903 13243 3909 13277
rect 3975 13243 3977 13277
rect 4011 13243 4013 13277
rect 4079 13243 4085 13277
rect 4147 13243 4157 13277
rect 4215 13243 4264 13277
rect 3724 13190 4264 13243
rect 5682 13276 6222 13330
rect 5682 13242 5732 13276
rect 5790 13242 5800 13276
rect 5862 13242 5868 13276
rect 5934 13242 5936 13276
rect 5970 13242 5972 13276
rect 6038 13242 6044 13276
rect 6106 13242 6116 13276
rect 6174 13242 6222 13276
rect 5682 13190 6222 13242
rect 3120 13109 3154 13128
rect 3120 13041 3154 13043
rect 3120 13005 3154 13007
rect 3120 12920 3154 12939
rect 3278 13109 3312 13128
rect 3278 13041 3312 13043
rect 3278 13005 3312 13007
rect 3278 12920 3312 12939
rect 3742 13119 3776 13138
rect 3742 13051 3776 13053
rect 3742 13015 3776 13017
rect 3742 12930 3776 12949
rect 3900 13119 3934 13138
rect 3900 13051 3934 13053
rect 3900 13015 3934 13017
rect 3900 12930 3934 12949
rect 4050 13119 4084 13138
rect 4050 13051 4084 13053
rect 4050 13015 4084 13017
rect 4050 12930 4084 12949
rect 4208 13119 4242 13138
rect 4208 13051 4242 13053
rect 4208 13015 4242 13017
rect 4208 12930 4242 12949
rect 4402 13119 4436 13138
rect 4402 13051 4436 13053
rect 4402 13015 4436 13017
rect 4402 12930 4436 12949
rect 4560 13119 4594 13138
rect 4560 13051 4594 13053
rect 4560 13015 4594 13017
rect 4560 12930 4594 12949
rect 4710 13119 4744 13138
rect 4710 13051 4744 13053
rect 4710 13015 4744 13017
rect 4710 12930 4744 12949
rect 4868 13119 4902 13138
rect 4868 13051 4902 13053
rect 4868 13015 4902 13017
rect 4868 12930 4902 12949
rect 5700 13120 5734 13138
rect 5700 13052 5734 13054
rect 5700 13016 5734 13018
rect 5700 12930 5734 12950
rect 5858 13120 5892 13138
rect 5858 13052 5892 13054
rect 5858 13016 5892 13018
rect 5858 12930 5892 12950
rect 6008 13120 6042 13138
rect 6008 13052 6042 13054
rect 6008 13016 6042 13018
rect 6008 12930 6042 12950
rect 6166 13120 6200 13138
rect 6166 13052 6200 13054
rect 6166 13016 6200 13018
rect 6166 12930 6200 12950
rect 6360 13120 6394 13138
rect 6360 13052 6394 13054
rect 6360 13016 6394 13018
rect 6360 12930 6394 12950
rect 6518 13120 6552 13138
rect 6518 13052 6552 13054
rect 6518 13016 6552 13018
rect 6518 12930 6552 12950
rect 6668 13120 6702 13138
rect 6668 13052 6702 13054
rect 6668 13016 6702 13018
rect 6668 12930 6702 12950
rect 6826 13120 6860 13138
rect 6826 13052 6860 13054
rect 6826 13016 6860 13018
rect 6826 12930 6860 12950
rect 3670 12894 3704 12907
rect 3668 12891 3707 12894
rect 1773 12821 1807 12830
rect 2261 12823 2319 12835
rect 2625 12824 2703 12838
rect 2850 12833 2857 12867
rect 2891 12833 2898 12867
rect 3013 12833 3029 12867
rect 3063 12833 3079 12867
rect 3668 12857 3670 12891
rect 3704 12857 3707 12891
rect 3984 12885 4018 12898
rect 5628 12894 5662 12908
rect 3668 12855 3707 12857
rect 3982 12882 4021 12885
rect 3670 12841 3704 12855
rect 3982 12848 3984 12882
rect 4018 12848 4021 12882
rect 3982 12846 4021 12848
rect 4306 12877 4340 12892
rect 4306 12876 4341 12877
rect 2850 12826 2898 12833
rect 1255 12807 1318 12819
rect 2271 12817 2309 12823
rect 1410 12753 1444 12790
rect 556 12664 616 12680
rect 556 12640 565 12664
rect 606 12640 616 12664
rect 702 12664 762 12680
rect 702 12640 712 12664
rect 753 12640 762 12664
rect 846 12669 906 12686
rect 846 12646 856 12669
rect 897 12646 906 12669
rect 1000 12670 1060 12686
rect 1410 12682 1444 12719
rect 1568 12753 1602 12790
rect 1568 12682 1602 12719
rect 1698 12753 1732 12790
rect 1698 12682 1732 12719
rect 1856 12753 1890 12790
rect 1856 12682 1890 12719
rect 2030 12753 2064 12790
rect 2030 12682 2064 12719
rect 2188 12753 2222 12790
rect 2188 12682 2222 12719
rect 2352 12753 2420 12796
rect 2352 12719 2372 12753
rect 2406 12719 2420 12753
rect 1000 12646 1010 12670
rect 1051 12646 1060 12670
rect 540 12624 565 12640
rect 606 12624 632 12640
rect 540 12606 569 12624
rect 603 12606 632 12624
rect 686 12624 712 12640
rect 753 12624 778 12640
rect 686 12606 715 12624
rect 749 12606 778 12624
rect 830 12629 856 12646
rect 897 12629 922 12646
rect 830 12612 859 12629
rect 893 12612 922 12629
rect 984 12630 1010 12646
rect 1051 12630 1076 12646
rect 984 12612 1013 12630
rect 1047 12612 1076 12630
rect 1324 12576 1960 12640
rect 1324 12542 1353 12576
rect 1407 12542 1421 12576
rect 1479 12542 1489 12576
rect 1551 12542 1557 12576
rect 1623 12542 1625 12576
rect 1659 12542 1661 12576
rect 1727 12542 1733 12576
rect 1795 12542 1805 12576
rect 1863 12542 1877 12576
rect 1931 12542 1960 12576
rect 1324 12500 1960 12542
rect 2352 12551 2420 12719
rect 2530 12753 2564 12790
rect 2530 12682 2564 12719
rect 2352 12517 2369 12551
rect 2403 12517 2420 12551
rect 2352 12500 2420 12517
rect 2642 12455 2696 12824
rect 2857 12817 2891 12826
rect 3019 12823 3073 12833
rect 3984 12832 4018 12846
rect 4340 12842 4341 12876
rect 4621 12860 4637 12894
rect 4671 12860 4687 12894
rect 5626 12892 5666 12894
rect 5626 12858 5628 12892
rect 5662 12858 5666 12892
rect 5942 12886 5976 12898
rect 5626 12856 5666 12858
rect 5940 12882 5980 12886
rect 5628 12842 5662 12856
rect 5940 12848 5942 12882
rect 5976 12848 5980 12882
rect 5940 12846 5980 12848
rect 6264 12878 6298 12892
rect 6264 12876 6300 12878
rect 4306 12826 4340 12842
rect 5942 12832 5976 12846
rect 6298 12842 6300 12876
rect 6580 12860 6596 12894
rect 6630 12860 6646 12894
rect 6264 12826 6298 12842
rect 2776 12753 2810 12790
rect 2776 12682 2810 12719
rect 2934 12753 2968 12790
rect 2934 12682 2968 12719
rect 3120 12753 3154 12790
rect 3120 12682 3154 12719
rect 3278 12753 3312 12790
rect 3278 12682 3312 12719
rect 3742 12763 3776 12800
rect 3742 12692 3776 12729
rect 3900 12763 3934 12800
rect 3900 12692 3934 12729
rect 4050 12763 4084 12800
rect 4050 12692 4084 12729
rect 4208 12763 4242 12800
rect 4208 12692 4242 12729
rect 4402 12765 4436 12802
rect 4402 12694 4436 12731
rect 4560 12765 4594 12802
rect 4560 12694 4594 12731
rect 4710 12765 4744 12802
rect 4710 12694 4744 12731
rect 4868 12765 4902 12802
rect 4868 12694 4902 12731
rect 5700 12764 5734 12800
rect 5700 12692 5734 12730
rect 5858 12764 5892 12800
rect 5858 12692 5892 12730
rect 6008 12764 6042 12800
rect 6008 12692 6042 12730
rect 6166 12764 6200 12800
rect 6166 12692 6200 12730
rect 6360 12766 6394 12802
rect 6360 12694 6394 12732
rect 6518 12766 6552 12802
rect 6518 12694 6552 12732
rect 6668 12766 6702 12802
rect 6668 12694 6702 12732
rect 6826 12766 6860 12802
rect 6826 12694 6860 12732
rect 3704 12587 4244 12640
rect 3704 12553 3741 12587
rect 3787 12553 3813 12587
rect 3855 12553 3885 12587
rect 3923 12553 3957 12587
rect 3991 12553 4025 12587
rect 4063 12553 4093 12587
rect 4135 12553 4161 12587
rect 4207 12553 4244 12587
rect 3704 12500 4244 12553
rect 5662 12588 6202 12640
rect 5662 12554 5700 12588
rect 5746 12554 5772 12588
rect 5814 12554 5844 12588
rect 5882 12554 5916 12588
rect 5950 12554 5984 12588
rect 6022 12554 6052 12588
rect 6094 12554 6120 12588
rect 6166 12554 6202 12588
rect 5662 12500 6202 12554
rect 1348 12050 1880 12102
rect 1348 12016 1383 12050
rect 1429 12016 1455 12050
rect 1497 12016 1527 12050
rect 1565 12016 1599 12050
rect 1633 12016 1667 12050
rect 1705 12016 1735 12050
rect 1777 12016 1803 12050
rect 1849 12016 1880 12050
rect 3724 12049 4264 12102
rect 540 11964 569 11980
rect 603 11964 632 11980
rect 540 11946 566 11964
rect 607 11946 632 11964
rect 686 11964 715 11980
rect 749 11964 778 11980
rect 686 11946 710 11964
rect 751 11946 778 11964
rect 830 11969 859 11986
rect 893 11969 922 11986
rect 830 11952 856 11969
rect 897 11952 922 11969
rect 984 11969 1013 11986
rect 1047 11969 1076 11986
rect 984 11952 1009 11969
rect 1050 11952 1076 11969
rect 1348 11962 1880 12016
rect 2627 11969 3073 12023
rect 556 11924 566 11946
rect 607 11924 616 11946
rect 556 11906 616 11924
rect 702 11924 710 11946
rect 751 11924 762 11946
rect 702 11906 762 11924
rect 846 11929 856 11952
rect 897 11929 906 11952
rect 846 11912 906 11929
rect 1000 11929 1009 11952
rect 1050 11929 1060 11952
rect 1000 11912 1060 11929
rect 1410 11881 1444 11900
rect 1410 11813 1444 11815
rect 1410 11777 1444 11779
rect 1410 11692 1444 11711
rect 1568 11881 1602 11900
rect 1568 11813 1602 11815
rect 1568 11777 1602 11779
rect 1568 11692 1602 11711
rect 1698 11881 1732 11900
rect 1698 11813 1732 11815
rect 1698 11777 1732 11779
rect 1698 11692 1732 11711
rect 1856 11881 1890 11900
rect 1856 11813 1890 11815
rect 1856 11777 1890 11779
rect 1856 11692 1890 11711
rect 2030 11881 2064 11900
rect 2030 11813 2064 11815
rect 2030 11777 2064 11779
rect 2030 11692 2064 11711
rect 2188 11881 2222 11900
rect 2188 11813 2222 11815
rect 2188 11777 2222 11779
rect 2188 11692 2222 11711
rect 2372 11881 2406 11900
rect 2372 11813 2406 11815
rect 2372 11777 2406 11779
rect 2372 11692 2406 11711
rect 2530 11881 2564 11900
rect 2627 11819 2681 11969
rect 2776 11881 2810 11900
rect 2530 11813 2564 11815
rect 2530 11777 2564 11779
rect 2530 11692 2564 11711
rect 2625 11797 2703 11819
rect 2625 11763 2647 11797
rect 2681 11763 2703 11797
rect 1255 11662 1318 11674
rect 1251 11643 1322 11662
rect 2625 11659 2703 11763
rect 2776 11813 2810 11815
rect 2776 11777 2810 11779
rect 2776 11692 2810 11711
rect 2934 11881 2968 11900
rect 2934 11813 2968 11815
rect 2934 11777 2968 11779
rect 2934 11692 2968 11711
rect 1773 11650 1807 11659
rect 2271 11653 2309 11659
rect 1251 11609 1269 11643
rect 1303 11609 1322 11643
rect 1251 11591 1322 11609
rect 1766 11643 1814 11650
rect 1766 11609 1773 11643
rect 1807 11609 1814 11643
rect 1766 11602 1814 11609
rect 2261 11641 2319 11653
rect 2261 11607 2273 11641
rect 2307 11607 2319 11641
rect 2615 11651 2713 11659
rect 2615 11617 2647 11651
rect 2681 11617 2713 11651
rect 2857 11646 2891 11655
rect 2615 11610 2713 11617
rect 2850 11639 2898 11646
rect 3019 11639 3073 11969
rect 3724 12015 3773 12049
rect 3831 12015 3841 12049
rect 3903 12015 3909 12049
rect 3975 12015 3977 12049
rect 4011 12015 4013 12049
rect 4079 12015 4085 12049
rect 4147 12015 4157 12049
rect 4215 12015 4264 12049
rect 3724 11962 4264 12015
rect 5682 12048 6222 12102
rect 5682 12014 5732 12048
rect 5790 12014 5800 12048
rect 5862 12014 5868 12048
rect 5934 12014 5936 12048
rect 5970 12014 5972 12048
rect 6038 12014 6044 12048
rect 6106 12014 6116 12048
rect 6174 12014 6222 12048
rect 5682 11962 6222 12014
rect 3120 11881 3154 11900
rect 3120 11813 3154 11815
rect 3120 11777 3154 11779
rect 3120 11692 3154 11711
rect 3278 11881 3312 11900
rect 3278 11813 3312 11815
rect 3278 11777 3312 11779
rect 3278 11692 3312 11711
rect 3742 11891 3776 11910
rect 3742 11823 3776 11825
rect 3742 11787 3776 11789
rect 3742 11702 3776 11721
rect 3900 11891 3934 11910
rect 3900 11823 3934 11825
rect 3900 11787 3934 11789
rect 3900 11702 3934 11721
rect 4050 11891 4084 11910
rect 4050 11823 4084 11825
rect 4050 11787 4084 11789
rect 4050 11702 4084 11721
rect 4208 11891 4242 11910
rect 4208 11823 4242 11825
rect 4208 11787 4242 11789
rect 4208 11702 4242 11721
rect 4402 11891 4436 11910
rect 4402 11823 4436 11825
rect 4402 11787 4436 11789
rect 4402 11702 4436 11721
rect 4560 11891 4594 11910
rect 4560 11823 4594 11825
rect 4560 11787 4594 11789
rect 4560 11702 4594 11721
rect 4710 11891 4744 11910
rect 4710 11823 4744 11825
rect 4710 11787 4744 11789
rect 4710 11702 4744 11721
rect 4868 11891 4902 11910
rect 4868 11823 4902 11825
rect 4868 11787 4902 11789
rect 4868 11702 4902 11721
rect 5700 11892 5734 11910
rect 5700 11824 5734 11826
rect 5700 11788 5734 11790
rect 5700 11702 5734 11722
rect 5858 11892 5892 11910
rect 5858 11824 5892 11826
rect 5858 11788 5892 11790
rect 5858 11702 5892 11722
rect 6008 11892 6042 11910
rect 6008 11824 6042 11826
rect 6008 11788 6042 11790
rect 6008 11702 6042 11722
rect 6166 11892 6200 11910
rect 6166 11824 6200 11826
rect 6166 11788 6200 11790
rect 6166 11702 6200 11722
rect 6360 11892 6394 11910
rect 6360 11824 6394 11826
rect 6360 11788 6394 11790
rect 6360 11702 6394 11722
rect 6518 11892 6552 11910
rect 6518 11824 6552 11826
rect 6518 11788 6552 11790
rect 6518 11702 6552 11722
rect 6668 11892 6702 11910
rect 6668 11824 6702 11826
rect 6668 11788 6702 11790
rect 6668 11702 6702 11722
rect 6826 11892 6860 11910
rect 6826 11824 6860 11826
rect 6826 11788 6860 11790
rect 6826 11702 6860 11722
rect 3670 11666 3704 11679
rect 3668 11663 3707 11666
rect 1773 11593 1807 11602
rect 2261 11595 2319 11607
rect 2625 11596 2703 11610
rect 2850 11605 2857 11639
rect 2891 11605 2898 11639
rect 3013 11605 3029 11639
rect 3063 11605 3079 11639
rect 3668 11629 3670 11663
rect 3704 11629 3707 11663
rect 3984 11657 4018 11670
rect 5628 11666 5662 11680
rect 3668 11627 3707 11629
rect 3982 11654 4021 11657
rect 3670 11613 3704 11627
rect 3982 11620 3984 11654
rect 4018 11620 4021 11654
rect 3982 11618 4021 11620
rect 4306 11649 4340 11664
rect 4306 11648 4341 11649
rect 2850 11598 2898 11605
rect 1255 11579 1318 11591
rect 2271 11589 2309 11595
rect 1410 11525 1444 11562
rect 556 11436 616 11452
rect 556 11412 565 11436
rect 606 11412 616 11436
rect 702 11436 762 11452
rect 702 11412 712 11436
rect 753 11412 762 11436
rect 846 11441 906 11458
rect 846 11418 856 11441
rect 897 11418 906 11441
rect 1000 11442 1060 11458
rect 1410 11454 1444 11491
rect 1568 11525 1602 11562
rect 1568 11454 1602 11491
rect 1698 11525 1732 11562
rect 1698 11454 1732 11491
rect 1856 11525 1890 11562
rect 1856 11454 1890 11491
rect 2030 11525 2064 11562
rect 2030 11454 2064 11491
rect 2188 11525 2222 11562
rect 2188 11454 2222 11491
rect 2352 11525 2420 11568
rect 2352 11491 2372 11525
rect 2406 11491 2420 11525
rect 1000 11418 1010 11442
rect 1051 11418 1060 11442
rect 540 11396 565 11412
rect 606 11396 632 11412
rect 540 11378 569 11396
rect 603 11378 632 11396
rect 686 11396 712 11412
rect 753 11396 778 11412
rect 686 11378 715 11396
rect 749 11378 778 11396
rect 830 11401 856 11418
rect 897 11401 922 11418
rect 830 11384 859 11401
rect 893 11384 922 11401
rect 984 11402 1010 11418
rect 1051 11402 1076 11418
rect 984 11384 1013 11402
rect 1047 11384 1076 11402
rect 1324 11348 1960 11412
rect 1324 11314 1353 11348
rect 1407 11314 1421 11348
rect 1479 11314 1489 11348
rect 1551 11314 1557 11348
rect 1623 11314 1625 11348
rect 1659 11314 1661 11348
rect 1727 11314 1733 11348
rect 1795 11314 1805 11348
rect 1863 11314 1877 11348
rect 1931 11314 1960 11348
rect 1324 11272 1960 11314
rect 2352 11323 2420 11491
rect 2530 11525 2564 11562
rect 2530 11454 2564 11491
rect 2352 11289 2369 11323
rect 2403 11289 2420 11323
rect 2352 11272 2420 11289
rect 2642 11227 2696 11596
rect 2857 11589 2891 11598
rect 3019 11595 3073 11605
rect 3984 11604 4018 11618
rect 4340 11614 4341 11648
rect 4621 11632 4637 11666
rect 4671 11632 4687 11666
rect 5626 11664 5666 11666
rect 5626 11630 5628 11664
rect 5662 11630 5666 11664
rect 5942 11658 5976 11670
rect 5626 11628 5666 11630
rect 5940 11654 5980 11658
rect 5628 11614 5662 11628
rect 5940 11620 5942 11654
rect 5976 11620 5980 11654
rect 5940 11618 5980 11620
rect 6264 11650 6298 11664
rect 6264 11648 6300 11650
rect 4306 11598 4340 11614
rect 5942 11604 5976 11618
rect 6298 11614 6300 11648
rect 6580 11632 6596 11666
rect 6630 11632 6646 11666
rect 6264 11598 6298 11614
rect 2776 11525 2810 11562
rect 2776 11454 2810 11491
rect 2934 11525 2968 11562
rect 2934 11454 2968 11491
rect 3120 11525 3154 11562
rect 3120 11454 3154 11491
rect 3278 11525 3312 11562
rect 3278 11454 3312 11491
rect 3742 11535 3776 11572
rect 3742 11464 3776 11501
rect 3900 11535 3934 11572
rect 3900 11464 3934 11501
rect 4050 11535 4084 11572
rect 4050 11464 4084 11501
rect 4208 11535 4242 11572
rect 4208 11464 4242 11501
rect 4402 11537 4436 11574
rect 4402 11466 4436 11503
rect 4560 11537 4594 11574
rect 4560 11466 4594 11503
rect 4710 11537 4744 11574
rect 4710 11466 4744 11503
rect 4868 11537 4902 11574
rect 4868 11466 4902 11503
rect 5700 11536 5734 11572
rect 5700 11464 5734 11502
rect 5858 11536 5892 11572
rect 5858 11464 5892 11502
rect 6008 11536 6042 11572
rect 6008 11464 6042 11502
rect 6166 11536 6200 11572
rect 6166 11464 6200 11502
rect 6360 11538 6394 11574
rect 6360 11466 6394 11504
rect 6518 11538 6552 11574
rect 6518 11466 6552 11504
rect 6668 11538 6702 11574
rect 6668 11466 6702 11504
rect 6826 11538 6860 11574
rect 6826 11466 6860 11504
rect 3704 11359 4244 11412
rect 3704 11325 3741 11359
rect 3787 11325 3813 11359
rect 3855 11325 3885 11359
rect 3923 11325 3957 11359
rect 3991 11325 4025 11359
rect 4063 11325 4093 11359
rect 4135 11325 4161 11359
rect 4207 11325 4244 11359
rect 3704 11272 4244 11325
rect 5662 11360 6202 11412
rect 5662 11326 5700 11360
rect 5746 11326 5772 11360
rect 5814 11326 5844 11360
rect 5882 11326 5916 11360
rect 5950 11326 5984 11360
rect 6022 11326 6052 11360
rect 6094 11326 6120 11360
rect 6166 11326 6202 11360
rect 5662 11272 6202 11326
rect 1348 10822 1880 10874
rect 1348 10788 1383 10822
rect 1429 10788 1455 10822
rect 1497 10788 1527 10822
rect 1565 10788 1599 10822
rect 1633 10788 1667 10822
rect 1705 10788 1735 10822
rect 1777 10788 1803 10822
rect 1849 10788 1880 10822
rect 3724 10821 4264 10874
rect 540 10736 569 10752
rect 603 10736 632 10752
rect 540 10718 566 10736
rect 607 10718 632 10736
rect 686 10736 715 10752
rect 749 10736 778 10752
rect 686 10718 710 10736
rect 751 10718 778 10736
rect 830 10741 859 10758
rect 893 10741 922 10758
rect 830 10724 856 10741
rect 897 10724 922 10741
rect 984 10741 1013 10758
rect 1047 10741 1076 10758
rect 984 10724 1009 10741
rect 1050 10724 1076 10741
rect 1348 10734 1880 10788
rect 2627 10741 3073 10795
rect 556 10696 566 10718
rect 607 10696 616 10718
rect 556 10678 616 10696
rect 702 10696 710 10718
rect 751 10696 762 10718
rect 702 10678 762 10696
rect 846 10701 856 10724
rect 897 10701 906 10724
rect 846 10684 906 10701
rect 1000 10701 1009 10724
rect 1050 10701 1060 10724
rect 1000 10684 1060 10701
rect 1410 10653 1444 10672
rect 1410 10585 1444 10587
rect 1410 10549 1444 10551
rect 1410 10464 1444 10483
rect 1568 10653 1602 10672
rect 1568 10585 1602 10587
rect 1568 10549 1602 10551
rect 1568 10464 1602 10483
rect 1698 10653 1732 10672
rect 1698 10585 1732 10587
rect 1698 10549 1732 10551
rect 1698 10464 1732 10483
rect 1856 10653 1890 10672
rect 1856 10585 1890 10587
rect 1856 10549 1890 10551
rect 1856 10464 1890 10483
rect 2030 10653 2064 10672
rect 2030 10585 2064 10587
rect 2030 10549 2064 10551
rect 2030 10464 2064 10483
rect 2188 10653 2222 10672
rect 2188 10585 2222 10587
rect 2188 10549 2222 10551
rect 2188 10464 2222 10483
rect 2372 10653 2406 10672
rect 2372 10585 2406 10587
rect 2372 10549 2406 10551
rect 2372 10464 2406 10483
rect 2530 10653 2564 10672
rect 2627 10591 2681 10741
rect 2776 10653 2810 10672
rect 2530 10585 2564 10587
rect 2530 10549 2564 10551
rect 2530 10464 2564 10483
rect 2625 10569 2703 10591
rect 2625 10535 2647 10569
rect 2681 10535 2703 10569
rect 1255 10434 1318 10446
rect 1251 10415 1322 10434
rect 2625 10431 2703 10535
rect 2776 10585 2810 10587
rect 2776 10549 2810 10551
rect 2776 10464 2810 10483
rect 2934 10653 2968 10672
rect 2934 10585 2968 10587
rect 2934 10549 2968 10551
rect 2934 10464 2968 10483
rect 1773 10422 1807 10431
rect 2271 10425 2309 10431
rect 1251 10381 1269 10415
rect 1303 10381 1322 10415
rect 1251 10363 1322 10381
rect 1766 10415 1814 10422
rect 1766 10381 1773 10415
rect 1807 10381 1814 10415
rect 1766 10374 1814 10381
rect 2261 10413 2319 10425
rect 2261 10379 2273 10413
rect 2307 10379 2319 10413
rect 2615 10423 2713 10431
rect 2615 10389 2647 10423
rect 2681 10389 2713 10423
rect 2857 10418 2891 10427
rect 2615 10382 2713 10389
rect 2850 10411 2898 10418
rect 3019 10411 3073 10741
rect 3724 10787 3773 10821
rect 3831 10787 3841 10821
rect 3903 10787 3909 10821
rect 3975 10787 3977 10821
rect 4011 10787 4013 10821
rect 4079 10787 4085 10821
rect 4147 10787 4157 10821
rect 4215 10787 4264 10821
rect 3724 10734 4264 10787
rect 5682 10820 6222 10874
rect 5682 10786 5732 10820
rect 5790 10786 5800 10820
rect 5862 10786 5868 10820
rect 5934 10786 5936 10820
rect 5970 10786 5972 10820
rect 6038 10786 6044 10820
rect 6106 10786 6116 10820
rect 6174 10786 6222 10820
rect 5682 10734 6222 10786
rect 3120 10653 3154 10672
rect 3120 10585 3154 10587
rect 3120 10549 3154 10551
rect 3120 10464 3154 10483
rect 3278 10653 3312 10672
rect 3278 10585 3312 10587
rect 3278 10549 3312 10551
rect 3278 10464 3312 10483
rect 3742 10663 3776 10682
rect 3742 10595 3776 10597
rect 3742 10559 3776 10561
rect 3742 10474 3776 10493
rect 3900 10663 3934 10682
rect 3900 10595 3934 10597
rect 3900 10559 3934 10561
rect 3900 10474 3934 10493
rect 4050 10663 4084 10682
rect 4050 10595 4084 10597
rect 4050 10559 4084 10561
rect 4050 10474 4084 10493
rect 4208 10663 4242 10682
rect 4208 10595 4242 10597
rect 4208 10559 4242 10561
rect 4208 10474 4242 10493
rect 4402 10663 4436 10682
rect 4402 10595 4436 10597
rect 4402 10559 4436 10561
rect 4402 10474 4436 10493
rect 4560 10663 4594 10682
rect 4560 10595 4594 10597
rect 4560 10559 4594 10561
rect 4560 10474 4594 10493
rect 4710 10663 4744 10682
rect 4710 10595 4744 10597
rect 4710 10559 4744 10561
rect 4710 10474 4744 10493
rect 4868 10663 4902 10682
rect 4868 10595 4902 10597
rect 4868 10559 4902 10561
rect 4868 10474 4902 10493
rect 5700 10664 5734 10682
rect 5700 10596 5734 10598
rect 5700 10560 5734 10562
rect 5700 10474 5734 10494
rect 5858 10664 5892 10682
rect 5858 10596 5892 10598
rect 5858 10560 5892 10562
rect 5858 10474 5892 10494
rect 6008 10664 6042 10682
rect 6008 10596 6042 10598
rect 6008 10560 6042 10562
rect 6008 10474 6042 10494
rect 6166 10664 6200 10682
rect 6166 10596 6200 10598
rect 6166 10560 6200 10562
rect 6166 10474 6200 10494
rect 6360 10664 6394 10682
rect 6360 10596 6394 10598
rect 6360 10560 6394 10562
rect 6360 10474 6394 10494
rect 6518 10664 6552 10682
rect 6518 10596 6552 10598
rect 6518 10560 6552 10562
rect 6518 10474 6552 10494
rect 6668 10664 6702 10682
rect 6668 10596 6702 10598
rect 6668 10560 6702 10562
rect 6668 10474 6702 10494
rect 6826 10664 6860 10682
rect 6826 10596 6860 10598
rect 6826 10560 6860 10562
rect 6826 10474 6860 10494
rect 3670 10438 3704 10451
rect 3668 10435 3707 10438
rect 1773 10365 1807 10374
rect 2261 10367 2319 10379
rect 2625 10368 2703 10382
rect 2850 10377 2857 10411
rect 2891 10377 2898 10411
rect 3013 10377 3029 10411
rect 3063 10377 3079 10411
rect 3668 10401 3670 10435
rect 3704 10401 3707 10435
rect 3984 10429 4018 10442
rect 5628 10438 5662 10452
rect 3668 10399 3707 10401
rect 3982 10426 4021 10429
rect 3670 10385 3704 10399
rect 3982 10392 3984 10426
rect 4018 10392 4021 10426
rect 3982 10390 4021 10392
rect 4306 10421 4340 10436
rect 4306 10420 4341 10421
rect 2850 10370 2898 10377
rect 1255 10351 1318 10363
rect 2271 10361 2309 10367
rect 1410 10297 1444 10334
rect 556 10208 616 10224
rect 556 10184 565 10208
rect 606 10184 616 10208
rect 702 10208 762 10224
rect 702 10184 712 10208
rect 753 10184 762 10208
rect 846 10213 906 10230
rect 846 10190 856 10213
rect 897 10190 906 10213
rect 1000 10214 1060 10230
rect 1410 10226 1444 10263
rect 1568 10297 1602 10334
rect 1568 10226 1602 10263
rect 1698 10297 1732 10334
rect 1698 10226 1732 10263
rect 1856 10297 1890 10334
rect 1856 10226 1890 10263
rect 2030 10297 2064 10334
rect 2030 10226 2064 10263
rect 2188 10297 2222 10334
rect 2188 10226 2222 10263
rect 2352 10297 2420 10340
rect 2352 10263 2372 10297
rect 2406 10263 2420 10297
rect 1000 10190 1010 10214
rect 1051 10190 1060 10214
rect 540 10168 565 10184
rect 606 10168 632 10184
rect 540 10150 569 10168
rect 603 10150 632 10168
rect 686 10168 712 10184
rect 753 10168 778 10184
rect 686 10150 715 10168
rect 749 10150 778 10168
rect 830 10173 856 10190
rect 897 10173 922 10190
rect 830 10156 859 10173
rect 893 10156 922 10173
rect 984 10174 1010 10190
rect 1051 10174 1076 10190
rect 984 10156 1013 10174
rect 1047 10156 1076 10174
rect 1324 10120 1960 10184
rect 1324 10086 1353 10120
rect 1407 10086 1421 10120
rect 1479 10086 1489 10120
rect 1551 10086 1557 10120
rect 1623 10086 1625 10120
rect 1659 10086 1661 10120
rect 1727 10086 1733 10120
rect 1795 10086 1805 10120
rect 1863 10086 1877 10120
rect 1931 10086 1960 10120
rect 1324 10044 1960 10086
rect 2352 10095 2420 10263
rect 2530 10297 2564 10334
rect 2530 10226 2564 10263
rect 2352 10061 2369 10095
rect 2403 10061 2420 10095
rect 2352 10044 2420 10061
rect 2642 9999 2696 10368
rect 2857 10361 2891 10370
rect 3019 10367 3073 10377
rect 3984 10376 4018 10390
rect 4340 10386 4341 10420
rect 4621 10404 4637 10438
rect 4671 10404 4687 10438
rect 5626 10436 5666 10438
rect 5626 10402 5628 10436
rect 5662 10402 5666 10436
rect 5942 10430 5976 10442
rect 5626 10400 5666 10402
rect 5940 10426 5980 10430
rect 5628 10386 5662 10400
rect 5940 10392 5942 10426
rect 5976 10392 5980 10426
rect 5940 10390 5980 10392
rect 6264 10422 6298 10436
rect 6264 10420 6300 10422
rect 4306 10370 4340 10386
rect 5942 10376 5976 10390
rect 6298 10386 6300 10420
rect 6580 10404 6596 10438
rect 6630 10404 6646 10438
rect 6264 10370 6298 10386
rect 2776 10297 2810 10334
rect 2776 10226 2810 10263
rect 2934 10297 2968 10334
rect 2934 10226 2968 10263
rect 3120 10297 3154 10334
rect 3120 10226 3154 10263
rect 3278 10297 3312 10334
rect 3278 10226 3312 10263
rect 3742 10307 3776 10344
rect 3742 10236 3776 10273
rect 3900 10307 3934 10344
rect 3900 10236 3934 10273
rect 4050 10307 4084 10344
rect 4050 10236 4084 10273
rect 4208 10307 4242 10344
rect 4208 10236 4242 10273
rect 4402 10309 4436 10346
rect 4402 10238 4436 10275
rect 4560 10309 4594 10346
rect 4560 10238 4594 10275
rect 4710 10309 4744 10346
rect 4710 10238 4744 10275
rect 4868 10309 4902 10346
rect 4868 10238 4902 10275
rect 5700 10308 5734 10344
rect 5700 10236 5734 10274
rect 5858 10308 5892 10344
rect 5858 10236 5892 10274
rect 6008 10308 6042 10344
rect 6008 10236 6042 10274
rect 6166 10308 6200 10344
rect 6166 10236 6200 10274
rect 6360 10310 6394 10346
rect 6360 10238 6394 10276
rect 6518 10310 6552 10346
rect 6518 10238 6552 10276
rect 6668 10310 6702 10346
rect 6668 10238 6702 10276
rect 6826 10310 6860 10346
rect 6826 10238 6860 10276
rect 3704 10131 4244 10184
rect 3704 10097 3741 10131
rect 3787 10097 3813 10131
rect 3855 10097 3885 10131
rect 3923 10097 3957 10131
rect 3991 10097 4025 10131
rect 4063 10097 4093 10131
rect 4135 10097 4161 10131
rect 4207 10097 4244 10131
rect 3704 10044 4244 10097
rect 5662 10132 6202 10184
rect 5662 10098 5700 10132
rect 5746 10098 5772 10132
rect 5814 10098 5844 10132
rect 5882 10098 5916 10132
rect 5950 10098 5984 10132
rect 6022 10098 6052 10132
rect 6094 10098 6120 10132
rect 6166 10098 6202 10132
rect 5662 10044 6202 10098
rect 1348 9594 1880 9646
rect 1348 9560 1383 9594
rect 1429 9560 1455 9594
rect 1497 9560 1527 9594
rect 1565 9560 1599 9594
rect 1633 9560 1667 9594
rect 1705 9560 1735 9594
rect 1777 9560 1803 9594
rect 1849 9560 1880 9594
rect 3724 9593 4264 9646
rect 540 9508 569 9524
rect 603 9508 632 9524
rect 540 9490 566 9508
rect 607 9490 632 9508
rect 686 9508 715 9524
rect 749 9508 778 9524
rect 686 9490 710 9508
rect 751 9490 778 9508
rect 830 9513 859 9530
rect 893 9513 922 9530
rect 830 9496 856 9513
rect 897 9496 922 9513
rect 984 9513 1013 9530
rect 1047 9513 1076 9530
rect 984 9496 1009 9513
rect 1050 9496 1076 9513
rect 1348 9506 1880 9560
rect 2627 9513 3073 9567
rect 556 9468 566 9490
rect 607 9468 616 9490
rect 556 9450 616 9468
rect 702 9468 710 9490
rect 751 9468 762 9490
rect 702 9450 762 9468
rect 846 9473 856 9496
rect 897 9473 906 9496
rect 846 9456 906 9473
rect 1000 9473 1009 9496
rect 1050 9473 1060 9496
rect 1000 9456 1060 9473
rect 1410 9425 1444 9444
rect 1410 9357 1444 9359
rect 1410 9321 1444 9323
rect 1410 9236 1444 9255
rect 1568 9425 1602 9444
rect 1568 9357 1602 9359
rect 1568 9321 1602 9323
rect 1568 9236 1602 9255
rect 1698 9425 1732 9444
rect 1698 9357 1732 9359
rect 1698 9321 1732 9323
rect 1698 9236 1732 9255
rect 1856 9425 1890 9444
rect 1856 9357 1890 9359
rect 1856 9321 1890 9323
rect 1856 9236 1890 9255
rect 2030 9425 2064 9444
rect 2030 9357 2064 9359
rect 2030 9321 2064 9323
rect 2030 9236 2064 9255
rect 2188 9425 2222 9444
rect 2188 9357 2222 9359
rect 2188 9321 2222 9323
rect 2188 9236 2222 9255
rect 2372 9425 2406 9444
rect 2372 9357 2406 9359
rect 2372 9321 2406 9323
rect 2372 9236 2406 9255
rect 2530 9425 2564 9444
rect 2627 9363 2681 9513
rect 2776 9425 2810 9444
rect 2530 9357 2564 9359
rect 2530 9321 2564 9323
rect 2530 9236 2564 9255
rect 2625 9341 2703 9363
rect 2625 9307 2647 9341
rect 2681 9307 2703 9341
rect 1255 9206 1318 9218
rect 1251 9187 1322 9206
rect 2625 9203 2703 9307
rect 2776 9357 2810 9359
rect 2776 9321 2810 9323
rect 2776 9236 2810 9255
rect 2934 9425 2968 9444
rect 2934 9357 2968 9359
rect 2934 9321 2968 9323
rect 2934 9236 2968 9255
rect 1773 9194 1807 9203
rect 2271 9197 2309 9203
rect 1251 9153 1269 9187
rect 1303 9153 1322 9187
rect 1251 9135 1322 9153
rect 1766 9187 1814 9194
rect 1766 9153 1773 9187
rect 1807 9153 1814 9187
rect 1766 9146 1814 9153
rect 2261 9185 2319 9197
rect 2261 9151 2273 9185
rect 2307 9151 2319 9185
rect 2615 9195 2713 9203
rect 2615 9161 2647 9195
rect 2681 9161 2713 9195
rect 2857 9190 2891 9199
rect 2615 9154 2713 9161
rect 2850 9183 2898 9190
rect 3019 9183 3073 9513
rect 3724 9559 3773 9593
rect 3831 9559 3841 9593
rect 3903 9559 3909 9593
rect 3975 9559 3977 9593
rect 4011 9559 4013 9593
rect 4079 9559 4085 9593
rect 4147 9559 4157 9593
rect 4215 9559 4264 9593
rect 3724 9506 4264 9559
rect 5682 9592 6222 9646
rect 5682 9558 5732 9592
rect 5790 9558 5800 9592
rect 5862 9558 5868 9592
rect 5934 9558 5936 9592
rect 5970 9558 5972 9592
rect 6038 9558 6044 9592
rect 6106 9558 6116 9592
rect 6174 9558 6222 9592
rect 5682 9506 6222 9558
rect 3120 9425 3154 9444
rect 3120 9357 3154 9359
rect 3120 9321 3154 9323
rect 3120 9236 3154 9255
rect 3278 9425 3312 9444
rect 3278 9357 3312 9359
rect 3278 9321 3312 9323
rect 3278 9236 3312 9255
rect 3742 9435 3776 9454
rect 3742 9367 3776 9369
rect 3742 9331 3776 9333
rect 3742 9246 3776 9265
rect 3900 9435 3934 9454
rect 3900 9367 3934 9369
rect 3900 9331 3934 9333
rect 3900 9246 3934 9265
rect 4050 9435 4084 9454
rect 4050 9367 4084 9369
rect 4050 9331 4084 9333
rect 4050 9246 4084 9265
rect 4208 9435 4242 9454
rect 4208 9367 4242 9369
rect 4208 9331 4242 9333
rect 4208 9246 4242 9265
rect 4402 9435 4436 9454
rect 4402 9367 4436 9369
rect 4402 9331 4436 9333
rect 4402 9246 4436 9265
rect 4560 9435 4594 9454
rect 4560 9367 4594 9369
rect 4560 9331 4594 9333
rect 4560 9246 4594 9265
rect 4710 9435 4744 9454
rect 4710 9367 4744 9369
rect 4710 9331 4744 9333
rect 4710 9246 4744 9265
rect 4868 9435 4902 9454
rect 4868 9367 4902 9369
rect 4868 9331 4902 9333
rect 4868 9246 4902 9265
rect 5700 9436 5734 9454
rect 5700 9368 5734 9370
rect 5700 9332 5734 9334
rect 5700 9246 5734 9266
rect 5858 9436 5892 9454
rect 5858 9368 5892 9370
rect 5858 9332 5892 9334
rect 5858 9246 5892 9266
rect 6008 9436 6042 9454
rect 6008 9368 6042 9370
rect 6008 9332 6042 9334
rect 6008 9246 6042 9266
rect 6166 9436 6200 9454
rect 6166 9368 6200 9370
rect 6166 9332 6200 9334
rect 6166 9246 6200 9266
rect 6360 9436 6394 9454
rect 6360 9368 6394 9370
rect 6360 9332 6394 9334
rect 6360 9246 6394 9266
rect 6518 9436 6552 9454
rect 6518 9368 6552 9370
rect 6518 9332 6552 9334
rect 6518 9246 6552 9266
rect 6668 9436 6702 9454
rect 6668 9368 6702 9370
rect 6668 9332 6702 9334
rect 6668 9246 6702 9266
rect 6826 9436 6860 9454
rect 6826 9368 6860 9370
rect 6826 9332 6860 9334
rect 6826 9246 6860 9266
rect 3670 9210 3704 9223
rect 3668 9207 3707 9210
rect 1773 9137 1807 9146
rect 2261 9139 2319 9151
rect 2625 9140 2703 9154
rect 2850 9149 2857 9183
rect 2891 9149 2898 9183
rect 3013 9149 3029 9183
rect 3063 9149 3079 9183
rect 3668 9173 3670 9207
rect 3704 9173 3707 9207
rect 3984 9201 4018 9214
rect 5628 9210 5662 9224
rect 3668 9171 3707 9173
rect 3982 9198 4021 9201
rect 3670 9157 3704 9171
rect 3982 9164 3984 9198
rect 4018 9164 4021 9198
rect 3982 9162 4021 9164
rect 4306 9193 4340 9208
rect 4306 9192 4341 9193
rect 2850 9142 2898 9149
rect 1255 9123 1318 9135
rect 2271 9133 2309 9139
rect 1410 9069 1444 9106
rect 556 8980 616 8996
rect 556 8956 565 8980
rect 606 8956 616 8980
rect 702 8980 762 8996
rect 702 8956 712 8980
rect 753 8956 762 8980
rect 846 8985 906 9002
rect 846 8962 856 8985
rect 897 8962 906 8985
rect 1000 8986 1060 9002
rect 1410 8998 1444 9035
rect 1568 9069 1602 9106
rect 1568 8998 1602 9035
rect 1698 9069 1732 9106
rect 1698 8998 1732 9035
rect 1856 9069 1890 9106
rect 1856 8998 1890 9035
rect 2030 9069 2064 9106
rect 2030 8998 2064 9035
rect 2188 9069 2222 9106
rect 2188 8998 2222 9035
rect 2352 9069 2420 9112
rect 2352 9035 2372 9069
rect 2406 9035 2420 9069
rect 1000 8962 1010 8986
rect 1051 8962 1060 8986
rect 540 8940 565 8956
rect 606 8940 632 8956
rect 540 8922 569 8940
rect 603 8922 632 8940
rect 686 8940 712 8956
rect 753 8940 778 8956
rect 686 8922 715 8940
rect 749 8922 778 8940
rect 830 8945 856 8962
rect 897 8945 922 8962
rect 830 8928 859 8945
rect 893 8928 922 8945
rect 984 8946 1010 8962
rect 1051 8946 1076 8962
rect 984 8928 1013 8946
rect 1047 8928 1076 8946
rect 1324 8892 1960 8956
rect 1324 8858 1353 8892
rect 1407 8858 1421 8892
rect 1479 8858 1489 8892
rect 1551 8858 1557 8892
rect 1623 8858 1625 8892
rect 1659 8858 1661 8892
rect 1727 8858 1733 8892
rect 1795 8858 1805 8892
rect 1863 8858 1877 8892
rect 1931 8858 1960 8892
rect 1324 8816 1960 8858
rect 2352 8867 2420 9035
rect 2530 9069 2564 9106
rect 2530 8998 2564 9035
rect 2352 8833 2369 8867
rect 2403 8833 2420 8867
rect 2352 8816 2420 8833
rect 2642 8771 2696 9140
rect 2857 9133 2891 9142
rect 3019 9139 3073 9149
rect 3984 9148 4018 9162
rect 4340 9158 4341 9192
rect 4621 9176 4637 9210
rect 4671 9176 4687 9210
rect 5626 9208 5666 9210
rect 5626 9174 5628 9208
rect 5662 9174 5666 9208
rect 5942 9202 5976 9214
rect 5626 9172 5666 9174
rect 5940 9198 5980 9202
rect 5628 9158 5662 9172
rect 5940 9164 5942 9198
rect 5976 9164 5980 9198
rect 5940 9162 5980 9164
rect 6264 9194 6298 9208
rect 6264 9192 6300 9194
rect 4306 9142 4340 9158
rect 5942 9148 5976 9162
rect 6298 9158 6300 9192
rect 6580 9176 6596 9210
rect 6630 9176 6646 9210
rect 6264 9142 6298 9158
rect 2776 9069 2810 9106
rect 2776 8998 2810 9035
rect 2934 9069 2968 9106
rect 2934 8998 2968 9035
rect 3120 9069 3154 9106
rect 3120 8998 3154 9035
rect 3278 9069 3312 9106
rect 3278 8998 3312 9035
rect 3742 9079 3776 9116
rect 3742 9008 3776 9045
rect 3900 9079 3934 9116
rect 3900 9008 3934 9045
rect 4050 9079 4084 9116
rect 4050 9008 4084 9045
rect 4208 9079 4242 9116
rect 4208 9008 4242 9045
rect 4402 9081 4436 9118
rect 4402 9010 4436 9047
rect 4560 9081 4594 9118
rect 4560 9010 4594 9047
rect 4710 9081 4744 9118
rect 4710 9010 4744 9047
rect 4868 9081 4902 9118
rect 4868 9010 4902 9047
rect 5700 9080 5734 9116
rect 5700 9008 5734 9046
rect 5858 9080 5892 9116
rect 5858 9008 5892 9046
rect 6008 9080 6042 9116
rect 6008 9008 6042 9046
rect 6166 9080 6200 9116
rect 6166 9008 6200 9046
rect 6360 9082 6394 9118
rect 6360 9010 6394 9048
rect 6518 9082 6552 9118
rect 6518 9010 6552 9048
rect 6668 9082 6702 9118
rect 6668 9010 6702 9048
rect 6826 9082 6860 9118
rect 6826 9010 6860 9048
rect 3704 8903 4244 8956
rect 3704 8869 3741 8903
rect 3787 8869 3813 8903
rect 3855 8869 3885 8903
rect 3923 8869 3957 8903
rect 3991 8869 4025 8903
rect 4063 8869 4093 8903
rect 4135 8869 4161 8903
rect 4207 8869 4244 8903
rect 3704 8816 4244 8869
rect 5662 8904 6202 8956
rect 5662 8870 5700 8904
rect 5746 8870 5772 8904
rect 5814 8870 5844 8904
rect 5882 8870 5916 8904
rect 5950 8870 5984 8904
rect 6022 8870 6052 8904
rect 6094 8870 6120 8904
rect 6166 8870 6202 8904
rect 5662 8816 6202 8870
rect 1348 8366 1880 8418
rect 1348 8332 1383 8366
rect 1429 8332 1455 8366
rect 1497 8332 1527 8366
rect 1565 8332 1599 8366
rect 1633 8332 1667 8366
rect 1705 8332 1735 8366
rect 1777 8332 1803 8366
rect 1849 8332 1880 8366
rect 3724 8365 4264 8418
rect 540 8280 569 8296
rect 603 8280 632 8296
rect 540 8262 566 8280
rect 607 8262 632 8280
rect 686 8280 715 8296
rect 749 8280 778 8296
rect 686 8262 710 8280
rect 751 8262 778 8280
rect 830 8285 859 8302
rect 893 8285 922 8302
rect 830 8268 856 8285
rect 897 8268 922 8285
rect 984 8285 1013 8302
rect 1047 8285 1076 8302
rect 984 8268 1009 8285
rect 1050 8268 1076 8285
rect 1348 8278 1880 8332
rect 2627 8285 3073 8339
rect 556 8240 566 8262
rect 607 8240 616 8262
rect 556 8222 616 8240
rect 702 8240 710 8262
rect 751 8240 762 8262
rect 702 8222 762 8240
rect 846 8245 856 8268
rect 897 8245 906 8268
rect 846 8228 906 8245
rect 1000 8245 1009 8268
rect 1050 8245 1060 8268
rect 1000 8228 1060 8245
rect 1410 8197 1444 8216
rect 1410 8129 1444 8131
rect 1410 8093 1444 8095
rect 1410 8008 1444 8027
rect 1568 8197 1602 8216
rect 1568 8129 1602 8131
rect 1568 8093 1602 8095
rect 1568 8008 1602 8027
rect 1698 8197 1732 8216
rect 1698 8129 1732 8131
rect 1698 8093 1732 8095
rect 1698 8008 1732 8027
rect 1856 8197 1890 8216
rect 1856 8129 1890 8131
rect 1856 8093 1890 8095
rect 1856 8008 1890 8027
rect 2030 8197 2064 8216
rect 2030 8129 2064 8131
rect 2030 8093 2064 8095
rect 2030 8008 2064 8027
rect 2188 8197 2222 8216
rect 2188 8129 2222 8131
rect 2188 8093 2222 8095
rect 2188 8008 2222 8027
rect 2372 8197 2406 8216
rect 2372 8129 2406 8131
rect 2372 8093 2406 8095
rect 2372 8008 2406 8027
rect 2530 8197 2564 8216
rect 2627 8135 2681 8285
rect 2776 8197 2810 8216
rect 2530 8129 2564 8131
rect 2530 8093 2564 8095
rect 2530 8008 2564 8027
rect 2625 8113 2703 8135
rect 2625 8079 2647 8113
rect 2681 8079 2703 8113
rect 1255 7978 1318 7990
rect 1251 7959 1322 7978
rect 2625 7975 2703 8079
rect 2776 8129 2810 8131
rect 2776 8093 2810 8095
rect 2776 8008 2810 8027
rect 2934 8197 2968 8216
rect 2934 8129 2968 8131
rect 2934 8093 2968 8095
rect 2934 8008 2968 8027
rect 1773 7966 1807 7975
rect 2271 7969 2309 7975
rect 1251 7925 1269 7959
rect 1303 7925 1322 7959
rect 1251 7907 1322 7925
rect 1766 7959 1814 7966
rect 1766 7925 1773 7959
rect 1807 7925 1814 7959
rect 1766 7918 1814 7925
rect 2261 7957 2319 7969
rect 2261 7923 2273 7957
rect 2307 7923 2319 7957
rect 2615 7967 2713 7975
rect 2615 7933 2647 7967
rect 2681 7933 2713 7967
rect 2857 7962 2891 7971
rect 2615 7926 2713 7933
rect 2850 7955 2898 7962
rect 3019 7955 3073 8285
rect 3724 8331 3773 8365
rect 3831 8331 3841 8365
rect 3903 8331 3909 8365
rect 3975 8331 3977 8365
rect 4011 8331 4013 8365
rect 4079 8331 4085 8365
rect 4147 8331 4157 8365
rect 4215 8331 4264 8365
rect 3724 8278 4264 8331
rect 5682 8364 6222 8418
rect 5682 8330 5732 8364
rect 5790 8330 5800 8364
rect 5862 8330 5868 8364
rect 5934 8330 5936 8364
rect 5970 8330 5972 8364
rect 6038 8330 6044 8364
rect 6106 8330 6116 8364
rect 6174 8330 6222 8364
rect 5682 8278 6222 8330
rect 3120 8197 3154 8216
rect 3120 8129 3154 8131
rect 3120 8093 3154 8095
rect 3120 8008 3154 8027
rect 3278 8197 3312 8216
rect 3278 8129 3312 8131
rect 3278 8093 3312 8095
rect 3278 8008 3312 8027
rect 3742 8207 3776 8226
rect 3742 8139 3776 8141
rect 3742 8103 3776 8105
rect 3742 8018 3776 8037
rect 3900 8207 3934 8226
rect 3900 8139 3934 8141
rect 3900 8103 3934 8105
rect 3900 8018 3934 8037
rect 4050 8207 4084 8226
rect 4050 8139 4084 8141
rect 4050 8103 4084 8105
rect 4050 8018 4084 8037
rect 4208 8207 4242 8226
rect 4208 8139 4242 8141
rect 4208 8103 4242 8105
rect 4208 8018 4242 8037
rect 4402 8207 4436 8226
rect 4402 8139 4436 8141
rect 4402 8103 4436 8105
rect 4402 8018 4436 8037
rect 4560 8207 4594 8226
rect 4560 8139 4594 8141
rect 4560 8103 4594 8105
rect 4560 8018 4594 8037
rect 4710 8207 4744 8226
rect 4710 8139 4744 8141
rect 4710 8103 4744 8105
rect 4710 8018 4744 8037
rect 4868 8207 4902 8226
rect 4868 8139 4902 8141
rect 4868 8103 4902 8105
rect 4868 8018 4902 8037
rect 5700 8208 5734 8226
rect 5700 8140 5734 8142
rect 5700 8104 5734 8106
rect 5700 8018 5734 8038
rect 5858 8208 5892 8226
rect 5858 8140 5892 8142
rect 5858 8104 5892 8106
rect 5858 8018 5892 8038
rect 6008 8208 6042 8226
rect 6008 8140 6042 8142
rect 6008 8104 6042 8106
rect 6008 8018 6042 8038
rect 6166 8208 6200 8226
rect 6166 8140 6200 8142
rect 6166 8104 6200 8106
rect 6166 8018 6200 8038
rect 6360 8208 6394 8226
rect 6360 8140 6394 8142
rect 6360 8104 6394 8106
rect 6360 8018 6394 8038
rect 6518 8208 6552 8226
rect 6518 8140 6552 8142
rect 6518 8104 6552 8106
rect 6518 8018 6552 8038
rect 6668 8208 6702 8226
rect 6668 8140 6702 8142
rect 6668 8104 6702 8106
rect 6668 8018 6702 8038
rect 6826 8208 6860 8226
rect 6826 8140 6860 8142
rect 6826 8104 6860 8106
rect 6826 8018 6860 8038
rect 3670 7982 3704 7995
rect 3668 7979 3707 7982
rect 1773 7909 1807 7918
rect 2261 7911 2319 7923
rect 2625 7912 2703 7926
rect 2850 7921 2857 7955
rect 2891 7921 2898 7955
rect 3013 7921 3029 7955
rect 3063 7921 3079 7955
rect 3668 7945 3670 7979
rect 3704 7945 3707 7979
rect 3984 7973 4018 7986
rect 5628 7982 5662 7996
rect 3668 7943 3707 7945
rect 3982 7970 4021 7973
rect 3670 7929 3704 7943
rect 3982 7936 3984 7970
rect 4018 7936 4021 7970
rect 3982 7934 4021 7936
rect 4306 7965 4340 7980
rect 4306 7964 4341 7965
rect 2850 7914 2898 7921
rect 1255 7895 1318 7907
rect 2271 7905 2309 7911
rect 1410 7841 1444 7878
rect 556 7752 616 7768
rect 556 7728 565 7752
rect 606 7728 616 7752
rect 702 7752 762 7768
rect 702 7728 712 7752
rect 753 7728 762 7752
rect 846 7757 906 7774
rect 846 7734 856 7757
rect 897 7734 906 7757
rect 1000 7758 1060 7774
rect 1410 7770 1444 7807
rect 1568 7841 1602 7878
rect 1568 7770 1602 7807
rect 1698 7841 1732 7878
rect 1698 7770 1732 7807
rect 1856 7841 1890 7878
rect 1856 7770 1890 7807
rect 2030 7841 2064 7878
rect 2030 7770 2064 7807
rect 2188 7841 2222 7878
rect 2188 7770 2222 7807
rect 2352 7841 2420 7884
rect 2352 7807 2372 7841
rect 2406 7807 2420 7841
rect 1000 7734 1010 7758
rect 1051 7734 1060 7758
rect 540 7712 565 7728
rect 606 7712 632 7728
rect 540 7694 569 7712
rect 603 7694 632 7712
rect 686 7712 712 7728
rect 753 7712 778 7728
rect 686 7694 715 7712
rect 749 7694 778 7712
rect 830 7717 856 7734
rect 897 7717 922 7734
rect 830 7700 859 7717
rect 893 7700 922 7717
rect 984 7718 1010 7734
rect 1051 7718 1076 7734
rect 984 7700 1013 7718
rect 1047 7700 1076 7718
rect 1324 7664 1960 7728
rect 1324 7630 1353 7664
rect 1407 7630 1421 7664
rect 1479 7630 1489 7664
rect 1551 7630 1557 7664
rect 1623 7630 1625 7664
rect 1659 7630 1661 7664
rect 1727 7630 1733 7664
rect 1795 7630 1805 7664
rect 1863 7630 1877 7664
rect 1931 7630 1960 7664
rect 1324 7588 1960 7630
rect 2352 7639 2420 7807
rect 2530 7841 2564 7878
rect 2530 7770 2564 7807
rect 2352 7605 2369 7639
rect 2403 7605 2420 7639
rect 2352 7588 2420 7605
rect 2642 7543 2696 7912
rect 2857 7905 2891 7914
rect 3019 7911 3073 7921
rect 3984 7920 4018 7934
rect 4340 7930 4341 7964
rect 4621 7948 4637 7982
rect 4671 7948 4687 7982
rect 5626 7980 5666 7982
rect 5626 7946 5628 7980
rect 5662 7946 5666 7980
rect 5942 7974 5976 7986
rect 5626 7944 5666 7946
rect 5940 7970 5980 7974
rect 5628 7930 5662 7944
rect 5940 7936 5942 7970
rect 5976 7936 5980 7970
rect 5940 7934 5980 7936
rect 6264 7966 6298 7980
rect 6264 7964 6300 7966
rect 4306 7914 4340 7930
rect 5942 7920 5976 7934
rect 6298 7930 6300 7964
rect 6580 7948 6596 7982
rect 6630 7948 6646 7982
rect 6264 7914 6298 7930
rect 2776 7841 2810 7878
rect 2776 7770 2810 7807
rect 2934 7841 2968 7878
rect 2934 7770 2968 7807
rect 3120 7841 3154 7878
rect 3120 7770 3154 7807
rect 3278 7841 3312 7878
rect 3278 7770 3312 7807
rect 3742 7851 3776 7888
rect 3742 7780 3776 7817
rect 3900 7851 3934 7888
rect 3900 7780 3934 7817
rect 4050 7851 4084 7888
rect 4050 7780 4084 7817
rect 4208 7851 4242 7888
rect 4208 7780 4242 7817
rect 4402 7853 4436 7890
rect 4402 7782 4436 7819
rect 4560 7853 4594 7890
rect 4560 7782 4594 7819
rect 4710 7853 4744 7890
rect 4710 7782 4744 7819
rect 4868 7853 4902 7890
rect 4868 7782 4902 7819
rect 5700 7852 5734 7888
rect 5700 7780 5734 7818
rect 5858 7852 5892 7888
rect 5858 7780 5892 7818
rect 6008 7852 6042 7888
rect 6008 7780 6042 7818
rect 6166 7852 6200 7888
rect 6166 7780 6200 7818
rect 6360 7854 6394 7890
rect 6360 7782 6394 7820
rect 6518 7854 6552 7890
rect 6518 7782 6552 7820
rect 6668 7854 6702 7890
rect 6668 7782 6702 7820
rect 6826 7854 6860 7890
rect 6826 7782 6860 7820
rect 3704 7675 4244 7728
rect 3704 7641 3741 7675
rect 3787 7641 3813 7675
rect 3855 7641 3885 7675
rect 3923 7641 3957 7675
rect 3991 7641 4025 7675
rect 4063 7641 4093 7675
rect 4135 7641 4161 7675
rect 4207 7641 4244 7675
rect 3704 7588 4244 7641
rect 5662 7676 6202 7728
rect 5662 7642 5700 7676
rect 5746 7642 5772 7676
rect 5814 7642 5844 7676
rect 5882 7642 5916 7676
rect 5950 7642 5984 7676
rect 6022 7642 6052 7676
rect 6094 7642 6120 7676
rect 6166 7642 6202 7676
rect 5662 7588 6202 7642
rect 1348 7138 1880 7190
rect 1348 7104 1383 7138
rect 1429 7104 1455 7138
rect 1497 7104 1527 7138
rect 1565 7104 1599 7138
rect 1633 7104 1667 7138
rect 1705 7104 1735 7138
rect 1777 7104 1803 7138
rect 1849 7104 1880 7138
rect 3724 7137 4264 7190
rect 540 7052 569 7068
rect 603 7052 632 7068
rect 540 7034 566 7052
rect 607 7034 632 7052
rect 686 7052 715 7068
rect 749 7052 778 7068
rect 686 7034 710 7052
rect 751 7034 778 7052
rect 830 7057 859 7074
rect 893 7057 922 7074
rect 830 7040 856 7057
rect 897 7040 922 7057
rect 984 7057 1013 7074
rect 1047 7057 1076 7074
rect 984 7040 1009 7057
rect 1050 7040 1076 7057
rect 1348 7050 1880 7104
rect 2627 7057 3073 7111
rect 556 7012 566 7034
rect 607 7012 616 7034
rect 556 6994 616 7012
rect 702 7012 710 7034
rect 751 7012 762 7034
rect 702 6994 762 7012
rect 846 7017 856 7040
rect 897 7017 906 7040
rect 846 7000 906 7017
rect 1000 7017 1009 7040
rect 1050 7017 1060 7040
rect 1000 7000 1060 7017
rect 1410 6969 1444 6988
rect 1410 6901 1444 6903
rect 1410 6865 1444 6867
rect 1410 6780 1444 6799
rect 1568 6969 1602 6988
rect 1568 6901 1602 6903
rect 1568 6865 1602 6867
rect 1568 6780 1602 6799
rect 1698 6969 1732 6988
rect 1698 6901 1732 6903
rect 1698 6865 1732 6867
rect 1698 6780 1732 6799
rect 1856 6969 1890 6988
rect 1856 6901 1890 6903
rect 1856 6865 1890 6867
rect 1856 6780 1890 6799
rect 2030 6969 2064 6988
rect 2030 6901 2064 6903
rect 2030 6865 2064 6867
rect 2030 6780 2064 6799
rect 2188 6969 2222 6988
rect 2188 6901 2222 6903
rect 2188 6865 2222 6867
rect 2188 6780 2222 6799
rect 2372 6969 2406 6988
rect 2372 6901 2406 6903
rect 2372 6865 2406 6867
rect 2372 6780 2406 6799
rect 2530 6969 2564 6988
rect 2627 6907 2681 7057
rect 2776 6969 2810 6988
rect 2530 6901 2564 6903
rect 2530 6865 2564 6867
rect 2530 6780 2564 6799
rect 2625 6885 2703 6907
rect 2625 6851 2647 6885
rect 2681 6851 2703 6885
rect 1255 6750 1318 6762
rect 1251 6731 1322 6750
rect 2625 6747 2703 6851
rect 2776 6901 2810 6903
rect 2776 6865 2810 6867
rect 2776 6780 2810 6799
rect 2934 6969 2968 6988
rect 2934 6901 2968 6903
rect 2934 6865 2968 6867
rect 2934 6780 2968 6799
rect 1773 6738 1807 6747
rect 2271 6741 2309 6747
rect 1251 6697 1269 6731
rect 1303 6697 1322 6731
rect 1251 6679 1322 6697
rect 1766 6731 1814 6738
rect 1766 6697 1773 6731
rect 1807 6697 1814 6731
rect 1766 6690 1814 6697
rect 2261 6729 2319 6741
rect 2261 6695 2273 6729
rect 2307 6695 2319 6729
rect 2615 6739 2713 6747
rect 2615 6705 2647 6739
rect 2681 6705 2713 6739
rect 2857 6734 2891 6743
rect 2615 6698 2713 6705
rect 2850 6727 2898 6734
rect 3019 6727 3073 7057
rect 3724 7103 3773 7137
rect 3831 7103 3841 7137
rect 3903 7103 3909 7137
rect 3975 7103 3977 7137
rect 4011 7103 4013 7137
rect 4079 7103 4085 7137
rect 4147 7103 4157 7137
rect 4215 7103 4264 7137
rect 3724 7050 4264 7103
rect 5682 7136 6222 7190
rect 5682 7102 5732 7136
rect 5790 7102 5800 7136
rect 5862 7102 5868 7136
rect 5934 7102 5936 7136
rect 5970 7102 5972 7136
rect 6038 7102 6044 7136
rect 6106 7102 6116 7136
rect 6174 7102 6222 7136
rect 5682 7050 6222 7102
rect 3120 6969 3154 6988
rect 3120 6901 3154 6903
rect 3120 6865 3154 6867
rect 3120 6780 3154 6799
rect 3278 6969 3312 6988
rect 3278 6901 3312 6903
rect 3278 6865 3312 6867
rect 3278 6780 3312 6799
rect 3742 6979 3776 6998
rect 3742 6911 3776 6913
rect 3742 6875 3776 6877
rect 3742 6790 3776 6809
rect 3900 6979 3934 6998
rect 3900 6911 3934 6913
rect 3900 6875 3934 6877
rect 3900 6790 3934 6809
rect 4050 6979 4084 6998
rect 4050 6911 4084 6913
rect 4050 6875 4084 6877
rect 4050 6790 4084 6809
rect 4208 6979 4242 6998
rect 4208 6911 4242 6913
rect 4208 6875 4242 6877
rect 4208 6790 4242 6809
rect 4402 6979 4436 6998
rect 4402 6911 4436 6913
rect 4402 6875 4436 6877
rect 4402 6790 4436 6809
rect 4560 6979 4594 6998
rect 4560 6911 4594 6913
rect 4560 6875 4594 6877
rect 4560 6790 4594 6809
rect 4710 6979 4744 6998
rect 4710 6911 4744 6913
rect 4710 6875 4744 6877
rect 4710 6790 4744 6809
rect 4868 6979 4902 6998
rect 4868 6911 4902 6913
rect 4868 6875 4902 6877
rect 4868 6790 4902 6809
rect 5700 6980 5734 6998
rect 5700 6912 5734 6914
rect 5700 6876 5734 6878
rect 5700 6790 5734 6810
rect 5858 6980 5892 6998
rect 5858 6912 5892 6914
rect 5858 6876 5892 6878
rect 5858 6790 5892 6810
rect 6008 6980 6042 6998
rect 6008 6912 6042 6914
rect 6008 6876 6042 6878
rect 6008 6790 6042 6810
rect 6166 6980 6200 6998
rect 6166 6912 6200 6914
rect 6166 6876 6200 6878
rect 6166 6790 6200 6810
rect 6360 6980 6394 6998
rect 6360 6912 6394 6914
rect 6360 6876 6394 6878
rect 6360 6790 6394 6810
rect 6518 6980 6552 6998
rect 6518 6912 6552 6914
rect 6518 6876 6552 6878
rect 6518 6790 6552 6810
rect 6668 6980 6702 6998
rect 6668 6912 6702 6914
rect 6668 6876 6702 6878
rect 6668 6790 6702 6810
rect 6826 6980 6860 6998
rect 6826 6912 6860 6914
rect 6826 6876 6860 6878
rect 6826 6790 6860 6810
rect 3670 6754 3704 6767
rect 3668 6751 3707 6754
rect 1773 6681 1807 6690
rect 2261 6683 2319 6695
rect 2625 6684 2703 6698
rect 2850 6693 2857 6727
rect 2891 6693 2898 6727
rect 3013 6693 3029 6727
rect 3063 6693 3079 6727
rect 3668 6717 3670 6751
rect 3704 6717 3707 6751
rect 3984 6745 4018 6758
rect 5628 6754 5662 6768
rect 3668 6715 3707 6717
rect 3982 6742 4021 6745
rect 3670 6701 3704 6715
rect 3982 6708 3984 6742
rect 4018 6708 4021 6742
rect 3982 6706 4021 6708
rect 4306 6737 4340 6752
rect 4306 6736 4341 6737
rect 2850 6686 2898 6693
rect 1255 6667 1318 6679
rect 2271 6677 2309 6683
rect 1410 6613 1444 6650
rect 556 6524 616 6540
rect 556 6500 565 6524
rect 606 6500 616 6524
rect 702 6524 762 6540
rect 702 6500 712 6524
rect 753 6500 762 6524
rect 846 6529 906 6546
rect 846 6506 856 6529
rect 897 6506 906 6529
rect 1000 6530 1060 6546
rect 1410 6542 1444 6579
rect 1568 6613 1602 6650
rect 1568 6542 1602 6579
rect 1698 6613 1732 6650
rect 1698 6542 1732 6579
rect 1856 6613 1890 6650
rect 1856 6542 1890 6579
rect 2030 6613 2064 6650
rect 2030 6542 2064 6579
rect 2188 6613 2222 6650
rect 2188 6542 2222 6579
rect 2352 6613 2420 6656
rect 2352 6579 2372 6613
rect 2406 6579 2420 6613
rect 1000 6506 1010 6530
rect 1051 6506 1060 6530
rect 540 6484 565 6500
rect 606 6484 632 6500
rect 540 6466 569 6484
rect 603 6466 632 6484
rect 686 6484 712 6500
rect 753 6484 778 6500
rect 686 6466 715 6484
rect 749 6466 778 6484
rect 830 6489 856 6506
rect 897 6489 922 6506
rect 830 6472 859 6489
rect 893 6472 922 6489
rect 984 6490 1010 6506
rect 1051 6490 1076 6506
rect 984 6472 1013 6490
rect 1047 6472 1076 6490
rect 1324 6436 1960 6500
rect 1324 6402 1353 6436
rect 1407 6402 1421 6436
rect 1479 6402 1489 6436
rect 1551 6402 1557 6436
rect 1623 6402 1625 6436
rect 1659 6402 1661 6436
rect 1727 6402 1733 6436
rect 1795 6402 1805 6436
rect 1863 6402 1877 6436
rect 1931 6402 1960 6436
rect 1324 6360 1960 6402
rect 2352 6411 2420 6579
rect 2530 6613 2564 6650
rect 2530 6542 2564 6579
rect 2352 6377 2369 6411
rect 2403 6377 2420 6411
rect 2352 6360 2420 6377
rect 2642 6315 2696 6684
rect 2857 6677 2891 6686
rect 3019 6683 3073 6693
rect 3984 6692 4018 6706
rect 4340 6702 4341 6736
rect 4621 6720 4637 6754
rect 4671 6720 4687 6754
rect 5626 6752 5666 6754
rect 5626 6718 5628 6752
rect 5662 6718 5666 6752
rect 5942 6746 5976 6758
rect 5626 6716 5666 6718
rect 5940 6742 5980 6746
rect 5628 6702 5662 6716
rect 5940 6708 5942 6742
rect 5976 6708 5980 6742
rect 5940 6706 5980 6708
rect 6264 6738 6298 6752
rect 6264 6736 6300 6738
rect 4306 6686 4340 6702
rect 5942 6692 5976 6706
rect 6298 6702 6300 6736
rect 6580 6720 6596 6754
rect 6630 6720 6646 6754
rect 6264 6686 6298 6702
rect 2776 6613 2810 6650
rect 2776 6542 2810 6579
rect 2934 6613 2968 6650
rect 2934 6542 2968 6579
rect 3120 6613 3154 6650
rect 3120 6542 3154 6579
rect 3278 6613 3312 6650
rect 3278 6542 3312 6579
rect 3742 6623 3776 6660
rect 3742 6552 3776 6589
rect 3900 6623 3934 6660
rect 3900 6552 3934 6589
rect 4050 6623 4084 6660
rect 4050 6552 4084 6589
rect 4208 6623 4242 6660
rect 4208 6552 4242 6589
rect 4402 6625 4436 6662
rect 4402 6554 4436 6591
rect 4560 6625 4594 6662
rect 4560 6554 4594 6591
rect 4710 6625 4744 6662
rect 4710 6554 4744 6591
rect 4868 6625 4902 6662
rect 4868 6554 4902 6591
rect 5700 6624 5734 6660
rect 5700 6552 5734 6590
rect 5858 6624 5892 6660
rect 5858 6552 5892 6590
rect 6008 6624 6042 6660
rect 6008 6552 6042 6590
rect 6166 6624 6200 6660
rect 6166 6552 6200 6590
rect 6360 6626 6394 6662
rect 6360 6554 6394 6592
rect 6518 6626 6552 6662
rect 6518 6554 6552 6592
rect 6668 6626 6702 6662
rect 6668 6554 6702 6592
rect 6826 6626 6860 6662
rect 6826 6554 6860 6592
rect 3704 6447 4244 6500
rect 3704 6413 3741 6447
rect 3787 6413 3813 6447
rect 3855 6413 3885 6447
rect 3923 6413 3957 6447
rect 3991 6413 4025 6447
rect 4063 6413 4093 6447
rect 4135 6413 4161 6447
rect 4207 6413 4244 6447
rect 3704 6360 4244 6413
rect 5662 6448 6202 6500
rect 5662 6414 5700 6448
rect 5746 6414 5772 6448
rect 5814 6414 5844 6448
rect 5882 6414 5916 6448
rect 5950 6414 5984 6448
rect 6022 6414 6052 6448
rect 6094 6414 6120 6448
rect 6166 6414 6202 6448
rect 5662 6360 6202 6414
rect 1348 5910 1880 5962
rect 1348 5876 1383 5910
rect 1429 5876 1455 5910
rect 1497 5876 1527 5910
rect 1565 5876 1599 5910
rect 1633 5876 1667 5910
rect 1705 5876 1735 5910
rect 1777 5876 1803 5910
rect 1849 5876 1880 5910
rect 3724 5909 4264 5962
rect 540 5824 569 5840
rect 603 5824 632 5840
rect 540 5806 566 5824
rect 607 5806 632 5824
rect 686 5824 715 5840
rect 749 5824 778 5840
rect 686 5806 710 5824
rect 751 5806 778 5824
rect 830 5829 859 5846
rect 893 5829 922 5846
rect 830 5812 856 5829
rect 897 5812 922 5829
rect 984 5829 1013 5846
rect 1047 5829 1076 5846
rect 984 5812 1009 5829
rect 1050 5812 1076 5829
rect 1348 5822 1880 5876
rect 2627 5829 3073 5883
rect 556 5784 566 5806
rect 607 5784 616 5806
rect 556 5766 616 5784
rect 702 5784 710 5806
rect 751 5784 762 5806
rect 702 5766 762 5784
rect 846 5789 856 5812
rect 897 5789 906 5812
rect 846 5772 906 5789
rect 1000 5789 1009 5812
rect 1050 5789 1060 5812
rect 1000 5772 1060 5789
rect 1410 5741 1444 5760
rect 1410 5673 1444 5675
rect 1410 5637 1444 5639
rect 1410 5552 1444 5571
rect 1568 5741 1602 5760
rect 1568 5673 1602 5675
rect 1568 5637 1602 5639
rect 1568 5552 1602 5571
rect 1698 5741 1732 5760
rect 1698 5673 1732 5675
rect 1698 5637 1732 5639
rect 1698 5552 1732 5571
rect 1856 5741 1890 5760
rect 1856 5673 1890 5675
rect 1856 5637 1890 5639
rect 1856 5552 1890 5571
rect 2030 5741 2064 5760
rect 2030 5673 2064 5675
rect 2030 5637 2064 5639
rect 2030 5552 2064 5571
rect 2188 5741 2222 5760
rect 2188 5673 2222 5675
rect 2188 5637 2222 5639
rect 2188 5552 2222 5571
rect 2372 5741 2406 5760
rect 2372 5673 2406 5675
rect 2372 5637 2406 5639
rect 2372 5552 2406 5571
rect 2530 5741 2564 5760
rect 2627 5679 2681 5829
rect 2776 5741 2810 5760
rect 2530 5673 2564 5675
rect 2530 5637 2564 5639
rect 2530 5552 2564 5571
rect 2625 5657 2703 5679
rect 2625 5623 2647 5657
rect 2681 5623 2703 5657
rect 1255 5522 1318 5534
rect 1251 5503 1322 5522
rect 2625 5519 2703 5623
rect 2776 5673 2810 5675
rect 2776 5637 2810 5639
rect 2776 5552 2810 5571
rect 2934 5741 2968 5760
rect 2934 5673 2968 5675
rect 2934 5637 2968 5639
rect 2934 5552 2968 5571
rect 1773 5510 1807 5519
rect 2271 5513 2309 5519
rect 1251 5469 1269 5503
rect 1303 5469 1322 5503
rect 1251 5451 1322 5469
rect 1766 5503 1814 5510
rect 1766 5469 1773 5503
rect 1807 5469 1814 5503
rect 1766 5462 1814 5469
rect 2261 5501 2319 5513
rect 2261 5467 2273 5501
rect 2307 5467 2319 5501
rect 2615 5511 2713 5519
rect 2615 5477 2647 5511
rect 2681 5477 2713 5511
rect 2857 5506 2891 5515
rect 2615 5470 2713 5477
rect 2850 5499 2898 5506
rect 3019 5499 3073 5829
rect 3724 5875 3773 5909
rect 3831 5875 3841 5909
rect 3903 5875 3909 5909
rect 3975 5875 3977 5909
rect 4011 5875 4013 5909
rect 4079 5875 4085 5909
rect 4147 5875 4157 5909
rect 4215 5875 4264 5909
rect 3724 5822 4264 5875
rect 5682 5908 6222 5962
rect 5682 5874 5732 5908
rect 5790 5874 5800 5908
rect 5862 5874 5868 5908
rect 5934 5874 5936 5908
rect 5970 5874 5972 5908
rect 6038 5874 6044 5908
rect 6106 5874 6116 5908
rect 6174 5874 6222 5908
rect 5682 5822 6222 5874
rect 3120 5741 3154 5760
rect 3120 5673 3154 5675
rect 3120 5637 3154 5639
rect 3120 5552 3154 5571
rect 3278 5741 3312 5760
rect 3278 5673 3312 5675
rect 3278 5637 3312 5639
rect 3278 5552 3312 5571
rect 3742 5751 3776 5770
rect 3742 5683 3776 5685
rect 3742 5647 3776 5649
rect 3742 5562 3776 5581
rect 3900 5751 3934 5770
rect 3900 5683 3934 5685
rect 3900 5647 3934 5649
rect 3900 5562 3934 5581
rect 4050 5751 4084 5770
rect 4050 5683 4084 5685
rect 4050 5647 4084 5649
rect 4050 5562 4084 5581
rect 4208 5751 4242 5770
rect 4208 5683 4242 5685
rect 4208 5647 4242 5649
rect 4208 5562 4242 5581
rect 4402 5751 4436 5770
rect 4402 5683 4436 5685
rect 4402 5647 4436 5649
rect 4402 5562 4436 5581
rect 4560 5751 4594 5770
rect 4560 5683 4594 5685
rect 4560 5647 4594 5649
rect 4560 5562 4594 5581
rect 4710 5751 4744 5770
rect 4710 5683 4744 5685
rect 4710 5647 4744 5649
rect 4710 5562 4744 5581
rect 4868 5751 4902 5770
rect 4868 5683 4902 5685
rect 4868 5647 4902 5649
rect 4868 5562 4902 5581
rect 5700 5752 5734 5770
rect 5700 5684 5734 5686
rect 5700 5648 5734 5650
rect 5700 5562 5734 5582
rect 5858 5752 5892 5770
rect 5858 5684 5892 5686
rect 5858 5648 5892 5650
rect 5858 5562 5892 5582
rect 6008 5752 6042 5770
rect 6008 5684 6042 5686
rect 6008 5648 6042 5650
rect 6008 5562 6042 5582
rect 6166 5752 6200 5770
rect 6166 5684 6200 5686
rect 6166 5648 6200 5650
rect 6166 5562 6200 5582
rect 6360 5752 6394 5770
rect 6360 5684 6394 5686
rect 6360 5648 6394 5650
rect 6360 5562 6394 5582
rect 6518 5752 6552 5770
rect 6518 5684 6552 5686
rect 6518 5648 6552 5650
rect 6518 5562 6552 5582
rect 6668 5752 6702 5770
rect 6668 5684 6702 5686
rect 6668 5648 6702 5650
rect 6668 5562 6702 5582
rect 6826 5752 6860 5770
rect 6826 5684 6860 5686
rect 6826 5648 6860 5650
rect 6826 5562 6860 5582
rect 3670 5526 3704 5539
rect 3668 5523 3707 5526
rect 1773 5453 1807 5462
rect 2261 5455 2319 5467
rect 2625 5456 2703 5470
rect 2850 5465 2857 5499
rect 2891 5465 2898 5499
rect 3013 5465 3029 5499
rect 3063 5465 3079 5499
rect 3668 5489 3670 5523
rect 3704 5489 3707 5523
rect 3984 5517 4018 5530
rect 5628 5526 5662 5540
rect 3668 5487 3707 5489
rect 3982 5514 4021 5517
rect 3670 5473 3704 5487
rect 3982 5480 3984 5514
rect 4018 5480 4021 5514
rect 3982 5478 4021 5480
rect 4306 5509 4340 5524
rect 4306 5508 4341 5509
rect 2850 5458 2898 5465
rect 1255 5439 1318 5451
rect 2271 5449 2309 5455
rect 1410 5385 1444 5422
rect 556 5296 616 5312
rect 556 5272 565 5296
rect 606 5272 616 5296
rect 702 5296 762 5312
rect 702 5272 712 5296
rect 753 5272 762 5296
rect 846 5301 906 5318
rect 846 5278 856 5301
rect 897 5278 906 5301
rect 1000 5302 1060 5318
rect 1410 5314 1444 5351
rect 1568 5385 1602 5422
rect 1568 5314 1602 5351
rect 1698 5385 1732 5422
rect 1698 5314 1732 5351
rect 1856 5385 1890 5422
rect 1856 5314 1890 5351
rect 2030 5385 2064 5422
rect 2030 5314 2064 5351
rect 2188 5385 2222 5422
rect 2188 5314 2222 5351
rect 2352 5385 2420 5428
rect 2352 5351 2372 5385
rect 2406 5351 2420 5385
rect 1000 5278 1010 5302
rect 1051 5278 1060 5302
rect 540 5256 565 5272
rect 606 5256 632 5272
rect 540 5238 569 5256
rect 603 5238 632 5256
rect 686 5256 712 5272
rect 753 5256 778 5272
rect 686 5238 715 5256
rect 749 5238 778 5256
rect 830 5261 856 5278
rect 897 5261 922 5278
rect 830 5244 859 5261
rect 893 5244 922 5261
rect 984 5262 1010 5278
rect 1051 5262 1076 5278
rect 984 5244 1013 5262
rect 1047 5244 1076 5262
rect 1324 5208 1960 5272
rect 1324 5174 1353 5208
rect 1407 5174 1421 5208
rect 1479 5174 1489 5208
rect 1551 5174 1557 5208
rect 1623 5174 1625 5208
rect 1659 5174 1661 5208
rect 1727 5174 1733 5208
rect 1795 5174 1805 5208
rect 1863 5174 1877 5208
rect 1931 5174 1960 5208
rect 1324 5132 1960 5174
rect 2352 5183 2420 5351
rect 2530 5385 2564 5422
rect 2530 5314 2564 5351
rect 2352 5149 2369 5183
rect 2403 5149 2420 5183
rect 2352 5132 2420 5149
rect 2642 5087 2696 5456
rect 2857 5449 2891 5458
rect 3019 5455 3073 5465
rect 3984 5464 4018 5478
rect 4340 5474 4341 5508
rect 4621 5492 4637 5526
rect 4671 5492 4687 5526
rect 5626 5524 5666 5526
rect 5626 5490 5628 5524
rect 5662 5490 5666 5524
rect 5942 5518 5976 5530
rect 5626 5488 5666 5490
rect 5940 5514 5980 5518
rect 5628 5474 5662 5488
rect 5940 5480 5942 5514
rect 5976 5480 5980 5514
rect 5940 5478 5980 5480
rect 6264 5510 6298 5524
rect 6264 5508 6300 5510
rect 4306 5458 4340 5474
rect 5942 5464 5976 5478
rect 6298 5474 6300 5508
rect 6580 5492 6596 5526
rect 6630 5492 6646 5526
rect 6264 5458 6298 5474
rect 2776 5385 2810 5422
rect 2776 5314 2810 5351
rect 2934 5385 2968 5422
rect 2934 5314 2968 5351
rect 3120 5385 3154 5422
rect 3120 5314 3154 5351
rect 3278 5385 3312 5422
rect 3278 5314 3312 5351
rect 3742 5395 3776 5432
rect 3742 5324 3776 5361
rect 3900 5395 3934 5432
rect 3900 5324 3934 5361
rect 4050 5395 4084 5432
rect 4050 5324 4084 5361
rect 4208 5395 4242 5432
rect 4208 5324 4242 5361
rect 4402 5397 4436 5434
rect 4402 5326 4436 5363
rect 4560 5397 4594 5434
rect 4560 5326 4594 5363
rect 4710 5397 4744 5434
rect 4710 5326 4744 5363
rect 4868 5397 4902 5434
rect 4868 5326 4902 5363
rect 5700 5396 5734 5432
rect 5700 5324 5734 5362
rect 5858 5396 5892 5432
rect 5858 5324 5892 5362
rect 6008 5396 6042 5432
rect 6008 5324 6042 5362
rect 6166 5396 6200 5432
rect 6166 5324 6200 5362
rect 6360 5398 6394 5434
rect 6360 5326 6394 5364
rect 6518 5398 6552 5434
rect 6518 5326 6552 5364
rect 6668 5398 6702 5434
rect 6668 5326 6702 5364
rect 6826 5398 6860 5434
rect 6826 5326 6860 5364
rect 3704 5219 4244 5272
rect 3704 5185 3741 5219
rect 3787 5185 3813 5219
rect 3855 5185 3885 5219
rect 3923 5185 3957 5219
rect 3991 5185 4025 5219
rect 4063 5185 4093 5219
rect 4135 5185 4161 5219
rect 4207 5185 4244 5219
rect 3704 5132 4244 5185
rect 5662 5220 6202 5272
rect 5662 5186 5700 5220
rect 5746 5186 5772 5220
rect 5814 5186 5844 5220
rect 5882 5186 5916 5220
rect 5950 5186 5984 5220
rect 6022 5186 6052 5220
rect 6094 5186 6120 5220
rect 6166 5186 6202 5220
rect 5662 5132 6202 5186
rect 1348 4682 1880 4734
rect 1348 4648 1383 4682
rect 1429 4648 1455 4682
rect 1497 4648 1527 4682
rect 1565 4648 1599 4682
rect 1633 4648 1667 4682
rect 1705 4648 1735 4682
rect 1777 4648 1803 4682
rect 1849 4648 1880 4682
rect 3724 4681 4264 4734
rect 540 4596 569 4612
rect 603 4596 632 4612
rect 540 4578 566 4596
rect 607 4578 632 4596
rect 686 4596 715 4612
rect 749 4596 778 4612
rect 686 4578 710 4596
rect 751 4578 778 4596
rect 830 4601 859 4618
rect 893 4601 922 4618
rect 830 4584 856 4601
rect 897 4584 922 4601
rect 984 4601 1013 4618
rect 1047 4601 1076 4618
rect 984 4584 1009 4601
rect 1050 4584 1076 4601
rect 1348 4594 1880 4648
rect 2627 4601 3073 4655
rect 556 4556 566 4578
rect 607 4556 616 4578
rect 556 4538 616 4556
rect 702 4556 710 4578
rect 751 4556 762 4578
rect 702 4538 762 4556
rect 846 4561 856 4584
rect 897 4561 906 4584
rect 846 4544 906 4561
rect 1000 4561 1009 4584
rect 1050 4561 1060 4584
rect 1000 4544 1060 4561
rect 1410 4513 1444 4532
rect 1410 4445 1444 4447
rect 1410 4409 1444 4411
rect 1410 4324 1444 4343
rect 1568 4513 1602 4532
rect 1568 4445 1602 4447
rect 1568 4409 1602 4411
rect 1568 4324 1602 4343
rect 1698 4513 1732 4532
rect 1698 4445 1732 4447
rect 1698 4409 1732 4411
rect 1698 4324 1732 4343
rect 1856 4513 1890 4532
rect 1856 4445 1890 4447
rect 1856 4409 1890 4411
rect 1856 4324 1890 4343
rect 2030 4513 2064 4532
rect 2030 4445 2064 4447
rect 2030 4409 2064 4411
rect 2030 4324 2064 4343
rect 2188 4513 2222 4532
rect 2188 4445 2222 4447
rect 2188 4409 2222 4411
rect 2188 4324 2222 4343
rect 2372 4513 2406 4532
rect 2372 4445 2406 4447
rect 2372 4409 2406 4411
rect 2372 4324 2406 4343
rect 2530 4513 2564 4532
rect 2627 4451 2681 4601
rect 2776 4513 2810 4532
rect 2530 4445 2564 4447
rect 2530 4409 2564 4411
rect 2530 4324 2564 4343
rect 2625 4429 2703 4451
rect 2625 4395 2647 4429
rect 2681 4395 2703 4429
rect 1255 4294 1318 4306
rect 1251 4275 1322 4294
rect 2625 4291 2703 4395
rect 2776 4445 2810 4447
rect 2776 4409 2810 4411
rect 2776 4324 2810 4343
rect 2934 4513 2968 4532
rect 2934 4445 2968 4447
rect 2934 4409 2968 4411
rect 2934 4324 2968 4343
rect 1773 4282 1807 4291
rect 2271 4285 2309 4291
rect 1251 4241 1269 4275
rect 1303 4241 1322 4275
rect 1251 4223 1322 4241
rect 1766 4275 1814 4282
rect 1766 4241 1773 4275
rect 1807 4241 1814 4275
rect 1766 4234 1814 4241
rect 2261 4273 2319 4285
rect 2261 4239 2273 4273
rect 2307 4239 2319 4273
rect 2615 4283 2713 4291
rect 2615 4249 2647 4283
rect 2681 4249 2713 4283
rect 2857 4278 2891 4287
rect 2615 4242 2713 4249
rect 2850 4271 2898 4278
rect 3019 4271 3073 4601
rect 3724 4647 3773 4681
rect 3831 4647 3841 4681
rect 3903 4647 3909 4681
rect 3975 4647 3977 4681
rect 4011 4647 4013 4681
rect 4079 4647 4085 4681
rect 4147 4647 4157 4681
rect 4215 4647 4264 4681
rect 3724 4594 4264 4647
rect 5682 4680 6222 4734
rect 5682 4646 5732 4680
rect 5790 4646 5800 4680
rect 5862 4646 5868 4680
rect 5934 4646 5936 4680
rect 5970 4646 5972 4680
rect 6038 4646 6044 4680
rect 6106 4646 6116 4680
rect 6174 4646 6222 4680
rect 5682 4594 6222 4646
rect 3120 4513 3154 4532
rect 3120 4445 3154 4447
rect 3120 4409 3154 4411
rect 3120 4324 3154 4343
rect 3278 4513 3312 4532
rect 3278 4445 3312 4447
rect 3278 4409 3312 4411
rect 3278 4324 3312 4343
rect 3742 4523 3776 4542
rect 3742 4455 3776 4457
rect 3742 4419 3776 4421
rect 3742 4334 3776 4353
rect 3900 4523 3934 4542
rect 3900 4455 3934 4457
rect 3900 4419 3934 4421
rect 3900 4334 3934 4353
rect 4050 4523 4084 4542
rect 4050 4455 4084 4457
rect 4050 4419 4084 4421
rect 4050 4334 4084 4353
rect 4208 4523 4242 4542
rect 4208 4455 4242 4457
rect 4208 4419 4242 4421
rect 4208 4334 4242 4353
rect 4402 4523 4436 4542
rect 4402 4455 4436 4457
rect 4402 4419 4436 4421
rect 4402 4334 4436 4353
rect 4560 4523 4594 4542
rect 4560 4455 4594 4457
rect 4560 4419 4594 4421
rect 4560 4334 4594 4353
rect 4710 4523 4744 4542
rect 4710 4455 4744 4457
rect 4710 4419 4744 4421
rect 4710 4334 4744 4353
rect 4868 4523 4902 4542
rect 4868 4455 4902 4457
rect 4868 4419 4902 4421
rect 4868 4334 4902 4353
rect 5700 4524 5734 4542
rect 5700 4456 5734 4458
rect 5700 4420 5734 4422
rect 5700 4334 5734 4354
rect 5858 4524 5892 4542
rect 5858 4456 5892 4458
rect 5858 4420 5892 4422
rect 5858 4334 5892 4354
rect 6008 4524 6042 4542
rect 6008 4456 6042 4458
rect 6008 4420 6042 4422
rect 6008 4334 6042 4354
rect 6166 4524 6200 4542
rect 6166 4456 6200 4458
rect 6166 4420 6200 4422
rect 6166 4334 6200 4354
rect 6360 4524 6394 4542
rect 6360 4456 6394 4458
rect 6360 4420 6394 4422
rect 6360 4334 6394 4354
rect 6518 4524 6552 4542
rect 6518 4456 6552 4458
rect 6518 4420 6552 4422
rect 6518 4334 6552 4354
rect 6668 4524 6702 4542
rect 6668 4456 6702 4458
rect 6668 4420 6702 4422
rect 6668 4334 6702 4354
rect 6826 4524 6860 4542
rect 6826 4456 6860 4458
rect 6826 4420 6860 4422
rect 6826 4334 6860 4354
rect 3670 4298 3704 4311
rect 3668 4295 3707 4298
rect 1773 4225 1807 4234
rect 2261 4227 2319 4239
rect 2625 4228 2703 4242
rect 2850 4237 2857 4271
rect 2891 4237 2898 4271
rect 3013 4237 3029 4271
rect 3063 4237 3079 4271
rect 3668 4261 3670 4295
rect 3704 4261 3707 4295
rect 3984 4289 4018 4302
rect 5628 4298 5662 4312
rect 3668 4259 3707 4261
rect 3982 4286 4021 4289
rect 3670 4245 3704 4259
rect 3982 4252 3984 4286
rect 4018 4252 4021 4286
rect 3982 4250 4021 4252
rect 4306 4281 4340 4296
rect 4306 4280 4341 4281
rect 2850 4230 2898 4237
rect 1255 4211 1318 4223
rect 2271 4221 2309 4227
rect 1410 4157 1444 4194
rect 556 4068 616 4084
rect 556 4044 565 4068
rect 606 4044 616 4068
rect 702 4068 762 4084
rect 702 4044 712 4068
rect 753 4044 762 4068
rect 846 4073 906 4090
rect 846 4050 856 4073
rect 897 4050 906 4073
rect 1000 4074 1060 4090
rect 1410 4086 1444 4123
rect 1568 4157 1602 4194
rect 1568 4086 1602 4123
rect 1698 4157 1732 4194
rect 1698 4086 1732 4123
rect 1856 4157 1890 4194
rect 1856 4086 1890 4123
rect 2030 4157 2064 4194
rect 2030 4086 2064 4123
rect 2188 4157 2222 4194
rect 2188 4086 2222 4123
rect 2352 4157 2420 4200
rect 2352 4123 2372 4157
rect 2406 4123 2420 4157
rect 1000 4050 1010 4074
rect 1051 4050 1060 4074
rect 540 4028 565 4044
rect 606 4028 632 4044
rect 540 4010 569 4028
rect 603 4010 632 4028
rect 686 4028 712 4044
rect 753 4028 778 4044
rect 686 4010 715 4028
rect 749 4010 778 4028
rect 830 4033 856 4050
rect 897 4033 922 4050
rect 830 4016 859 4033
rect 893 4016 922 4033
rect 984 4034 1010 4050
rect 1051 4034 1076 4050
rect 984 4016 1013 4034
rect 1047 4016 1076 4034
rect 1324 3980 1960 4044
rect 1324 3946 1353 3980
rect 1407 3946 1421 3980
rect 1479 3946 1489 3980
rect 1551 3946 1557 3980
rect 1623 3946 1625 3980
rect 1659 3946 1661 3980
rect 1727 3946 1733 3980
rect 1795 3946 1805 3980
rect 1863 3946 1877 3980
rect 1931 3946 1960 3980
rect 1324 3904 1960 3946
rect 2352 3955 2420 4123
rect 2530 4157 2564 4194
rect 2530 4086 2564 4123
rect 2352 3921 2369 3955
rect 2403 3921 2420 3955
rect 2352 3904 2420 3921
rect 2642 3859 2696 4228
rect 2857 4221 2891 4230
rect 3019 4227 3073 4237
rect 3984 4236 4018 4250
rect 4340 4246 4341 4280
rect 4621 4264 4637 4298
rect 4671 4264 4687 4298
rect 5626 4296 5666 4298
rect 5626 4262 5628 4296
rect 5662 4262 5666 4296
rect 5942 4290 5976 4302
rect 5626 4260 5666 4262
rect 5940 4286 5980 4290
rect 5628 4246 5662 4260
rect 5940 4252 5942 4286
rect 5976 4252 5980 4286
rect 5940 4250 5980 4252
rect 6264 4282 6298 4296
rect 6264 4280 6300 4282
rect 4306 4230 4340 4246
rect 5942 4236 5976 4250
rect 6298 4246 6300 4280
rect 6580 4264 6596 4298
rect 6630 4264 6646 4298
rect 6264 4230 6298 4246
rect 2776 4157 2810 4194
rect 2776 4086 2810 4123
rect 2934 4157 2968 4194
rect 2934 4086 2968 4123
rect 3120 4157 3154 4194
rect 3120 4086 3154 4123
rect 3278 4157 3312 4194
rect 3278 4086 3312 4123
rect 3742 4167 3776 4204
rect 3742 4096 3776 4133
rect 3900 4167 3934 4204
rect 3900 4096 3934 4133
rect 4050 4167 4084 4204
rect 4050 4096 4084 4133
rect 4208 4167 4242 4204
rect 4208 4096 4242 4133
rect 4402 4169 4436 4206
rect 4402 4098 4436 4135
rect 4560 4169 4594 4206
rect 4560 4098 4594 4135
rect 4710 4169 4744 4206
rect 4710 4098 4744 4135
rect 4868 4169 4902 4206
rect 4868 4098 4902 4135
rect 5700 4168 5734 4204
rect 5700 4096 5734 4134
rect 5858 4168 5892 4204
rect 5858 4096 5892 4134
rect 6008 4168 6042 4204
rect 6008 4096 6042 4134
rect 6166 4168 6200 4204
rect 6166 4096 6200 4134
rect 6360 4170 6394 4206
rect 6360 4098 6394 4136
rect 6518 4170 6552 4206
rect 6518 4098 6552 4136
rect 6668 4170 6702 4206
rect 6668 4098 6702 4136
rect 6826 4170 6860 4206
rect 6826 4098 6860 4136
rect 3704 3991 4244 4044
rect 3704 3957 3741 3991
rect 3787 3957 3813 3991
rect 3855 3957 3885 3991
rect 3923 3957 3957 3991
rect 3991 3957 4025 3991
rect 4063 3957 4093 3991
rect 4135 3957 4161 3991
rect 4207 3957 4244 3991
rect 3704 3904 4244 3957
rect 5662 3992 6202 4044
rect 5662 3958 5700 3992
rect 5746 3958 5772 3992
rect 5814 3958 5844 3992
rect 5882 3958 5916 3992
rect 5950 3958 5984 3992
rect 6022 3958 6052 3992
rect 6094 3958 6120 3992
rect 6166 3958 6202 3992
rect 5662 3904 6202 3958
rect 1348 3454 1880 3506
rect 1348 3420 1383 3454
rect 1429 3420 1455 3454
rect 1497 3420 1527 3454
rect 1565 3420 1599 3454
rect 1633 3420 1667 3454
rect 1705 3420 1735 3454
rect 1777 3420 1803 3454
rect 1849 3420 1880 3454
rect 3724 3453 4264 3506
rect 540 3368 569 3384
rect 603 3368 632 3384
rect 540 3350 566 3368
rect 607 3350 632 3368
rect 686 3368 715 3384
rect 749 3368 778 3384
rect 686 3350 710 3368
rect 751 3350 778 3368
rect 830 3373 859 3390
rect 893 3373 922 3390
rect 830 3356 856 3373
rect 897 3356 922 3373
rect 984 3373 1013 3390
rect 1047 3373 1076 3390
rect 984 3356 1009 3373
rect 1050 3356 1076 3373
rect 1348 3366 1880 3420
rect 2627 3373 3073 3427
rect 556 3328 566 3350
rect 607 3328 616 3350
rect 556 3310 616 3328
rect 702 3328 710 3350
rect 751 3328 762 3350
rect 702 3310 762 3328
rect 846 3333 856 3356
rect 897 3333 906 3356
rect 846 3316 906 3333
rect 1000 3333 1009 3356
rect 1050 3333 1060 3356
rect 1000 3316 1060 3333
rect 1410 3285 1444 3304
rect 1410 3217 1444 3219
rect 1410 3181 1444 3183
rect 1410 3096 1444 3115
rect 1568 3285 1602 3304
rect 1568 3217 1602 3219
rect 1568 3181 1602 3183
rect 1568 3096 1602 3115
rect 1698 3285 1732 3304
rect 1698 3217 1732 3219
rect 1698 3181 1732 3183
rect 1698 3096 1732 3115
rect 1856 3285 1890 3304
rect 1856 3217 1890 3219
rect 1856 3181 1890 3183
rect 1856 3096 1890 3115
rect 2030 3285 2064 3304
rect 2030 3217 2064 3219
rect 2030 3181 2064 3183
rect 2030 3096 2064 3115
rect 2188 3285 2222 3304
rect 2188 3217 2222 3219
rect 2188 3181 2222 3183
rect 2188 3096 2222 3115
rect 2372 3285 2406 3304
rect 2372 3217 2406 3219
rect 2372 3181 2406 3183
rect 2372 3096 2406 3115
rect 2530 3285 2564 3304
rect 2627 3223 2681 3373
rect 2776 3285 2810 3304
rect 2530 3217 2564 3219
rect 2530 3181 2564 3183
rect 2530 3096 2564 3115
rect 2625 3201 2703 3223
rect 2625 3167 2647 3201
rect 2681 3167 2703 3201
rect 1255 3066 1318 3078
rect 1251 3047 1322 3066
rect 2625 3063 2703 3167
rect 2776 3217 2810 3219
rect 2776 3181 2810 3183
rect 2776 3096 2810 3115
rect 2934 3285 2968 3304
rect 2934 3217 2968 3219
rect 2934 3181 2968 3183
rect 2934 3096 2968 3115
rect 1773 3054 1807 3063
rect 2271 3057 2309 3063
rect 1251 3013 1269 3047
rect 1303 3013 1322 3047
rect 1251 2995 1322 3013
rect 1766 3047 1814 3054
rect 1766 3013 1773 3047
rect 1807 3013 1814 3047
rect 1766 3006 1814 3013
rect 2261 3045 2319 3057
rect 2261 3011 2273 3045
rect 2307 3011 2319 3045
rect 2615 3055 2713 3063
rect 2615 3021 2647 3055
rect 2681 3021 2713 3055
rect 2857 3050 2891 3059
rect 2615 3014 2713 3021
rect 2850 3043 2898 3050
rect 3019 3043 3073 3373
rect 3724 3419 3773 3453
rect 3831 3419 3841 3453
rect 3903 3419 3909 3453
rect 3975 3419 3977 3453
rect 4011 3419 4013 3453
rect 4079 3419 4085 3453
rect 4147 3419 4157 3453
rect 4215 3419 4264 3453
rect 3724 3366 4264 3419
rect 5682 3452 6222 3506
rect 5682 3418 5732 3452
rect 5790 3418 5800 3452
rect 5862 3418 5868 3452
rect 5934 3418 5936 3452
rect 5970 3418 5972 3452
rect 6038 3418 6044 3452
rect 6106 3418 6116 3452
rect 6174 3418 6222 3452
rect 5682 3366 6222 3418
rect 3120 3285 3154 3304
rect 3120 3217 3154 3219
rect 3120 3181 3154 3183
rect 3120 3096 3154 3115
rect 3278 3285 3312 3304
rect 3278 3217 3312 3219
rect 3278 3181 3312 3183
rect 3278 3096 3312 3115
rect 3742 3295 3776 3314
rect 3742 3227 3776 3229
rect 3742 3191 3776 3193
rect 3742 3106 3776 3125
rect 3900 3295 3934 3314
rect 3900 3227 3934 3229
rect 3900 3191 3934 3193
rect 3900 3106 3934 3125
rect 4050 3295 4084 3314
rect 4050 3227 4084 3229
rect 4050 3191 4084 3193
rect 4050 3106 4084 3125
rect 4208 3295 4242 3314
rect 4208 3227 4242 3229
rect 4208 3191 4242 3193
rect 4208 3106 4242 3125
rect 4402 3295 4436 3314
rect 4402 3227 4436 3229
rect 4402 3191 4436 3193
rect 4402 3106 4436 3125
rect 4560 3295 4594 3314
rect 4560 3227 4594 3229
rect 4560 3191 4594 3193
rect 4560 3106 4594 3125
rect 4710 3295 4744 3314
rect 4710 3227 4744 3229
rect 4710 3191 4744 3193
rect 4710 3106 4744 3125
rect 4868 3295 4902 3314
rect 4868 3227 4902 3229
rect 4868 3191 4902 3193
rect 4868 3106 4902 3125
rect 5700 3296 5734 3314
rect 5700 3228 5734 3230
rect 5700 3192 5734 3194
rect 5700 3106 5734 3126
rect 5858 3296 5892 3314
rect 5858 3228 5892 3230
rect 5858 3192 5892 3194
rect 5858 3106 5892 3126
rect 6008 3296 6042 3314
rect 6008 3228 6042 3230
rect 6008 3192 6042 3194
rect 6008 3106 6042 3126
rect 6166 3296 6200 3314
rect 6166 3228 6200 3230
rect 6166 3192 6200 3194
rect 6166 3106 6200 3126
rect 6360 3296 6394 3314
rect 6360 3228 6394 3230
rect 6360 3192 6394 3194
rect 6360 3106 6394 3126
rect 6518 3296 6552 3314
rect 6518 3228 6552 3230
rect 6518 3192 6552 3194
rect 6518 3106 6552 3126
rect 6668 3296 6702 3314
rect 6668 3228 6702 3230
rect 6668 3192 6702 3194
rect 6668 3106 6702 3126
rect 6826 3296 6860 3314
rect 6826 3228 6860 3230
rect 6826 3192 6860 3194
rect 6826 3106 6860 3126
rect 3670 3070 3704 3083
rect 3668 3067 3707 3070
rect 1773 2997 1807 3006
rect 2261 2999 2319 3011
rect 2625 3000 2703 3014
rect 2850 3009 2857 3043
rect 2891 3009 2898 3043
rect 3013 3009 3029 3043
rect 3063 3009 3079 3043
rect 3668 3033 3670 3067
rect 3704 3033 3707 3067
rect 3984 3061 4018 3074
rect 5628 3070 5662 3084
rect 3668 3031 3707 3033
rect 3982 3058 4021 3061
rect 3670 3017 3704 3031
rect 3982 3024 3984 3058
rect 4018 3024 4021 3058
rect 3982 3022 4021 3024
rect 4306 3053 4340 3068
rect 4306 3052 4341 3053
rect 2850 3002 2898 3009
rect 1255 2983 1318 2995
rect 2271 2993 2309 2999
rect 1410 2929 1444 2966
rect 556 2840 616 2856
rect 556 2816 565 2840
rect 606 2816 616 2840
rect 702 2840 762 2856
rect 702 2816 712 2840
rect 753 2816 762 2840
rect 846 2845 906 2862
rect 846 2822 856 2845
rect 897 2822 906 2845
rect 1000 2846 1060 2862
rect 1410 2858 1444 2895
rect 1568 2929 1602 2966
rect 1568 2858 1602 2895
rect 1698 2929 1732 2966
rect 1698 2858 1732 2895
rect 1856 2929 1890 2966
rect 1856 2858 1890 2895
rect 2030 2929 2064 2966
rect 2030 2858 2064 2895
rect 2188 2929 2222 2966
rect 2188 2858 2222 2895
rect 2352 2929 2420 2972
rect 2352 2895 2372 2929
rect 2406 2895 2420 2929
rect 1000 2822 1010 2846
rect 1051 2822 1060 2846
rect 540 2800 565 2816
rect 606 2800 632 2816
rect 540 2782 569 2800
rect 603 2782 632 2800
rect 686 2800 712 2816
rect 753 2800 778 2816
rect 686 2782 715 2800
rect 749 2782 778 2800
rect 830 2805 856 2822
rect 897 2805 922 2822
rect 830 2788 859 2805
rect 893 2788 922 2805
rect 984 2806 1010 2822
rect 1051 2806 1076 2822
rect 984 2788 1013 2806
rect 1047 2788 1076 2806
rect 1324 2752 1960 2816
rect 1324 2718 1353 2752
rect 1407 2718 1421 2752
rect 1479 2718 1489 2752
rect 1551 2718 1557 2752
rect 1623 2718 1625 2752
rect 1659 2718 1661 2752
rect 1727 2718 1733 2752
rect 1795 2718 1805 2752
rect 1863 2718 1877 2752
rect 1931 2718 1960 2752
rect 1324 2676 1960 2718
rect 2352 2727 2420 2895
rect 2530 2929 2564 2966
rect 2530 2858 2564 2895
rect 2352 2693 2369 2727
rect 2403 2693 2420 2727
rect 2352 2676 2420 2693
rect 2642 2631 2696 3000
rect 2857 2993 2891 3002
rect 3019 2999 3073 3009
rect 3984 3008 4018 3022
rect 4340 3018 4341 3052
rect 4621 3036 4637 3070
rect 4671 3036 4687 3070
rect 5626 3068 5666 3070
rect 5626 3034 5628 3068
rect 5662 3034 5666 3068
rect 5942 3062 5976 3074
rect 5626 3032 5666 3034
rect 5940 3058 5980 3062
rect 5628 3018 5662 3032
rect 5940 3024 5942 3058
rect 5976 3024 5980 3058
rect 5940 3022 5980 3024
rect 6264 3054 6298 3068
rect 6264 3052 6300 3054
rect 4306 3002 4340 3018
rect 5942 3008 5976 3022
rect 6298 3018 6300 3052
rect 6580 3036 6596 3070
rect 6630 3036 6646 3070
rect 6264 3002 6298 3018
rect 2776 2929 2810 2966
rect 2776 2858 2810 2895
rect 2934 2929 2968 2966
rect 2934 2858 2968 2895
rect 3120 2929 3154 2966
rect 3120 2858 3154 2895
rect 3278 2929 3312 2966
rect 3278 2858 3312 2895
rect 3742 2939 3776 2976
rect 3742 2868 3776 2905
rect 3900 2939 3934 2976
rect 3900 2868 3934 2905
rect 4050 2939 4084 2976
rect 4050 2868 4084 2905
rect 4208 2939 4242 2976
rect 4208 2868 4242 2905
rect 4402 2941 4436 2978
rect 4402 2870 4436 2907
rect 4560 2941 4594 2978
rect 4560 2870 4594 2907
rect 4710 2941 4744 2978
rect 4710 2870 4744 2907
rect 4868 2941 4902 2978
rect 4868 2870 4902 2907
rect 5700 2940 5734 2976
rect 5700 2868 5734 2906
rect 5858 2940 5892 2976
rect 5858 2868 5892 2906
rect 6008 2940 6042 2976
rect 6008 2868 6042 2906
rect 6166 2940 6200 2976
rect 6166 2868 6200 2906
rect 6360 2942 6394 2978
rect 6360 2870 6394 2908
rect 6518 2942 6552 2978
rect 6518 2870 6552 2908
rect 6668 2942 6702 2978
rect 6668 2870 6702 2908
rect 6826 2942 6860 2978
rect 6826 2870 6860 2908
rect 3704 2763 4244 2816
rect 3704 2729 3741 2763
rect 3787 2729 3813 2763
rect 3855 2729 3885 2763
rect 3923 2729 3957 2763
rect 3991 2729 4025 2763
rect 4063 2729 4093 2763
rect 4135 2729 4161 2763
rect 4207 2729 4244 2763
rect 3704 2676 4244 2729
rect 5662 2764 6202 2816
rect 5662 2730 5700 2764
rect 5746 2730 5772 2764
rect 5814 2730 5844 2764
rect 5882 2730 5916 2764
rect 5950 2730 5984 2764
rect 6022 2730 6052 2764
rect 6094 2730 6120 2764
rect 6166 2730 6202 2764
rect 5662 2676 6202 2730
rect 1348 2226 1880 2278
rect 1348 2192 1383 2226
rect 1429 2192 1455 2226
rect 1497 2192 1527 2226
rect 1565 2192 1599 2226
rect 1633 2192 1667 2226
rect 1705 2192 1735 2226
rect 1777 2192 1803 2226
rect 1849 2192 1880 2226
rect 3724 2225 4264 2278
rect 540 2140 569 2156
rect 603 2140 632 2156
rect 540 2122 566 2140
rect 607 2122 632 2140
rect 686 2140 715 2156
rect 749 2140 778 2156
rect 686 2122 710 2140
rect 751 2122 778 2140
rect 830 2145 859 2162
rect 893 2145 922 2162
rect 830 2128 856 2145
rect 897 2128 922 2145
rect 984 2145 1013 2162
rect 1047 2145 1076 2162
rect 984 2128 1009 2145
rect 1050 2128 1076 2145
rect 1348 2138 1880 2192
rect 2627 2145 3073 2199
rect 556 2100 566 2122
rect 607 2100 616 2122
rect 556 2082 616 2100
rect 702 2100 710 2122
rect 751 2100 762 2122
rect 702 2082 762 2100
rect 846 2105 856 2128
rect 897 2105 906 2128
rect 846 2088 906 2105
rect 1000 2105 1009 2128
rect 1050 2105 1060 2128
rect 1000 2088 1060 2105
rect 1410 2057 1444 2076
rect 1410 1989 1444 1991
rect 1410 1953 1444 1955
rect 1410 1868 1444 1887
rect 1568 2057 1602 2076
rect 1568 1989 1602 1991
rect 1568 1953 1602 1955
rect 1568 1868 1602 1887
rect 1698 2057 1732 2076
rect 1698 1989 1732 1991
rect 1698 1953 1732 1955
rect 1698 1868 1732 1887
rect 1856 2057 1890 2076
rect 1856 1989 1890 1991
rect 1856 1953 1890 1955
rect 1856 1868 1890 1887
rect 2030 2057 2064 2076
rect 2030 1989 2064 1991
rect 2030 1953 2064 1955
rect 2030 1868 2064 1887
rect 2188 2057 2222 2076
rect 2188 1989 2222 1991
rect 2188 1953 2222 1955
rect 2188 1868 2222 1887
rect 2372 2057 2406 2076
rect 2372 1989 2406 1991
rect 2372 1953 2406 1955
rect 2372 1868 2406 1887
rect 2530 2057 2564 2076
rect 2627 1995 2681 2145
rect 2776 2057 2810 2076
rect 2530 1989 2564 1991
rect 2530 1953 2564 1955
rect 2530 1868 2564 1887
rect 2625 1973 2703 1995
rect 2625 1939 2647 1973
rect 2681 1939 2703 1973
rect 1255 1838 1318 1850
rect 1251 1819 1322 1838
rect 2625 1835 2703 1939
rect 2776 1989 2810 1991
rect 2776 1953 2810 1955
rect 2776 1868 2810 1887
rect 2934 2057 2968 2076
rect 2934 1989 2968 1991
rect 2934 1953 2968 1955
rect 2934 1868 2968 1887
rect 1773 1826 1807 1835
rect 2271 1829 2309 1835
rect 1251 1785 1269 1819
rect 1303 1785 1322 1819
rect 1251 1767 1322 1785
rect 1766 1819 1814 1826
rect 1766 1785 1773 1819
rect 1807 1785 1814 1819
rect 1766 1778 1814 1785
rect 2261 1817 2319 1829
rect 2261 1783 2273 1817
rect 2307 1783 2319 1817
rect 2615 1827 2713 1835
rect 2615 1793 2647 1827
rect 2681 1793 2713 1827
rect 2857 1822 2891 1831
rect 2615 1786 2713 1793
rect 2850 1815 2898 1822
rect 3019 1815 3073 2145
rect 3724 2191 3773 2225
rect 3831 2191 3841 2225
rect 3903 2191 3909 2225
rect 3975 2191 3977 2225
rect 4011 2191 4013 2225
rect 4079 2191 4085 2225
rect 4147 2191 4157 2225
rect 4215 2191 4264 2225
rect 3724 2138 4264 2191
rect 5682 2224 6222 2278
rect 5682 2190 5732 2224
rect 5790 2190 5800 2224
rect 5862 2190 5868 2224
rect 5934 2190 5936 2224
rect 5970 2190 5972 2224
rect 6038 2190 6044 2224
rect 6106 2190 6116 2224
rect 6174 2190 6222 2224
rect 5682 2138 6222 2190
rect 3120 2057 3154 2076
rect 3120 1989 3154 1991
rect 3120 1953 3154 1955
rect 3120 1868 3154 1887
rect 3278 2057 3312 2076
rect 3278 1989 3312 1991
rect 3278 1953 3312 1955
rect 3278 1868 3312 1887
rect 3742 2067 3776 2086
rect 3742 1999 3776 2001
rect 3742 1963 3776 1965
rect 3742 1878 3776 1897
rect 3900 2067 3934 2086
rect 3900 1999 3934 2001
rect 3900 1963 3934 1965
rect 3900 1878 3934 1897
rect 4050 2067 4084 2086
rect 4050 1999 4084 2001
rect 4050 1963 4084 1965
rect 4050 1878 4084 1897
rect 4208 2067 4242 2086
rect 4208 1999 4242 2001
rect 4208 1963 4242 1965
rect 4208 1878 4242 1897
rect 4402 2067 4436 2086
rect 4402 1999 4436 2001
rect 4402 1963 4436 1965
rect 4402 1878 4436 1897
rect 4560 2067 4594 2086
rect 4560 1999 4594 2001
rect 4560 1963 4594 1965
rect 4560 1878 4594 1897
rect 4710 2067 4744 2086
rect 4710 1999 4744 2001
rect 4710 1963 4744 1965
rect 4710 1878 4744 1897
rect 4868 2067 4902 2086
rect 4868 1999 4902 2001
rect 4868 1963 4902 1965
rect 4868 1878 4902 1897
rect 5700 2068 5734 2086
rect 5700 2000 5734 2002
rect 5700 1964 5734 1966
rect 5700 1878 5734 1898
rect 5858 2068 5892 2086
rect 5858 2000 5892 2002
rect 5858 1964 5892 1966
rect 5858 1878 5892 1898
rect 6008 2068 6042 2086
rect 6008 2000 6042 2002
rect 6008 1964 6042 1966
rect 6008 1878 6042 1898
rect 6166 2068 6200 2086
rect 6166 2000 6200 2002
rect 6166 1964 6200 1966
rect 6166 1878 6200 1898
rect 6360 2068 6394 2086
rect 6360 2000 6394 2002
rect 6360 1964 6394 1966
rect 6360 1878 6394 1898
rect 6518 2068 6552 2086
rect 6518 2000 6552 2002
rect 6518 1964 6552 1966
rect 6518 1878 6552 1898
rect 6668 2068 6702 2086
rect 6668 2000 6702 2002
rect 6668 1964 6702 1966
rect 6668 1878 6702 1898
rect 6826 2068 6860 2086
rect 6826 2000 6860 2002
rect 6826 1964 6860 1966
rect 6826 1878 6860 1898
rect 3670 1842 3704 1855
rect 3668 1839 3707 1842
rect 1773 1769 1807 1778
rect 2261 1771 2319 1783
rect 2625 1772 2703 1786
rect 2850 1781 2857 1815
rect 2891 1781 2898 1815
rect 3013 1781 3029 1815
rect 3063 1781 3079 1815
rect 3668 1805 3670 1839
rect 3704 1805 3707 1839
rect 3984 1833 4018 1846
rect 5628 1842 5662 1856
rect 3668 1803 3707 1805
rect 3982 1830 4021 1833
rect 3670 1789 3704 1803
rect 3982 1796 3984 1830
rect 4018 1796 4021 1830
rect 3982 1794 4021 1796
rect 4306 1825 4340 1840
rect 4306 1824 4341 1825
rect 2850 1774 2898 1781
rect 1255 1755 1318 1767
rect 2271 1765 2309 1771
rect 1410 1701 1444 1738
rect 556 1612 616 1628
rect 556 1588 565 1612
rect 606 1588 616 1612
rect 702 1612 762 1628
rect 702 1588 712 1612
rect 753 1588 762 1612
rect 846 1617 906 1634
rect 846 1594 856 1617
rect 897 1594 906 1617
rect 1000 1618 1060 1634
rect 1410 1630 1444 1667
rect 1568 1701 1602 1738
rect 1568 1630 1602 1667
rect 1698 1701 1732 1738
rect 1698 1630 1732 1667
rect 1856 1701 1890 1738
rect 1856 1630 1890 1667
rect 2030 1701 2064 1738
rect 2030 1630 2064 1667
rect 2188 1701 2222 1738
rect 2188 1630 2222 1667
rect 2352 1701 2420 1744
rect 2352 1667 2372 1701
rect 2406 1667 2420 1701
rect 1000 1594 1010 1618
rect 1051 1594 1060 1618
rect 540 1572 565 1588
rect 606 1572 632 1588
rect 540 1554 569 1572
rect 603 1554 632 1572
rect 686 1572 712 1588
rect 753 1572 778 1588
rect 686 1554 715 1572
rect 749 1554 778 1572
rect 830 1577 856 1594
rect 897 1577 922 1594
rect 830 1560 859 1577
rect 893 1560 922 1577
rect 984 1578 1010 1594
rect 1051 1578 1076 1594
rect 984 1560 1013 1578
rect 1047 1560 1076 1578
rect 1324 1524 1960 1588
rect 1324 1490 1353 1524
rect 1407 1490 1421 1524
rect 1479 1490 1489 1524
rect 1551 1490 1557 1524
rect 1623 1490 1625 1524
rect 1659 1490 1661 1524
rect 1727 1490 1733 1524
rect 1795 1490 1805 1524
rect 1863 1490 1877 1524
rect 1931 1490 1960 1524
rect 1324 1448 1960 1490
rect 2352 1499 2420 1667
rect 2530 1701 2564 1738
rect 2530 1630 2564 1667
rect 2352 1465 2369 1499
rect 2403 1465 2420 1499
rect 2352 1448 2420 1465
rect 2642 1403 2696 1772
rect 2857 1765 2891 1774
rect 3019 1771 3073 1781
rect 3984 1780 4018 1794
rect 4340 1790 4341 1824
rect 4621 1808 4637 1842
rect 4671 1808 4687 1842
rect 5626 1840 5666 1842
rect 5626 1806 5628 1840
rect 5662 1806 5666 1840
rect 5942 1834 5976 1846
rect 5626 1804 5666 1806
rect 5940 1830 5980 1834
rect 5628 1790 5662 1804
rect 5940 1796 5942 1830
rect 5976 1796 5980 1830
rect 5940 1794 5980 1796
rect 6264 1826 6298 1840
rect 6264 1824 6300 1826
rect 4306 1774 4340 1790
rect 5942 1780 5976 1794
rect 6298 1790 6300 1824
rect 6580 1808 6596 1842
rect 6630 1808 6646 1842
rect 6264 1774 6298 1790
rect 2776 1701 2810 1738
rect 2776 1630 2810 1667
rect 2934 1701 2968 1738
rect 2934 1630 2968 1667
rect 3120 1701 3154 1738
rect 3120 1630 3154 1667
rect 3278 1701 3312 1738
rect 3278 1630 3312 1667
rect 3742 1711 3776 1748
rect 3742 1640 3776 1677
rect 3900 1711 3934 1748
rect 3900 1640 3934 1677
rect 4050 1711 4084 1748
rect 4050 1640 4084 1677
rect 4208 1711 4242 1748
rect 4208 1640 4242 1677
rect 4402 1713 4436 1750
rect 4402 1642 4436 1679
rect 4560 1713 4594 1750
rect 4560 1642 4594 1679
rect 4710 1713 4744 1750
rect 4710 1642 4744 1679
rect 4868 1713 4902 1750
rect 4868 1642 4902 1679
rect 5700 1712 5734 1748
rect 5700 1640 5734 1678
rect 5858 1712 5892 1748
rect 5858 1640 5892 1678
rect 6008 1712 6042 1748
rect 6008 1640 6042 1678
rect 6166 1712 6200 1748
rect 6166 1640 6200 1678
rect 6360 1714 6394 1750
rect 6360 1642 6394 1680
rect 6518 1714 6552 1750
rect 6518 1642 6552 1680
rect 6668 1714 6702 1750
rect 6668 1642 6702 1680
rect 6826 1714 6860 1750
rect 6826 1642 6860 1680
rect 3704 1535 4244 1588
rect 3704 1501 3741 1535
rect 3787 1501 3813 1535
rect 3855 1501 3885 1535
rect 3923 1501 3957 1535
rect 3991 1501 4025 1535
rect 4063 1501 4093 1535
rect 4135 1501 4161 1535
rect 4207 1501 4244 1535
rect 3704 1448 4244 1501
rect 5662 1536 6202 1588
rect 5662 1502 5700 1536
rect 5746 1502 5772 1536
rect 5814 1502 5844 1536
rect 5882 1502 5916 1536
rect 5950 1502 5984 1536
rect 6022 1502 6052 1536
rect 6094 1502 6120 1536
rect 6166 1502 6202 1536
rect 5662 1448 6202 1502
rect 1348 998 1880 1050
rect 1348 964 1383 998
rect 1429 964 1455 998
rect 1497 964 1527 998
rect 1565 964 1599 998
rect 1633 964 1667 998
rect 1705 964 1735 998
rect 1777 964 1803 998
rect 1849 964 1880 998
rect 3724 997 4264 1050
rect 540 912 569 928
rect 603 912 632 928
rect 540 894 566 912
rect 607 894 632 912
rect 686 912 715 928
rect 749 912 778 928
rect 686 894 710 912
rect 751 894 778 912
rect 830 917 859 934
rect 893 917 922 934
rect 830 900 856 917
rect 897 900 922 917
rect 984 917 1013 934
rect 1047 917 1076 934
rect 984 900 1009 917
rect 1050 900 1076 917
rect 1348 910 1880 964
rect 2627 917 3073 971
rect 556 872 566 894
rect 607 872 616 894
rect 556 854 616 872
rect 702 872 710 894
rect 751 872 762 894
rect 702 854 762 872
rect 846 877 856 900
rect 897 877 906 900
rect 846 860 906 877
rect 1000 877 1009 900
rect 1050 877 1060 900
rect 1000 860 1060 877
rect 1410 829 1444 848
rect 1410 761 1444 763
rect 1410 725 1444 727
rect 1410 640 1444 659
rect 1568 829 1602 848
rect 1568 761 1602 763
rect 1568 725 1602 727
rect 1568 640 1602 659
rect 1698 829 1732 848
rect 1698 761 1732 763
rect 1698 725 1732 727
rect 1698 640 1732 659
rect 1856 829 1890 848
rect 1856 761 1890 763
rect 1856 725 1890 727
rect 1856 640 1890 659
rect 2030 829 2064 848
rect 2030 761 2064 763
rect 2030 725 2064 727
rect 2030 640 2064 659
rect 2188 829 2222 848
rect 2188 761 2222 763
rect 2188 725 2222 727
rect 2188 640 2222 659
rect 2372 829 2406 848
rect 2372 761 2406 763
rect 2372 725 2406 727
rect 2372 640 2406 659
rect 2530 829 2564 848
rect 2627 767 2681 917
rect 2776 829 2810 848
rect 2530 761 2564 763
rect 2530 725 2564 727
rect 2530 640 2564 659
rect 2625 745 2703 767
rect 2625 711 2647 745
rect 2681 711 2703 745
rect 1255 610 1318 622
rect 1251 591 1322 610
rect 2625 607 2703 711
rect 2776 761 2810 763
rect 2776 725 2810 727
rect 2776 640 2810 659
rect 2934 829 2968 848
rect 2934 761 2968 763
rect 2934 725 2968 727
rect 2934 640 2968 659
rect 1773 598 1807 607
rect 2271 601 2309 607
rect 1251 557 1269 591
rect 1303 557 1322 591
rect 1251 539 1322 557
rect 1766 591 1814 598
rect 1766 557 1773 591
rect 1807 557 1814 591
rect 1766 550 1814 557
rect 2261 589 2319 601
rect 2261 555 2273 589
rect 2307 555 2319 589
rect 2615 599 2713 607
rect 2615 565 2647 599
rect 2681 565 2713 599
rect 2857 594 2891 603
rect 2615 558 2713 565
rect 2850 587 2898 594
rect 3019 587 3073 917
rect 3724 963 3773 997
rect 3831 963 3841 997
rect 3903 963 3909 997
rect 3975 963 3977 997
rect 4011 963 4013 997
rect 4079 963 4085 997
rect 4147 963 4157 997
rect 4215 963 4264 997
rect 3724 910 4264 963
rect 3120 829 3154 848
rect 3120 761 3154 763
rect 3120 725 3154 727
rect 3120 640 3154 659
rect 3278 829 3312 848
rect 3278 761 3312 763
rect 3278 725 3312 727
rect 3278 640 3312 659
rect 3742 839 3776 858
rect 3742 771 3776 773
rect 3742 735 3776 737
rect 3742 650 3776 669
rect 3900 839 3934 858
rect 3900 771 3934 773
rect 3900 735 3934 737
rect 3900 650 3934 669
rect 4050 839 4084 858
rect 4050 771 4084 773
rect 4050 735 4084 737
rect 4050 650 4084 669
rect 4208 839 4242 858
rect 4208 771 4242 773
rect 4208 735 4242 737
rect 4208 650 4242 669
rect 4402 839 4436 858
rect 4402 771 4436 773
rect 4402 735 4436 737
rect 4402 650 4436 669
rect 4560 839 4594 858
rect 4560 771 4594 773
rect 4560 735 4594 737
rect 4560 650 4594 669
rect 4710 839 4744 858
rect 4710 771 4744 773
rect 4710 735 4744 737
rect 4710 650 4744 669
rect 4868 839 4902 858
rect 4868 771 4902 773
rect 4868 735 4902 737
rect 4868 650 4902 669
rect 3670 614 3704 627
rect 3668 611 3707 614
rect 1773 541 1807 550
rect 2261 543 2319 555
rect 2625 544 2703 558
rect 2850 553 2857 587
rect 2891 553 2898 587
rect 3013 553 3029 587
rect 3063 553 3079 587
rect 3668 577 3670 611
rect 3704 577 3707 611
rect 3984 605 4018 618
rect 3668 575 3707 577
rect 3982 602 4021 605
rect 3670 561 3704 575
rect 3982 568 3984 602
rect 4018 568 4021 602
rect 3982 566 4021 568
rect 4306 597 4340 612
rect 4306 596 4341 597
rect 2850 546 2898 553
rect 1255 527 1318 539
rect 2271 537 2309 543
rect 1410 473 1444 510
rect 556 384 616 400
rect 556 360 565 384
rect 606 360 616 384
rect 702 384 762 400
rect 702 360 712 384
rect 753 360 762 384
rect 846 389 906 406
rect 846 366 856 389
rect 897 366 906 389
rect 1000 390 1060 406
rect 1410 402 1444 439
rect 1568 473 1602 510
rect 1568 402 1602 439
rect 1698 473 1732 510
rect 1698 402 1732 439
rect 1856 473 1890 510
rect 1856 402 1890 439
rect 2030 473 2064 510
rect 2030 402 2064 439
rect 2188 473 2222 510
rect 2188 402 2222 439
rect 2352 473 2420 516
rect 2352 439 2372 473
rect 2406 439 2420 473
rect 1000 366 1010 390
rect 1051 366 1060 390
rect 540 344 565 360
rect 606 344 632 360
rect 540 326 569 344
rect 603 326 632 344
rect 686 344 712 360
rect 753 344 778 360
rect 686 326 715 344
rect 749 326 778 344
rect 830 349 856 366
rect 897 349 922 366
rect 830 332 859 349
rect 893 332 922 349
rect 984 350 1010 366
rect 1051 350 1076 366
rect 984 332 1013 350
rect 1047 332 1076 350
rect 1324 296 1960 360
rect 1324 262 1353 296
rect 1407 262 1421 296
rect 1479 262 1489 296
rect 1551 262 1557 296
rect 1623 262 1625 296
rect 1659 262 1661 296
rect 1727 262 1733 296
rect 1795 262 1805 296
rect 1863 262 1877 296
rect 1931 262 1960 296
rect 1324 220 1960 262
rect 2352 271 2420 439
rect 2530 473 2564 510
rect 2530 402 2564 439
rect 2352 237 2369 271
rect 2403 237 2420 271
rect 2352 220 2420 237
rect 2642 175 2696 544
rect 2857 537 2891 546
rect 3019 543 3073 553
rect 3984 552 4018 566
rect 4340 562 4341 596
rect 4621 580 4637 614
rect 4671 580 4687 614
rect 4306 546 4340 562
rect 2776 473 2810 510
rect 2776 402 2810 439
rect 2934 473 2968 510
rect 2934 402 2968 439
rect 3120 473 3154 510
rect 3120 402 3154 439
rect 3278 473 3312 510
rect 3278 402 3312 439
rect 3742 483 3776 520
rect 3742 412 3776 449
rect 3900 483 3934 520
rect 3900 412 3934 449
rect 4050 483 4084 520
rect 4050 412 4084 449
rect 4208 483 4242 520
rect 4208 412 4242 449
rect 4402 485 4436 522
rect 4402 414 4436 451
rect 4560 485 4594 522
rect 4560 414 4594 451
rect 4710 485 4744 522
rect 4710 414 4744 451
rect 4868 485 4902 522
rect 4868 414 4902 451
rect 3704 307 4244 360
rect 3704 273 3741 307
rect 3787 273 3813 307
rect 3855 273 3885 307
rect 3923 273 3957 307
rect 3991 273 4025 307
rect 4063 273 4093 307
rect 4135 273 4161 307
rect 4207 273 4244 307
rect 3704 220 4244 273
<< viali >>
rect 1383 19384 1395 19418
rect 1395 19384 1417 19418
rect 1455 19384 1463 19418
rect 1463 19384 1489 19418
rect 1527 19384 1531 19418
rect 1531 19384 1561 19418
rect 1599 19384 1633 19418
rect 1671 19384 1701 19418
rect 1701 19384 1705 19418
rect 1743 19384 1769 19418
rect 1769 19384 1777 19418
rect 1815 19384 1837 19418
rect 1837 19384 1849 19418
rect 566 19314 569 19332
rect 569 19314 603 19332
rect 603 19314 607 19332
rect 710 19314 715 19332
rect 715 19314 749 19332
rect 749 19314 751 19332
rect 856 19320 859 19337
rect 859 19320 893 19337
rect 893 19320 897 19337
rect 1009 19320 1013 19337
rect 1013 19320 1047 19337
rect 1047 19320 1050 19337
rect 566 19292 607 19314
rect 710 19292 751 19314
rect 856 19297 897 19320
rect 1009 19297 1050 19320
rect 1410 19215 1444 19217
rect 1410 19183 1444 19215
rect 1410 19113 1444 19145
rect 1410 19111 1444 19113
rect 1568 19215 1602 19217
rect 1568 19183 1602 19215
rect 1568 19113 1602 19145
rect 1568 19111 1602 19113
rect 1698 19215 1732 19217
rect 1698 19183 1732 19215
rect 1698 19113 1732 19145
rect 1698 19111 1732 19113
rect 1856 19215 1890 19217
rect 1856 19183 1890 19215
rect 1856 19113 1890 19145
rect 1856 19111 1890 19113
rect 2030 19215 2064 19217
rect 2030 19183 2064 19215
rect 2030 19113 2064 19145
rect 2030 19111 2064 19113
rect 2188 19215 2222 19217
rect 2188 19183 2222 19215
rect 2188 19113 2222 19145
rect 2188 19111 2222 19113
rect 2372 19215 2406 19217
rect 2372 19183 2406 19215
rect 2372 19113 2406 19145
rect 2372 19111 2406 19113
rect 2530 19215 2564 19217
rect 2530 19183 2564 19215
rect 2776 19215 2810 19217
rect 2530 19113 2564 19145
rect 2530 19111 2564 19113
rect 2647 19131 2681 19165
rect 2776 19183 2810 19215
rect 2776 19113 2810 19145
rect 2776 19111 2810 19113
rect 2934 19215 2968 19217
rect 2934 19183 2968 19215
rect 2934 19113 2968 19145
rect 2934 19111 2968 19113
rect 1269 18977 1303 19011
rect 1773 18977 1807 19011
rect 2273 18975 2307 19009
rect 3797 19383 3807 19417
rect 3807 19383 3831 19417
rect 3869 19383 3875 19417
rect 3875 19383 3903 19417
rect 3941 19383 3943 19417
rect 3943 19383 3975 19417
rect 4013 19383 4045 19417
rect 4045 19383 4047 19417
rect 4085 19383 4113 19417
rect 4113 19383 4119 19417
rect 4157 19383 4181 19417
rect 4181 19383 4191 19417
rect 5756 19382 5766 19416
rect 5766 19382 5790 19416
rect 5828 19382 5834 19416
rect 5834 19382 5862 19416
rect 5900 19382 5902 19416
rect 5902 19382 5934 19416
rect 5972 19382 6004 19416
rect 6004 19382 6006 19416
rect 6044 19382 6072 19416
rect 6072 19382 6078 19416
rect 6116 19382 6140 19416
rect 6140 19382 6150 19416
rect 3120 19215 3154 19217
rect 3120 19183 3154 19215
rect 3120 19113 3154 19145
rect 3120 19111 3154 19113
rect 3278 19215 3312 19217
rect 3278 19183 3312 19215
rect 3278 19113 3312 19145
rect 3278 19111 3312 19113
rect 3742 19225 3776 19227
rect 3742 19193 3776 19225
rect 3742 19123 3776 19155
rect 3742 19121 3776 19123
rect 3900 19225 3934 19227
rect 3900 19193 3934 19225
rect 3900 19123 3934 19155
rect 3900 19121 3934 19123
rect 4050 19225 4084 19227
rect 4050 19193 4084 19225
rect 4050 19123 4084 19155
rect 4050 19121 4084 19123
rect 4208 19225 4242 19227
rect 4208 19193 4242 19225
rect 4208 19123 4242 19155
rect 4208 19121 4242 19123
rect 4402 19225 4436 19227
rect 4402 19193 4436 19225
rect 4402 19123 4436 19155
rect 4402 19121 4436 19123
rect 4560 19225 4594 19227
rect 4560 19193 4594 19225
rect 4560 19123 4594 19155
rect 4560 19121 4594 19123
rect 4710 19225 4744 19227
rect 4710 19193 4744 19225
rect 4710 19123 4744 19155
rect 4710 19121 4744 19123
rect 4868 19225 4902 19227
rect 4868 19193 4902 19225
rect 4868 19123 4902 19155
rect 4868 19121 4902 19123
rect 5700 19226 5734 19228
rect 5700 19194 5734 19226
rect 5700 19124 5734 19156
rect 5700 19122 5734 19124
rect 5858 19226 5892 19228
rect 5858 19194 5892 19226
rect 5858 19124 5892 19156
rect 5858 19122 5892 19124
rect 6008 19226 6042 19228
rect 6008 19194 6042 19226
rect 6008 19124 6042 19156
rect 6008 19122 6042 19124
rect 6166 19226 6200 19228
rect 6166 19194 6200 19226
rect 6166 19124 6200 19156
rect 6166 19122 6200 19124
rect 6360 19226 6394 19228
rect 6360 19194 6394 19226
rect 6360 19124 6394 19156
rect 6360 19122 6394 19124
rect 6518 19226 6552 19228
rect 6518 19194 6552 19226
rect 6518 19124 6552 19156
rect 6518 19122 6552 19124
rect 6668 19226 6702 19228
rect 6668 19194 6702 19226
rect 6668 19124 6702 19156
rect 6668 19122 6702 19124
rect 6826 19226 6860 19228
rect 6826 19194 6860 19226
rect 6826 19124 6860 19156
rect 6826 19122 6860 19124
rect 2857 18973 2891 19007
rect 3670 18997 3704 19031
rect 3984 18988 4018 19022
rect 1410 18859 1444 18893
rect 565 18780 606 18804
rect 712 18780 753 18804
rect 856 18786 897 18809
rect 1568 18859 1602 18893
rect 1698 18859 1732 18893
rect 1856 18859 1890 18893
rect 2030 18859 2064 18893
rect 2188 18859 2222 18893
rect 2372 18859 2406 18893
rect 1010 18786 1051 18810
rect 565 18764 569 18780
rect 569 18764 603 18780
rect 603 18764 606 18780
rect 712 18764 715 18780
rect 715 18764 749 18780
rect 749 18764 753 18780
rect 856 18769 859 18786
rect 859 18769 893 18786
rect 893 18769 897 18786
rect 1010 18770 1013 18786
rect 1013 18770 1047 18786
rect 1047 18770 1051 18786
rect 1373 18682 1387 18716
rect 1387 18682 1407 18716
rect 1445 18682 1455 18716
rect 1455 18682 1479 18716
rect 1517 18682 1523 18716
rect 1523 18682 1551 18716
rect 1589 18682 1591 18716
rect 1591 18682 1623 18716
rect 1661 18682 1693 18716
rect 1693 18682 1695 18716
rect 1733 18682 1761 18716
rect 1761 18682 1767 18716
rect 1805 18682 1829 18716
rect 1829 18682 1839 18716
rect 1877 18682 1897 18716
rect 1897 18682 1911 18716
rect 2530 18859 2564 18893
rect 2369 18657 2403 18691
rect 4306 18982 4340 19016
rect 4637 19000 4671 19034
rect 5628 18998 5662 19032
rect 5942 18988 5976 19022
rect 6264 18982 6298 19016
rect 6596 19000 6630 19034
rect 2776 18859 2810 18893
rect 2934 18859 2968 18893
rect 3120 18859 3154 18893
rect 3278 18859 3312 18893
rect 3742 18869 3776 18903
rect 3900 18869 3934 18903
rect 4050 18869 4084 18903
rect 4208 18869 4242 18903
rect 4402 18871 4436 18905
rect 4560 18871 4594 18905
rect 4710 18871 4744 18905
rect 4868 18871 4902 18905
rect 5700 18870 5734 18904
rect 5858 18870 5892 18904
rect 6008 18870 6042 18904
rect 6166 18870 6200 18904
rect 6360 18872 6394 18906
rect 6518 18872 6552 18906
rect 6668 18872 6702 18906
rect 6826 18872 6860 18906
rect 3741 18693 3753 18727
rect 3753 18693 3775 18727
rect 3813 18693 3821 18727
rect 3821 18693 3847 18727
rect 3885 18693 3889 18727
rect 3889 18693 3919 18727
rect 3957 18693 3991 18727
rect 4029 18693 4059 18727
rect 4059 18693 4063 18727
rect 4101 18693 4127 18727
rect 4127 18693 4135 18727
rect 4173 18693 4195 18727
rect 4195 18693 4207 18727
rect 5700 18694 5712 18728
rect 5712 18694 5734 18728
rect 5772 18694 5780 18728
rect 5780 18694 5806 18728
rect 5844 18694 5848 18728
rect 5848 18694 5878 18728
rect 5916 18694 5950 18728
rect 5988 18694 6018 18728
rect 6018 18694 6022 18728
rect 6060 18694 6086 18728
rect 6086 18694 6094 18728
rect 6132 18694 6154 18728
rect 6154 18694 6166 18728
rect 2642 18541 2696 18595
rect 1383 18156 1395 18190
rect 1395 18156 1417 18190
rect 1455 18156 1463 18190
rect 1463 18156 1489 18190
rect 1527 18156 1531 18190
rect 1531 18156 1561 18190
rect 1599 18156 1633 18190
rect 1671 18156 1701 18190
rect 1701 18156 1705 18190
rect 1743 18156 1769 18190
rect 1769 18156 1777 18190
rect 1815 18156 1837 18190
rect 1837 18156 1849 18190
rect 566 18086 569 18104
rect 569 18086 603 18104
rect 603 18086 607 18104
rect 710 18086 715 18104
rect 715 18086 749 18104
rect 749 18086 751 18104
rect 856 18092 859 18109
rect 859 18092 893 18109
rect 893 18092 897 18109
rect 1009 18092 1013 18109
rect 1013 18092 1047 18109
rect 1047 18092 1050 18109
rect 566 18064 607 18086
rect 710 18064 751 18086
rect 856 18069 897 18092
rect 1009 18069 1050 18092
rect 1410 17987 1444 17989
rect 1410 17955 1444 17987
rect 1410 17885 1444 17917
rect 1410 17883 1444 17885
rect 1568 17987 1602 17989
rect 1568 17955 1602 17987
rect 1568 17885 1602 17917
rect 1568 17883 1602 17885
rect 1698 17987 1732 17989
rect 1698 17955 1732 17987
rect 1698 17885 1732 17917
rect 1698 17883 1732 17885
rect 1856 17987 1890 17989
rect 1856 17955 1890 17987
rect 1856 17885 1890 17917
rect 1856 17883 1890 17885
rect 2030 17987 2064 17989
rect 2030 17955 2064 17987
rect 2030 17885 2064 17917
rect 2030 17883 2064 17885
rect 2188 17987 2222 17989
rect 2188 17955 2222 17987
rect 2188 17885 2222 17917
rect 2188 17883 2222 17885
rect 2372 17987 2406 17989
rect 2372 17955 2406 17987
rect 2372 17885 2406 17917
rect 2372 17883 2406 17885
rect 2530 17987 2564 17989
rect 2530 17955 2564 17987
rect 2776 17987 2810 17989
rect 2530 17885 2564 17917
rect 2530 17883 2564 17885
rect 2647 17903 2681 17937
rect 2776 17955 2810 17987
rect 2776 17885 2810 17917
rect 2776 17883 2810 17885
rect 2934 17987 2968 17989
rect 2934 17955 2968 17987
rect 2934 17885 2968 17917
rect 2934 17883 2968 17885
rect 1269 17749 1303 17783
rect 1773 17749 1807 17783
rect 2273 17747 2307 17781
rect 3797 18155 3807 18189
rect 3807 18155 3831 18189
rect 3869 18155 3875 18189
rect 3875 18155 3903 18189
rect 3941 18155 3943 18189
rect 3943 18155 3975 18189
rect 4013 18155 4045 18189
rect 4045 18155 4047 18189
rect 4085 18155 4113 18189
rect 4113 18155 4119 18189
rect 4157 18155 4181 18189
rect 4181 18155 4191 18189
rect 5756 18154 5766 18188
rect 5766 18154 5790 18188
rect 5828 18154 5834 18188
rect 5834 18154 5862 18188
rect 5900 18154 5902 18188
rect 5902 18154 5934 18188
rect 5972 18154 6004 18188
rect 6004 18154 6006 18188
rect 6044 18154 6072 18188
rect 6072 18154 6078 18188
rect 6116 18154 6140 18188
rect 6140 18154 6150 18188
rect 3120 17987 3154 17989
rect 3120 17955 3154 17987
rect 3120 17885 3154 17917
rect 3120 17883 3154 17885
rect 3278 17987 3312 17989
rect 3278 17955 3312 17987
rect 3278 17885 3312 17917
rect 3278 17883 3312 17885
rect 3742 17997 3776 17999
rect 3742 17965 3776 17997
rect 3742 17895 3776 17927
rect 3742 17893 3776 17895
rect 3900 17997 3934 17999
rect 3900 17965 3934 17997
rect 3900 17895 3934 17927
rect 3900 17893 3934 17895
rect 4050 17997 4084 17999
rect 4050 17965 4084 17997
rect 4050 17895 4084 17927
rect 4050 17893 4084 17895
rect 4208 17997 4242 17999
rect 4208 17965 4242 17997
rect 4208 17895 4242 17927
rect 4208 17893 4242 17895
rect 4402 17997 4436 17999
rect 4402 17965 4436 17997
rect 4402 17895 4436 17927
rect 4402 17893 4436 17895
rect 4560 17997 4594 17999
rect 4560 17965 4594 17997
rect 4560 17895 4594 17927
rect 4560 17893 4594 17895
rect 4710 17997 4744 17999
rect 4710 17965 4744 17997
rect 4710 17895 4744 17927
rect 4710 17893 4744 17895
rect 4868 17997 4902 17999
rect 4868 17965 4902 17997
rect 4868 17895 4902 17927
rect 4868 17893 4902 17895
rect 5700 17998 5734 18000
rect 5700 17966 5734 17998
rect 5700 17896 5734 17928
rect 5700 17894 5734 17896
rect 5858 17998 5892 18000
rect 5858 17966 5892 17998
rect 5858 17896 5892 17928
rect 5858 17894 5892 17896
rect 6008 17998 6042 18000
rect 6008 17966 6042 17998
rect 6008 17896 6042 17928
rect 6008 17894 6042 17896
rect 6166 17998 6200 18000
rect 6166 17966 6200 17998
rect 6166 17896 6200 17928
rect 6166 17894 6200 17896
rect 6360 17998 6394 18000
rect 6360 17966 6394 17998
rect 6360 17896 6394 17928
rect 6360 17894 6394 17896
rect 6518 17998 6552 18000
rect 6518 17966 6552 17998
rect 6518 17896 6552 17928
rect 6518 17894 6552 17896
rect 6668 17998 6702 18000
rect 6668 17966 6702 17998
rect 6668 17896 6702 17928
rect 6668 17894 6702 17896
rect 6826 17998 6860 18000
rect 6826 17966 6860 17998
rect 6826 17896 6860 17928
rect 6826 17894 6860 17896
rect 2857 17745 2891 17779
rect 3670 17769 3704 17803
rect 3984 17760 4018 17794
rect 1410 17631 1444 17665
rect 565 17552 606 17576
rect 712 17552 753 17576
rect 856 17558 897 17581
rect 1568 17631 1602 17665
rect 1698 17631 1732 17665
rect 1856 17631 1890 17665
rect 2030 17631 2064 17665
rect 2188 17631 2222 17665
rect 2372 17631 2406 17665
rect 1010 17558 1051 17582
rect 565 17536 569 17552
rect 569 17536 603 17552
rect 603 17536 606 17552
rect 712 17536 715 17552
rect 715 17536 749 17552
rect 749 17536 753 17552
rect 856 17541 859 17558
rect 859 17541 893 17558
rect 893 17541 897 17558
rect 1010 17542 1013 17558
rect 1013 17542 1047 17558
rect 1047 17542 1051 17558
rect 1373 17454 1387 17488
rect 1387 17454 1407 17488
rect 1445 17454 1455 17488
rect 1455 17454 1479 17488
rect 1517 17454 1523 17488
rect 1523 17454 1551 17488
rect 1589 17454 1591 17488
rect 1591 17454 1623 17488
rect 1661 17454 1693 17488
rect 1693 17454 1695 17488
rect 1733 17454 1761 17488
rect 1761 17454 1767 17488
rect 1805 17454 1829 17488
rect 1829 17454 1839 17488
rect 1877 17454 1897 17488
rect 1897 17454 1911 17488
rect 2530 17631 2564 17665
rect 2369 17429 2403 17463
rect 4306 17754 4340 17788
rect 4637 17772 4671 17806
rect 5628 17770 5662 17804
rect 5942 17760 5976 17794
rect 6264 17754 6298 17788
rect 6596 17772 6630 17806
rect 2776 17631 2810 17665
rect 2934 17631 2968 17665
rect 3120 17631 3154 17665
rect 3278 17631 3312 17665
rect 3742 17641 3776 17675
rect 3900 17641 3934 17675
rect 4050 17641 4084 17675
rect 4208 17641 4242 17675
rect 4402 17643 4436 17677
rect 4560 17643 4594 17677
rect 4710 17643 4744 17677
rect 4868 17643 4902 17677
rect 5700 17642 5734 17676
rect 5858 17642 5892 17676
rect 6008 17642 6042 17676
rect 6166 17642 6200 17676
rect 6360 17644 6394 17678
rect 6518 17644 6552 17678
rect 6668 17644 6702 17678
rect 6826 17644 6860 17678
rect 3741 17465 3753 17499
rect 3753 17465 3775 17499
rect 3813 17465 3821 17499
rect 3821 17465 3847 17499
rect 3885 17465 3889 17499
rect 3889 17465 3919 17499
rect 3957 17465 3991 17499
rect 4029 17465 4059 17499
rect 4059 17465 4063 17499
rect 4101 17465 4127 17499
rect 4127 17465 4135 17499
rect 4173 17465 4195 17499
rect 4195 17465 4207 17499
rect 5700 17466 5712 17500
rect 5712 17466 5734 17500
rect 5772 17466 5780 17500
rect 5780 17466 5806 17500
rect 5844 17466 5848 17500
rect 5848 17466 5878 17500
rect 5916 17466 5950 17500
rect 5988 17466 6018 17500
rect 6018 17466 6022 17500
rect 6060 17466 6086 17500
rect 6086 17466 6094 17500
rect 6132 17466 6154 17500
rect 6154 17466 6166 17500
rect 2642 17313 2696 17367
rect 1383 16928 1395 16962
rect 1395 16928 1417 16962
rect 1455 16928 1463 16962
rect 1463 16928 1489 16962
rect 1527 16928 1531 16962
rect 1531 16928 1561 16962
rect 1599 16928 1633 16962
rect 1671 16928 1701 16962
rect 1701 16928 1705 16962
rect 1743 16928 1769 16962
rect 1769 16928 1777 16962
rect 1815 16928 1837 16962
rect 1837 16928 1849 16962
rect 566 16858 569 16876
rect 569 16858 603 16876
rect 603 16858 607 16876
rect 710 16858 715 16876
rect 715 16858 749 16876
rect 749 16858 751 16876
rect 856 16864 859 16881
rect 859 16864 893 16881
rect 893 16864 897 16881
rect 1009 16864 1013 16881
rect 1013 16864 1047 16881
rect 1047 16864 1050 16881
rect 566 16836 607 16858
rect 710 16836 751 16858
rect 856 16841 897 16864
rect 1009 16841 1050 16864
rect 1410 16759 1444 16761
rect 1410 16727 1444 16759
rect 1410 16657 1444 16689
rect 1410 16655 1444 16657
rect 1568 16759 1602 16761
rect 1568 16727 1602 16759
rect 1568 16657 1602 16689
rect 1568 16655 1602 16657
rect 1698 16759 1732 16761
rect 1698 16727 1732 16759
rect 1698 16657 1732 16689
rect 1698 16655 1732 16657
rect 1856 16759 1890 16761
rect 1856 16727 1890 16759
rect 1856 16657 1890 16689
rect 1856 16655 1890 16657
rect 2030 16759 2064 16761
rect 2030 16727 2064 16759
rect 2030 16657 2064 16689
rect 2030 16655 2064 16657
rect 2188 16759 2222 16761
rect 2188 16727 2222 16759
rect 2188 16657 2222 16689
rect 2188 16655 2222 16657
rect 2372 16759 2406 16761
rect 2372 16727 2406 16759
rect 2372 16657 2406 16689
rect 2372 16655 2406 16657
rect 2530 16759 2564 16761
rect 2530 16727 2564 16759
rect 2776 16759 2810 16761
rect 2530 16657 2564 16689
rect 2530 16655 2564 16657
rect 2647 16675 2681 16709
rect 2776 16727 2810 16759
rect 2776 16657 2810 16689
rect 2776 16655 2810 16657
rect 2934 16759 2968 16761
rect 2934 16727 2968 16759
rect 2934 16657 2968 16689
rect 2934 16655 2968 16657
rect 1269 16521 1303 16555
rect 1773 16521 1807 16555
rect 2273 16519 2307 16553
rect 3797 16927 3807 16961
rect 3807 16927 3831 16961
rect 3869 16927 3875 16961
rect 3875 16927 3903 16961
rect 3941 16927 3943 16961
rect 3943 16927 3975 16961
rect 4013 16927 4045 16961
rect 4045 16927 4047 16961
rect 4085 16927 4113 16961
rect 4113 16927 4119 16961
rect 4157 16927 4181 16961
rect 4181 16927 4191 16961
rect 5756 16926 5766 16960
rect 5766 16926 5790 16960
rect 5828 16926 5834 16960
rect 5834 16926 5862 16960
rect 5900 16926 5902 16960
rect 5902 16926 5934 16960
rect 5972 16926 6004 16960
rect 6004 16926 6006 16960
rect 6044 16926 6072 16960
rect 6072 16926 6078 16960
rect 6116 16926 6140 16960
rect 6140 16926 6150 16960
rect 3120 16759 3154 16761
rect 3120 16727 3154 16759
rect 3120 16657 3154 16689
rect 3120 16655 3154 16657
rect 3278 16759 3312 16761
rect 3278 16727 3312 16759
rect 3278 16657 3312 16689
rect 3278 16655 3312 16657
rect 3742 16769 3776 16771
rect 3742 16737 3776 16769
rect 3742 16667 3776 16699
rect 3742 16665 3776 16667
rect 3900 16769 3934 16771
rect 3900 16737 3934 16769
rect 3900 16667 3934 16699
rect 3900 16665 3934 16667
rect 4050 16769 4084 16771
rect 4050 16737 4084 16769
rect 4050 16667 4084 16699
rect 4050 16665 4084 16667
rect 4208 16769 4242 16771
rect 4208 16737 4242 16769
rect 4208 16667 4242 16699
rect 4208 16665 4242 16667
rect 4402 16769 4436 16771
rect 4402 16737 4436 16769
rect 4402 16667 4436 16699
rect 4402 16665 4436 16667
rect 4560 16769 4594 16771
rect 4560 16737 4594 16769
rect 4560 16667 4594 16699
rect 4560 16665 4594 16667
rect 4710 16769 4744 16771
rect 4710 16737 4744 16769
rect 4710 16667 4744 16699
rect 4710 16665 4744 16667
rect 4868 16769 4902 16771
rect 4868 16737 4902 16769
rect 4868 16667 4902 16699
rect 4868 16665 4902 16667
rect 5700 16770 5734 16772
rect 5700 16738 5734 16770
rect 5700 16668 5734 16700
rect 5700 16666 5734 16668
rect 5858 16770 5892 16772
rect 5858 16738 5892 16770
rect 5858 16668 5892 16700
rect 5858 16666 5892 16668
rect 6008 16770 6042 16772
rect 6008 16738 6042 16770
rect 6008 16668 6042 16700
rect 6008 16666 6042 16668
rect 6166 16770 6200 16772
rect 6166 16738 6200 16770
rect 6166 16668 6200 16700
rect 6166 16666 6200 16668
rect 6360 16770 6394 16772
rect 6360 16738 6394 16770
rect 6360 16668 6394 16700
rect 6360 16666 6394 16668
rect 6518 16770 6552 16772
rect 6518 16738 6552 16770
rect 6518 16668 6552 16700
rect 6518 16666 6552 16668
rect 6668 16770 6702 16772
rect 6668 16738 6702 16770
rect 6668 16668 6702 16700
rect 6668 16666 6702 16668
rect 6826 16770 6860 16772
rect 6826 16738 6860 16770
rect 6826 16668 6860 16700
rect 6826 16666 6860 16668
rect 2857 16517 2891 16551
rect 3670 16541 3704 16575
rect 3984 16532 4018 16566
rect 1410 16403 1444 16437
rect 565 16324 606 16348
rect 712 16324 753 16348
rect 856 16330 897 16353
rect 1568 16403 1602 16437
rect 1698 16403 1732 16437
rect 1856 16403 1890 16437
rect 2030 16403 2064 16437
rect 2188 16403 2222 16437
rect 2372 16403 2406 16437
rect 1010 16330 1051 16354
rect 565 16308 569 16324
rect 569 16308 603 16324
rect 603 16308 606 16324
rect 712 16308 715 16324
rect 715 16308 749 16324
rect 749 16308 753 16324
rect 856 16313 859 16330
rect 859 16313 893 16330
rect 893 16313 897 16330
rect 1010 16314 1013 16330
rect 1013 16314 1047 16330
rect 1047 16314 1051 16330
rect 1373 16226 1387 16260
rect 1387 16226 1407 16260
rect 1445 16226 1455 16260
rect 1455 16226 1479 16260
rect 1517 16226 1523 16260
rect 1523 16226 1551 16260
rect 1589 16226 1591 16260
rect 1591 16226 1623 16260
rect 1661 16226 1693 16260
rect 1693 16226 1695 16260
rect 1733 16226 1761 16260
rect 1761 16226 1767 16260
rect 1805 16226 1829 16260
rect 1829 16226 1839 16260
rect 1877 16226 1897 16260
rect 1897 16226 1911 16260
rect 2530 16403 2564 16437
rect 2369 16201 2403 16235
rect 4306 16526 4340 16560
rect 4637 16544 4671 16578
rect 5628 16542 5662 16576
rect 5942 16532 5976 16566
rect 6264 16526 6298 16560
rect 6596 16544 6630 16578
rect 2776 16403 2810 16437
rect 2934 16403 2968 16437
rect 3120 16403 3154 16437
rect 3278 16403 3312 16437
rect 3742 16413 3776 16447
rect 3900 16413 3934 16447
rect 4050 16413 4084 16447
rect 4208 16413 4242 16447
rect 4402 16415 4436 16449
rect 4560 16415 4594 16449
rect 4710 16415 4744 16449
rect 4868 16415 4902 16449
rect 5700 16414 5734 16448
rect 5858 16414 5892 16448
rect 6008 16414 6042 16448
rect 6166 16414 6200 16448
rect 6360 16416 6394 16450
rect 6518 16416 6552 16450
rect 6668 16416 6702 16450
rect 6826 16416 6860 16450
rect 3741 16237 3753 16271
rect 3753 16237 3775 16271
rect 3813 16237 3821 16271
rect 3821 16237 3847 16271
rect 3885 16237 3889 16271
rect 3889 16237 3919 16271
rect 3957 16237 3991 16271
rect 4029 16237 4059 16271
rect 4059 16237 4063 16271
rect 4101 16237 4127 16271
rect 4127 16237 4135 16271
rect 4173 16237 4195 16271
rect 4195 16237 4207 16271
rect 5700 16238 5712 16272
rect 5712 16238 5734 16272
rect 5772 16238 5780 16272
rect 5780 16238 5806 16272
rect 5844 16238 5848 16272
rect 5848 16238 5878 16272
rect 5916 16238 5950 16272
rect 5988 16238 6018 16272
rect 6018 16238 6022 16272
rect 6060 16238 6086 16272
rect 6086 16238 6094 16272
rect 6132 16238 6154 16272
rect 6154 16238 6166 16272
rect 2642 16085 2696 16139
rect 1383 15700 1395 15734
rect 1395 15700 1417 15734
rect 1455 15700 1463 15734
rect 1463 15700 1489 15734
rect 1527 15700 1531 15734
rect 1531 15700 1561 15734
rect 1599 15700 1633 15734
rect 1671 15700 1701 15734
rect 1701 15700 1705 15734
rect 1743 15700 1769 15734
rect 1769 15700 1777 15734
rect 1815 15700 1837 15734
rect 1837 15700 1849 15734
rect 566 15630 569 15648
rect 569 15630 603 15648
rect 603 15630 607 15648
rect 710 15630 715 15648
rect 715 15630 749 15648
rect 749 15630 751 15648
rect 856 15636 859 15653
rect 859 15636 893 15653
rect 893 15636 897 15653
rect 1009 15636 1013 15653
rect 1013 15636 1047 15653
rect 1047 15636 1050 15653
rect 566 15608 607 15630
rect 710 15608 751 15630
rect 856 15613 897 15636
rect 1009 15613 1050 15636
rect 1410 15531 1444 15533
rect 1410 15499 1444 15531
rect 1410 15429 1444 15461
rect 1410 15427 1444 15429
rect 1568 15531 1602 15533
rect 1568 15499 1602 15531
rect 1568 15429 1602 15461
rect 1568 15427 1602 15429
rect 1698 15531 1732 15533
rect 1698 15499 1732 15531
rect 1698 15429 1732 15461
rect 1698 15427 1732 15429
rect 1856 15531 1890 15533
rect 1856 15499 1890 15531
rect 1856 15429 1890 15461
rect 1856 15427 1890 15429
rect 2030 15531 2064 15533
rect 2030 15499 2064 15531
rect 2030 15429 2064 15461
rect 2030 15427 2064 15429
rect 2188 15531 2222 15533
rect 2188 15499 2222 15531
rect 2188 15429 2222 15461
rect 2188 15427 2222 15429
rect 2372 15531 2406 15533
rect 2372 15499 2406 15531
rect 2372 15429 2406 15461
rect 2372 15427 2406 15429
rect 2530 15531 2564 15533
rect 2530 15499 2564 15531
rect 2776 15531 2810 15533
rect 2530 15429 2564 15461
rect 2530 15427 2564 15429
rect 2647 15447 2681 15481
rect 2776 15499 2810 15531
rect 2776 15429 2810 15461
rect 2776 15427 2810 15429
rect 2934 15531 2968 15533
rect 2934 15499 2968 15531
rect 2934 15429 2968 15461
rect 2934 15427 2968 15429
rect 1269 15293 1303 15327
rect 1773 15293 1807 15327
rect 2273 15291 2307 15325
rect 3797 15699 3807 15733
rect 3807 15699 3831 15733
rect 3869 15699 3875 15733
rect 3875 15699 3903 15733
rect 3941 15699 3943 15733
rect 3943 15699 3975 15733
rect 4013 15699 4045 15733
rect 4045 15699 4047 15733
rect 4085 15699 4113 15733
rect 4113 15699 4119 15733
rect 4157 15699 4181 15733
rect 4181 15699 4191 15733
rect 5756 15698 5766 15732
rect 5766 15698 5790 15732
rect 5828 15698 5834 15732
rect 5834 15698 5862 15732
rect 5900 15698 5902 15732
rect 5902 15698 5934 15732
rect 5972 15698 6004 15732
rect 6004 15698 6006 15732
rect 6044 15698 6072 15732
rect 6072 15698 6078 15732
rect 6116 15698 6140 15732
rect 6140 15698 6150 15732
rect 3120 15531 3154 15533
rect 3120 15499 3154 15531
rect 3120 15429 3154 15461
rect 3120 15427 3154 15429
rect 3278 15531 3312 15533
rect 3278 15499 3312 15531
rect 3278 15429 3312 15461
rect 3278 15427 3312 15429
rect 3742 15541 3776 15543
rect 3742 15509 3776 15541
rect 3742 15439 3776 15471
rect 3742 15437 3776 15439
rect 3900 15541 3934 15543
rect 3900 15509 3934 15541
rect 3900 15439 3934 15471
rect 3900 15437 3934 15439
rect 4050 15541 4084 15543
rect 4050 15509 4084 15541
rect 4050 15439 4084 15471
rect 4050 15437 4084 15439
rect 4208 15541 4242 15543
rect 4208 15509 4242 15541
rect 4208 15439 4242 15471
rect 4208 15437 4242 15439
rect 4402 15541 4436 15543
rect 4402 15509 4436 15541
rect 4402 15439 4436 15471
rect 4402 15437 4436 15439
rect 4560 15541 4594 15543
rect 4560 15509 4594 15541
rect 4560 15439 4594 15471
rect 4560 15437 4594 15439
rect 4710 15541 4744 15543
rect 4710 15509 4744 15541
rect 4710 15439 4744 15471
rect 4710 15437 4744 15439
rect 4868 15541 4902 15543
rect 4868 15509 4902 15541
rect 4868 15439 4902 15471
rect 4868 15437 4902 15439
rect 5700 15542 5734 15544
rect 5700 15510 5734 15542
rect 5700 15440 5734 15472
rect 5700 15438 5734 15440
rect 5858 15542 5892 15544
rect 5858 15510 5892 15542
rect 5858 15440 5892 15472
rect 5858 15438 5892 15440
rect 6008 15542 6042 15544
rect 6008 15510 6042 15542
rect 6008 15440 6042 15472
rect 6008 15438 6042 15440
rect 6166 15542 6200 15544
rect 6166 15510 6200 15542
rect 6166 15440 6200 15472
rect 6166 15438 6200 15440
rect 6360 15542 6394 15544
rect 6360 15510 6394 15542
rect 6360 15440 6394 15472
rect 6360 15438 6394 15440
rect 6518 15542 6552 15544
rect 6518 15510 6552 15542
rect 6518 15440 6552 15472
rect 6518 15438 6552 15440
rect 6668 15542 6702 15544
rect 6668 15510 6702 15542
rect 6668 15440 6702 15472
rect 6668 15438 6702 15440
rect 6826 15542 6860 15544
rect 6826 15510 6860 15542
rect 6826 15440 6860 15472
rect 6826 15438 6860 15440
rect 2857 15289 2891 15323
rect 3670 15313 3704 15347
rect 3984 15304 4018 15338
rect 1410 15175 1444 15209
rect 565 15096 606 15120
rect 712 15096 753 15120
rect 856 15102 897 15125
rect 1568 15175 1602 15209
rect 1698 15175 1732 15209
rect 1856 15175 1890 15209
rect 2030 15175 2064 15209
rect 2188 15175 2222 15209
rect 2372 15175 2406 15209
rect 1010 15102 1051 15126
rect 565 15080 569 15096
rect 569 15080 603 15096
rect 603 15080 606 15096
rect 712 15080 715 15096
rect 715 15080 749 15096
rect 749 15080 753 15096
rect 856 15085 859 15102
rect 859 15085 893 15102
rect 893 15085 897 15102
rect 1010 15086 1013 15102
rect 1013 15086 1047 15102
rect 1047 15086 1051 15102
rect 1373 14998 1387 15032
rect 1387 14998 1407 15032
rect 1445 14998 1455 15032
rect 1455 14998 1479 15032
rect 1517 14998 1523 15032
rect 1523 14998 1551 15032
rect 1589 14998 1591 15032
rect 1591 14998 1623 15032
rect 1661 14998 1693 15032
rect 1693 14998 1695 15032
rect 1733 14998 1761 15032
rect 1761 14998 1767 15032
rect 1805 14998 1829 15032
rect 1829 14998 1839 15032
rect 1877 14998 1897 15032
rect 1897 14998 1911 15032
rect 2530 15175 2564 15209
rect 2369 14973 2403 15007
rect 4306 15298 4340 15332
rect 4637 15316 4671 15350
rect 5628 15314 5662 15348
rect 5942 15304 5976 15338
rect 6264 15298 6298 15332
rect 6596 15316 6630 15350
rect 2776 15175 2810 15209
rect 2934 15175 2968 15209
rect 3120 15175 3154 15209
rect 3278 15175 3312 15209
rect 3742 15185 3776 15219
rect 3900 15185 3934 15219
rect 4050 15185 4084 15219
rect 4208 15185 4242 15219
rect 4402 15187 4436 15221
rect 4560 15187 4594 15221
rect 4710 15187 4744 15221
rect 4868 15187 4902 15221
rect 5700 15186 5734 15220
rect 5858 15186 5892 15220
rect 6008 15186 6042 15220
rect 6166 15186 6200 15220
rect 6360 15188 6394 15222
rect 6518 15188 6552 15222
rect 6668 15188 6702 15222
rect 6826 15188 6860 15222
rect 3741 15009 3753 15043
rect 3753 15009 3775 15043
rect 3813 15009 3821 15043
rect 3821 15009 3847 15043
rect 3885 15009 3889 15043
rect 3889 15009 3919 15043
rect 3957 15009 3991 15043
rect 4029 15009 4059 15043
rect 4059 15009 4063 15043
rect 4101 15009 4127 15043
rect 4127 15009 4135 15043
rect 4173 15009 4195 15043
rect 4195 15009 4207 15043
rect 5700 15010 5712 15044
rect 5712 15010 5734 15044
rect 5772 15010 5780 15044
rect 5780 15010 5806 15044
rect 5844 15010 5848 15044
rect 5848 15010 5878 15044
rect 5916 15010 5950 15044
rect 5988 15010 6018 15044
rect 6018 15010 6022 15044
rect 6060 15010 6086 15044
rect 6086 15010 6094 15044
rect 6132 15010 6154 15044
rect 6154 15010 6166 15044
rect 2642 14857 2696 14911
rect 1383 14472 1395 14506
rect 1395 14472 1417 14506
rect 1455 14472 1463 14506
rect 1463 14472 1489 14506
rect 1527 14472 1531 14506
rect 1531 14472 1561 14506
rect 1599 14472 1633 14506
rect 1671 14472 1701 14506
rect 1701 14472 1705 14506
rect 1743 14472 1769 14506
rect 1769 14472 1777 14506
rect 1815 14472 1837 14506
rect 1837 14472 1849 14506
rect 566 14402 569 14420
rect 569 14402 603 14420
rect 603 14402 607 14420
rect 710 14402 715 14420
rect 715 14402 749 14420
rect 749 14402 751 14420
rect 856 14408 859 14425
rect 859 14408 893 14425
rect 893 14408 897 14425
rect 1009 14408 1013 14425
rect 1013 14408 1047 14425
rect 1047 14408 1050 14425
rect 566 14380 607 14402
rect 710 14380 751 14402
rect 856 14385 897 14408
rect 1009 14385 1050 14408
rect 1410 14303 1444 14305
rect 1410 14271 1444 14303
rect 1410 14201 1444 14233
rect 1410 14199 1444 14201
rect 1568 14303 1602 14305
rect 1568 14271 1602 14303
rect 1568 14201 1602 14233
rect 1568 14199 1602 14201
rect 1698 14303 1732 14305
rect 1698 14271 1732 14303
rect 1698 14201 1732 14233
rect 1698 14199 1732 14201
rect 1856 14303 1890 14305
rect 1856 14271 1890 14303
rect 1856 14201 1890 14233
rect 1856 14199 1890 14201
rect 2030 14303 2064 14305
rect 2030 14271 2064 14303
rect 2030 14201 2064 14233
rect 2030 14199 2064 14201
rect 2188 14303 2222 14305
rect 2188 14271 2222 14303
rect 2188 14201 2222 14233
rect 2188 14199 2222 14201
rect 2372 14303 2406 14305
rect 2372 14271 2406 14303
rect 2372 14201 2406 14233
rect 2372 14199 2406 14201
rect 2530 14303 2564 14305
rect 2530 14271 2564 14303
rect 2776 14303 2810 14305
rect 2530 14201 2564 14233
rect 2530 14199 2564 14201
rect 2647 14219 2681 14253
rect 2776 14271 2810 14303
rect 2776 14201 2810 14233
rect 2776 14199 2810 14201
rect 2934 14303 2968 14305
rect 2934 14271 2968 14303
rect 2934 14201 2968 14233
rect 2934 14199 2968 14201
rect 1269 14065 1303 14099
rect 1773 14065 1807 14099
rect 2273 14063 2307 14097
rect 3797 14471 3807 14505
rect 3807 14471 3831 14505
rect 3869 14471 3875 14505
rect 3875 14471 3903 14505
rect 3941 14471 3943 14505
rect 3943 14471 3975 14505
rect 4013 14471 4045 14505
rect 4045 14471 4047 14505
rect 4085 14471 4113 14505
rect 4113 14471 4119 14505
rect 4157 14471 4181 14505
rect 4181 14471 4191 14505
rect 5756 14470 5766 14504
rect 5766 14470 5790 14504
rect 5828 14470 5834 14504
rect 5834 14470 5862 14504
rect 5900 14470 5902 14504
rect 5902 14470 5934 14504
rect 5972 14470 6004 14504
rect 6004 14470 6006 14504
rect 6044 14470 6072 14504
rect 6072 14470 6078 14504
rect 6116 14470 6140 14504
rect 6140 14470 6150 14504
rect 3120 14303 3154 14305
rect 3120 14271 3154 14303
rect 3120 14201 3154 14233
rect 3120 14199 3154 14201
rect 3278 14303 3312 14305
rect 3278 14271 3312 14303
rect 3278 14201 3312 14233
rect 3278 14199 3312 14201
rect 3742 14313 3776 14315
rect 3742 14281 3776 14313
rect 3742 14211 3776 14243
rect 3742 14209 3776 14211
rect 3900 14313 3934 14315
rect 3900 14281 3934 14313
rect 3900 14211 3934 14243
rect 3900 14209 3934 14211
rect 4050 14313 4084 14315
rect 4050 14281 4084 14313
rect 4050 14211 4084 14243
rect 4050 14209 4084 14211
rect 4208 14313 4242 14315
rect 4208 14281 4242 14313
rect 4208 14211 4242 14243
rect 4208 14209 4242 14211
rect 4402 14313 4436 14315
rect 4402 14281 4436 14313
rect 4402 14211 4436 14243
rect 4402 14209 4436 14211
rect 4560 14313 4594 14315
rect 4560 14281 4594 14313
rect 4560 14211 4594 14243
rect 4560 14209 4594 14211
rect 4710 14313 4744 14315
rect 4710 14281 4744 14313
rect 4710 14211 4744 14243
rect 4710 14209 4744 14211
rect 4868 14313 4902 14315
rect 4868 14281 4902 14313
rect 4868 14211 4902 14243
rect 4868 14209 4902 14211
rect 5700 14314 5734 14316
rect 5700 14282 5734 14314
rect 5700 14212 5734 14244
rect 5700 14210 5734 14212
rect 5858 14314 5892 14316
rect 5858 14282 5892 14314
rect 5858 14212 5892 14244
rect 5858 14210 5892 14212
rect 6008 14314 6042 14316
rect 6008 14282 6042 14314
rect 6008 14212 6042 14244
rect 6008 14210 6042 14212
rect 6166 14314 6200 14316
rect 6166 14282 6200 14314
rect 6166 14212 6200 14244
rect 6166 14210 6200 14212
rect 6360 14314 6394 14316
rect 6360 14282 6394 14314
rect 6360 14212 6394 14244
rect 6360 14210 6394 14212
rect 6518 14314 6552 14316
rect 6518 14282 6552 14314
rect 6518 14212 6552 14244
rect 6518 14210 6552 14212
rect 6668 14314 6702 14316
rect 6668 14282 6702 14314
rect 6668 14212 6702 14244
rect 6668 14210 6702 14212
rect 6826 14314 6860 14316
rect 6826 14282 6860 14314
rect 6826 14212 6860 14244
rect 6826 14210 6860 14212
rect 2857 14061 2891 14095
rect 3670 14085 3704 14119
rect 3984 14076 4018 14110
rect 1410 13947 1444 13981
rect 565 13868 606 13892
rect 712 13868 753 13892
rect 856 13874 897 13897
rect 1568 13947 1602 13981
rect 1698 13947 1732 13981
rect 1856 13947 1890 13981
rect 2030 13947 2064 13981
rect 2188 13947 2222 13981
rect 2372 13947 2406 13981
rect 1010 13874 1051 13898
rect 565 13852 569 13868
rect 569 13852 603 13868
rect 603 13852 606 13868
rect 712 13852 715 13868
rect 715 13852 749 13868
rect 749 13852 753 13868
rect 856 13857 859 13874
rect 859 13857 893 13874
rect 893 13857 897 13874
rect 1010 13858 1013 13874
rect 1013 13858 1047 13874
rect 1047 13858 1051 13874
rect 1373 13770 1387 13804
rect 1387 13770 1407 13804
rect 1445 13770 1455 13804
rect 1455 13770 1479 13804
rect 1517 13770 1523 13804
rect 1523 13770 1551 13804
rect 1589 13770 1591 13804
rect 1591 13770 1623 13804
rect 1661 13770 1693 13804
rect 1693 13770 1695 13804
rect 1733 13770 1761 13804
rect 1761 13770 1767 13804
rect 1805 13770 1829 13804
rect 1829 13770 1839 13804
rect 1877 13770 1897 13804
rect 1897 13770 1911 13804
rect 2530 13947 2564 13981
rect 2369 13745 2403 13779
rect 4306 14070 4340 14104
rect 4637 14088 4671 14122
rect 5628 14086 5662 14120
rect 5942 14076 5976 14110
rect 6264 14070 6298 14104
rect 6596 14088 6630 14122
rect 2776 13947 2810 13981
rect 2934 13947 2968 13981
rect 3120 13947 3154 13981
rect 3278 13947 3312 13981
rect 3742 13957 3776 13991
rect 3900 13957 3934 13991
rect 4050 13957 4084 13991
rect 4208 13957 4242 13991
rect 4402 13959 4436 13993
rect 4560 13959 4594 13993
rect 4710 13959 4744 13993
rect 4868 13959 4902 13993
rect 5700 13958 5734 13992
rect 5858 13958 5892 13992
rect 6008 13958 6042 13992
rect 6166 13958 6200 13992
rect 6360 13960 6394 13994
rect 6518 13960 6552 13994
rect 6668 13960 6702 13994
rect 6826 13960 6860 13994
rect 3741 13781 3753 13815
rect 3753 13781 3775 13815
rect 3813 13781 3821 13815
rect 3821 13781 3847 13815
rect 3885 13781 3889 13815
rect 3889 13781 3919 13815
rect 3957 13781 3991 13815
rect 4029 13781 4059 13815
rect 4059 13781 4063 13815
rect 4101 13781 4127 13815
rect 4127 13781 4135 13815
rect 4173 13781 4195 13815
rect 4195 13781 4207 13815
rect 5700 13782 5712 13816
rect 5712 13782 5734 13816
rect 5772 13782 5780 13816
rect 5780 13782 5806 13816
rect 5844 13782 5848 13816
rect 5848 13782 5878 13816
rect 5916 13782 5950 13816
rect 5988 13782 6018 13816
rect 6018 13782 6022 13816
rect 6060 13782 6086 13816
rect 6086 13782 6094 13816
rect 6132 13782 6154 13816
rect 6154 13782 6166 13816
rect 2642 13629 2696 13683
rect 1383 13244 1395 13278
rect 1395 13244 1417 13278
rect 1455 13244 1463 13278
rect 1463 13244 1489 13278
rect 1527 13244 1531 13278
rect 1531 13244 1561 13278
rect 1599 13244 1633 13278
rect 1671 13244 1701 13278
rect 1701 13244 1705 13278
rect 1743 13244 1769 13278
rect 1769 13244 1777 13278
rect 1815 13244 1837 13278
rect 1837 13244 1849 13278
rect 566 13174 569 13192
rect 569 13174 603 13192
rect 603 13174 607 13192
rect 710 13174 715 13192
rect 715 13174 749 13192
rect 749 13174 751 13192
rect 856 13180 859 13197
rect 859 13180 893 13197
rect 893 13180 897 13197
rect 1009 13180 1013 13197
rect 1013 13180 1047 13197
rect 1047 13180 1050 13197
rect 566 13152 607 13174
rect 710 13152 751 13174
rect 856 13157 897 13180
rect 1009 13157 1050 13180
rect 1410 13075 1444 13077
rect 1410 13043 1444 13075
rect 1410 12973 1444 13005
rect 1410 12971 1444 12973
rect 1568 13075 1602 13077
rect 1568 13043 1602 13075
rect 1568 12973 1602 13005
rect 1568 12971 1602 12973
rect 1698 13075 1732 13077
rect 1698 13043 1732 13075
rect 1698 12973 1732 13005
rect 1698 12971 1732 12973
rect 1856 13075 1890 13077
rect 1856 13043 1890 13075
rect 1856 12973 1890 13005
rect 1856 12971 1890 12973
rect 2030 13075 2064 13077
rect 2030 13043 2064 13075
rect 2030 12973 2064 13005
rect 2030 12971 2064 12973
rect 2188 13075 2222 13077
rect 2188 13043 2222 13075
rect 2188 12973 2222 13005
rect 2188 12971 2222 12973
rect 2372 13075 2406 13077
rect 2372 13043 2406 13075
rect 2372 12973 2406 13005
rect 2372 12971 2406 12973
rect 2530 13075 2564 13077
rect 2530 13043 2564 13075
rect 2776 13075 2810 13077
rect 2530 12973 2564 13005
rect 2530 12971 2564 12973
rect 2647 12991 2681 13025
rect 2776 13043 2810 13075
rect 2776 12973 2810 13005
rect 2776 12971 2810 12973
rect 2934 13075 2968 13077
rect 2934 13043 2968 13075
rect 2934 12973 2968 13005
rect 2934 12971 2968 12973
rect 1269 12837 1303 12871
rect 1773 12837 1807 12871
rect 2273 12835 2307 12869
rect 3797 13243 3807 13277
rect 3807 13243 3831 13277
rect 3869 13243 3875 13277
rect 3875 13243 3903 13277
rect 3941 13243 3943 13277
rect 3943 13243 3975 13277
rect 4013 13243 4045 13277
rect 4045 13243 4047 13277
rect 4085 13243 4113 13277
rect 4113 13243 4119 13277
rect 4157 13243 4181 13277
rect 4181 13243 4191 13277
rect 5756 13242 5766 13276
rect 5766 13242 5790 13276
rect 5828 13242 5834 13276
rect 5834 13242 5862 13276
rect 5900 13242 5902 13276
rect 5902 13242 5934 13276
rect 5972 13242 6004 13276
rect 6004 13242 6006 13276
rect 6044 13242 6072 13276
rect 6072 13242 6078 13276
rect 6116 13242 6140 13276
rect 6140 13242 6150 13276
rect 3120 13075 3154 13077
rect 3120 13043 3154 13075
rect 3120 12973 3154 13005
rect 3120 12971 3154 12973
rect 3278 13075 3312 13077
rect 3278 13043 3312 13075
rect 3278 12973 3312 13005
rect 3278 12971 3312 12973
rect 3742 13085 3776 13087
rect 3742 13053 3776 13085
rect 3742 12983 3776 13015
rect 3742 12981 3776 12983
rect 3900 13085 3934 13087
rect 3900 13053 3934 13085
rect 3900 12983 3934 13015
rect 3900 12981 3934 12983
rect 4050 13085 4084 13087
rect 4050 13053 4084 13085
rect 4050 12983 4084 13015
rect 4050 12981 4084 12983
rect 4208 13085 4242 13087
rect 4208 13053 4242 13085
rect 4208 12983 4242 13015
rect 4208 12981 4242 12983
rect 4402 13085 4436 13087
rect 4402 13053 4436 13085
rect 4402 12983 4436 13015
rect 4402 12981 4436 12983
rect 4560 13085 4594 13087
rect 4560 13053 4594 13085
rect 4560 12983 4594 13015
rect 4560 12981 4594 12983
rect 4710 13085 4744 13087
rect 4710 13053 4744 13085
rect 4710 12983 4744 13015
rect 4710 12981 4744 12983
rect 4868 13085 4902 13087
rect 4868 13053 4902 13085
rect 4868 12983 4902 13015
rect 4868 12981 4902 12983
rect 5700 13086 5734 13088
rect 5700 13054 5734 13086
rect 5700 12984 5734 13016
rect 5700 12982 5734 12984
rect 5858 13086 5892 13088
rect 5858 13054 5892 13086
rect 5858 12984 5892 13016
rect 5858 12982 5892 12984
rect 6008 13086 6042 13088
rect 6008 13054 6042 13086
rect 6008 12984 6042 13016
rect 6008 12982 6042 12984
rect 6166 13086 6200 13088
rect 6166 13054 6200 13086
rect 6166 12984 6200 13016
rect 6166 12982 6200 12984
rect 6360 13086 6394 13088
rect 6360 13054 6394 13086
rect 6360 12984 6394 13016
rect 6360 12982 6394 12984
rect 6518 13086 6552 13088
rect 6518 13054 6552 13086
rect 6518 12984 6552 13016
rect 6518 12982 6552 12984
rect 6668 13086 6702 13088
rect 6668 13054 6702 13086
rect 6668 12984 6702 13016
rect 6668 12982 6702 12984
rect 6826 13086 6860 13088
rect 6826 13054 6860 13086
rect 6826 12984 6860 13016
rect 6826 12982 6860 12984
rect 2857 12833 2891 12867
rect 3670 12857 3704 12891
rect 3984 12848 4018 12882
rect 1410 12719 1444 12753
rect 565 12640 606 12664
rect 712 12640 753 12664
rect 856 12646 897 12669
rect 1568 12719 1602 12753
rect 1698 12719 1732 12753
rect 1856 12719 1890 12753
rect 2030 12719 2064 12753
rect 2188 12719 2222 12753
rect 2372 12719 2406 12753
rect 1010 12646 1051 12670
rect 565 12624 569 12640
rect 569 12624 603 12640
rect 603 12624 606 12640
rect 712 12624 715 12640
rect 715 12624 749 12640
rect 749 12624 753 12640
rect 856 12629 859 12646
rect 859 12629 893 12646
rect 893 12629 897 12646
rect 1010 12630 1013 12646
rect 1013 12630 1047 12646
rect 1047 12630 1051 12646
rect 1373 12542 1387 12576
rect 1387 12542 1407 12576
rect 1445 12542 1455 12576
rect 1455 12542 1479 12576
rect 1517 12542 1523 12576
rect 1523 12542 1551 12576
rect 1589 12542 1591 12576
rect 1591 12542 1623 12576
rect 1661 12542 1693 12576
rect 1693 12542 1695 12576
rect 1733 12542 1761 12576
rect 1761 12542 1767 12576
rect 1805 12542 1829 12576
rect 1829 12542 1839 12576
rect 1877 12542 1897 12576
rect 1897 12542 1911 12576
rect 2530 12719 2564 12753
rect 2369 12517 2403 12551
rect 4306 12842 4340 12876
rect 4637 12860 4671 12894
rect 5628 12858 5662 12892
rect 5942 12848 5976 12882
rect 6264 12842 6298 12876
rect 6596 12860 6630 12894
rect 2776 12719 2810 12753
rect 2934 12719 2968 12753
rect 3120 12719 3154 12753
rect 3278 12719 3312 12753
rect 3742 12729 3776 12763
rect 3900 12729 3934 12763
rect 4050 12729 4084 12763
rect 4208 12729 4242 12763
rect 4402 12731 4436 12765
rect 4560 12731 4594 12765
rect 4710 12731 4744 12765
rect 4868 12731 4902 12765
rect 5700 12730 5734 12764
rect 5858 12730 5892 12764
rect 6008 12730 6042 12764
rect 6166 12730 6200 12764
rect 6360 12732 6394 12766
rect 6518 12732 6552 12766
rect 6668 12732 6702 12766
rect 6826 12732 6860 12766
rect 3741 12553 3753 12587
rect 3753 12553 3775 12587
rect 3813 12553 3821 12587
rect 3821 12553 3847 12587
rect 3885 12553 3889 12587
rect 3889 12553 3919 12587
rect 3957 12553 3991 12587
rect 4029 12553 4059 12587
rect 4059 12553 4063 12587
rect 4101 12553 4127 12587
rect 4127 12553 4135 12587
rect 4173 12553 4195 12587
rect 4195 12553 4207 12587
rect 5700 12554 5712 12588
rect 5712 12554 5734 12588
rect 5772 12554 5780 12588
rect 5780 12554 5806 12588
rect 5844 12554 5848 12588
rect 5848 12554 5878 12588
rect 5916 12554 5950 12588
rect 5988 12554 6018 12588
rect 6018 12554 6022 12588
rect 6060 12554 6086 12588
rect 6086 12554 6094 12588
rect 6132 12554 6154 12588
rect 6154 12554 6166 12588
rect 2642 12401 2696 12455
rect 1383 12016 1395 12050
rect 1395 12016 1417 12050
rect 1455 12016 1463 12050
rect 1463 12016 1489 12050
rect 1527 12016 1531 12050
rect 1531 12016 1561 12050
rect 1599 12016 1633 12050
rect 1671 12016 1701 12050
rect 1701 12016 1705 12050
rect 1743 12016 1769 12050
rect 1769 12016 1777 12050
rect 1815 12016 1837 12050
rect 1837 12016 1849 12050
rect 566 11946 569 11964
rect 569 11946 603 11964
rect 603 11946 607 11964
rect 710 11946 715 11964
rect 715 11946 749 11964
rect 749 11946 751 11964
rect 856 11952 859 11969
rect 859 11952 893 11969
rect 893 11952 897 11969
rect 1009 11952 1013 11969
rect 1013 11952 1047 11969
rect 1047 11952 1050 11969
rect 566 11924 607 11946
rect 710 11924 751 11946
rect 856 11929 897 11952
rect 1009 11929 1050 11952
rect 1410 11847 1444 11849
rect 1410 11815 1444 11847
rect 1410 11745 1444 11777
rect 1410 11743 1444 11745
rect 1568 11847 1602 11849
rect 1568 11815 1602 11847
rect 1568 11745 1602 11777
rect 1568 11743 1602 11745
rect 1698 11847 1732 11849
rect 1698 11815 1732 11847
rect 1698 11745 1732 11777
rect 1698 11743 1732 11745
rect 1856 11847 1890 11849
rect 1856 11815 1890 11847
rect 1856 11745 1890 11777
rect 1856 11743 1890 11745
rect 2030 11847 2064 11849
rect 2030 11815 2064 11847
rect 2030 11745 2064 11777
rect 2030 11743 2064 11745
rect 2188 11847 2222 11849
rect 2188 11815 2222 11847
rect 2188 11745 2222 11777
rect 2188 11743 2222 11745
rect 2372 11847 2406 11849
rect 2372 11815 2406 11847
rect 2372 11745 2406 11777
rect 2372 11743 2406 11745
rect 2530 11847 2564 11849
rect 2530 11815 2564 11847
rect 2776 11847 2810 11849
rect 2530 11745 2564 11777
rect 2530 11743 2564 11745
rect 2647 11763 2681 11797
rect 2776 11815 2810 11847
rect 2776 11745 2810 11777
rect 2776 11743 2810 11745
rect 2934 11847 2968 11849
rect 2934 11815 2968 11847
rect 2934 11745 2968 11777
rect 2934 11743 2968 11745
rect 1269 11609 1303 11643
rect 1773 11609 1807 11643
rect 2273 11607 2307 11641
rect 3797 12015 3807 12049
rect 3807 12015 3831 12049
rect 3869 12015 3875 12049
rect 3875 12015 3903 12049
rect 3941 12015 3943 12049
rect 3943 12015 3975 12049
rect 4013 12015 4045 12049
rect 4045 12015 4047 12049
rect 4085 12015 4113 12049
rect 4113 12015 4119 12049
rect 4157 12015 4181 12049
rect 4181 12015 4191 12049
rect 5756 12014 5766 12048
rect 5766 12014 5790 12048
rect 5828 12014 5834 12048
rect 5834 12014 5862 12048
rect 5900 12014 5902 12048
rect 5902 12014 5934 12048
rect 5972 12014 6004 12048
rect 6004 12014 6006 12048
rect 6044 12014 6072 12048
rect 6072 12014 6078 12048
rect 6116 12014 6140 12048
rect 6140 12014 6150 12048
rect 3120 11847 3154 11849
rect 3120 11815 3154 11847
rect 3120 11745 3154 11777
rect 3120 11743 3154 11745
rect 3278 11847 3312 11849
rect 3278 11815 3312 11847
rect 3278 11745 3312 11777
rect 3278 11743 3312 11745
rect 3742 11857 3776 11859
rect 3742 11825 3776 11857
rect 3742 11755 3776 11787
rect 3742 11753 3776 11755
rect 3900 11857 3934 11859
rect 3900 11825 3934 11857
rect 3900 11755 3934 11787
rect 3900 11753 3934 11755
rect 4050 11857 4084 11859
rect 4050 11825 4084 11857
rect 4050 11755 4084 11787
rect 4050 11753 4084 11755
rect 4208 11857 4242 11859
rect 4208 11825 4242 11857
rect 4208 11755 4242 11787
rect 4208 11753 4242 11755
rect 4402 11857 4436 11859
rect 4402 11825 4436 11857
rect 4402 11755 4436 11787
rect 4402 11753 4436 11755
rect 4560 11857 4594 11859
rect 4560 11825 4594 11857
rect 4560 11755 4594 11787
rect 4560 11753 4594 11755
rect 4710 11857 4744 11859
rect 4710 11825 4744 11857
rect 4710 11755 4744 11787
rect 4710 11753 4744 11755
rect 4868 11857 4902 11859
rect 4868 11825 4902 11857
rect 4868 11755 4902 11787
rect 4868 11753 4902 11755
rect 5700 11858 5734 11860
rect 5700 11826 5734 11858
rect 5700 11756 5734 11788
rect 5700 11754 5734 11756
rect 5858 11858 5892 11860
rect 5858 11826 5892 11858
rect 5858 11756 5892 11788
rect 5858 11754 5892 11756
rect 6008 11858 6042 11860
rect 6008 11826 6042 11858
rect 6008 11756 6042 11788
rect 6008 11754 6042 11756
rect 6166 11858 6200 11860
rect 6166 11826 6200 11858
rect 6166 11756 6200 11788
rect 6166 11754 6200 11756
rect 6360 11858 6394 11860
rect 6360 11826 6394 11858
rect 6360 11756 6394 11788
rect 6360 11754 6394 11756
rect 6518 11858 6552 11860
rect 6518 11826 6552 11858
rect 6518 11756 6552 11788
rect 6518 11754 6552 11756
rect 6668 11858 6702 11860
rect 6668 11826 6702 11858
rect 6668 11756 6702 11788
rect 6668 11754 6702 11756
rect 6826 11858 6860 11860
rect 6826 11826 6860 11858
rect 6826 11756 6860 11788
rect 6826 11754 6860 11756
rect 2857 11605 2891 11639
rect 3670 11629 3704 11663
rect 3984 11620 4018 11654
rect 1410 11491 1444 11525
rect 565 11412 606 11436
rect 712 11412 753 11436
rect 856 11418 897 11441
rect 1568 11491 1602 11525
rect 1698 11491 1732 11525
rect 1856 11491 1890 11525
rect 2030 11491 2064 11525
rect 2188 11491 2222 11525
rect 2372 11491 2406 11525
rect 1010 11418 1051 11442
rect 565 11396 569 11412
rect 569 11396 603 11412
rect 603 11396 606 11412
rect 712 11396 715 11412
rect 715 11396 749 11412
rect 749 11396 753 11412
rect 856 11401 859 11418
rect 859 11401 893 11418
rect 893 11401 897 11418
rect 1010 11402 1013 11418
rect 1013 11402 1047 11418
rect 1047 11402 1051 11418
rect 1373 11314 1387 11348
rect 1387 11314 1407 11348
rect 1445 11314 1455 11348
rect 1455 11314 1479 11348
rect 1517 11314 1523 11348
rect 1523 11314 1551 11348
rect 1589 11314 1591 11348
rect 1591 11314 1623 11348
rect 1661 11314 1693 11348
rect 1693 11314 1695 11348
rect 1733 11314 1761 11348
rect 1761 11314 1767 11348
rect 1805 11314 1829 11348
rect 1829 11314 1839 11348
rect 1877 11314 1897 11348
rect 1897 11314 1911 11348
rect 2530 11491 2564 11525
rect 2369 11289 2403 11323
rect 4306 11614 4340 11648
rect 4637 11632 4671 11666
rect 5628 11630 5662 11664
rect 5942 11620 5976 11654
rect 6264 11614 6298 11648
rect 6596 11632 6630 11666
rect 2776 11491 2810 11525
rect 2934 11491 2968 11525
rect 3120 11491 3154 11525
rect 3278 11491 3312 11525
rect 3742 11501 3776 11535
rect 3900 11501 3934 11535
rect 4050 11501 4084 11535
rect 4208 11501 4242 11535
rect 4402 11503 4436 11537
rect 4560 11503 4594 11537
rect 4710 11503 4744 11537
rect 4868 11503 4902 11537
rect 5700 11502 5734 11536
rect 5858 11502 5892 11536
rect 6008 11502 6042 11536
rect 6166 11502 6200 11536
rect 6360 11504 6394 11538
rect 6518 11504 6552 11538
rect 6668 11504 6702 11538
rect 6826 11504 6860 11538
rect 3741 11325 3753 11359
rect 3753 11325 3775 11359
rect 3813 11325 3821 11359
rect 3821 11325 3847 11359
rect 3885 11325 3889 11359
rect 3889 11325 3919 11359
rect 3957 11325 3991 11359
rect 4029 11325 4059 11359
rect 4059 11325 4063 11359
rect 4101 11325 4127 11359
rect 4127 11325 4135 11359
rect 4173 11325 4195 11359
rect 4195 11325 4207 11359
rect 5700 11326 5712 11360
rect 5712 11326 5734 11360
rect 5772 11326 5780 11360
rect 5780 11326 5806 11360
rect 5844 11326 5848 11360
rect 5848 11326 5878 11360
rect 5916 11326 5950 11360
rect 5988 11326 6018 11360
rect 6018 11326 6022 11360
rect 6060 11326 6086 11360
rect 6086 11326 6094 11360
rect 6132 11326 6154 11360
rect 6154 11326 6166 11360
rect 2642 11173 2696 11227
rect 1383 10788 1395 10822
rect 1395 10788 1417 10822
rect 1455 10788 1463 10822
rect 1463 10788 1489 10822
rect 1527 10788 1531 10822
rect 1531 10788 1561 10822
rect 1599 10788 1633 10822
rect 1671 10788 1701 10822
rect 1701 10788 1705 10822
rect 1743 10788 1769 10822
rect 1769 10788 1777 10822
rect 1815 10788 1837 10822
rect 1837 10788 1849 10822
rect 566 10718 569 10736
rect 569 10718 603 10736
rect 603 10718 607 10736
rect 710 10718 715 10736
rect 715 10718 749 10736
rect 749 10718 751 10736
rect 856 10724 859 10741
rect 859 10724 893 10741
rect 893 10724 897 10741
rect 1009 10724 1013 10741
rect 1013 10724 1047 10741
rect 1047 10724 1050 10741
rect 566 10696 607 10718
rect 710 10696 751 10718
rect 856 10701 897 10724
rect 1009 10701 1050 10724
rect 1410 10619 1444 10621
rect 1410 10587 1444 10619
rect 1410 10517 1444 10549
rect 1410 10515 1444 10517
rect 1568 10619 1602 10621
rect 1568 10587 1602 10619
rect 1568 10517 1602 10549
rect 1568 10515 1602 10517
rect 1698 10619 1732 10621
rect 1698 10587 1732 10619
rect 1698 10517 1732 10549
rect 1698 10515 1732 10517
rect 1856 10619 1890 10621
rect 1856 10587 1890 10619
rect 1856 10517 1890 10549
rect 1856 10515 1890 10517
rect 2030 10619 2064 10621
rect 2030 10587 2064 10619
rect 2030 10517 2064 10549
rect 2030 10515 2064 10517
rect 2188 10619 2222 10621
rect 2188 10587 2222 10619
rect 2188 10517 2222 10549
rect 2188 10515 2222 10517
rect 2372 10619 2406 10621
rect 2372 10587 2406 10619
rect 2372 10517 2406 10549
rect 2372 10515 2406 10517
rect 2530 10619 2564 10621
rect 2530 10587 2564 10619
rect 2776 10619 2810 10621
rect 2530 10517 2564 10549
rect 2530 10515 2564 10517
rect 2647 10535 2681 10569
rect 2776 10587 2810 10619
rect 2776 10517 2810 10549
rect 2776 10515 2810 10517
rect 2934 10619 2968 10621
rect 2934 10587 2968 10619
rect 2934 10517 2968 10549
rect 2934 10515 2968 10517
rect 1269 10381 1303 10415
rect 1773 10381 1807 10415
rect 2273 10379 2307 10413
rect 3797 10787 3807 10821
rect 3807 10787 3831 10821
rect 3869 10787 3875 10821
rect 3875 10787 3903 10821
rect 3941 10787 3943 10821
rect 3943 10787 3975 10821
rect 4013 10787 4045 10821
rect 4045 10787 4047 10821
rect 4085 10787 4113 10821
rect 4113 10787 4119 10821
rect 4157 10787 4181 10821
rect 4181 10787 4191 10821
rect 5756 10786 5766 10820
rect 5766 10786 5790 10820
rect 5828 10786 5834 10820
rect 5834 10786 5862 10820
rect 5900 10786 5902 10820
rect 5902 10786 5934 10820
rect 5972 10786 6004 10820
rect 6004 10786 6006 10820
rect 6044 10786 6072 10820
rect 6072 10786 6078 10820
rect 6116 10786 6140 10820
rect 6140 10786 6150 10820
rect 3120 10619 3154 10621
rect 3120 10587 3154 10619
rect 3120 10517 3154 10549
rect 3120 10515 3154 10517
rect 3278 10619 3312 10621
rect 3278 10587 3312 10619
rect 3278 10517 3312 10549
rect 3278 10515 3312 10517
rect 3742 10629 3776 10631
rect 3742 10597 3776 10629
rect 3742 10527 3776 10559
rect 3742 10525 3776 10527
rect 3900 10629 3934 10631
rect 3900 10597 3934 10629
rect 3900 10527 3934 10559
rect 3900 10525 3934 10527
rect 4050 10629 4084 10631
rect 4050 10597 4084 10629
rect 4050 10527 4084 10559
rect 4050 10525 4084 10527
rect 4208 10629 4242 10631
rect 4208 10597 4242 10629
rect 4208 10527 4242 10559
rect 4208 10525 4242 10527
rect 4402 10629 4436 10631
rect 4402 10597 4436 10629
rect 4402 10527 4436 10559
rect 4402 10525 4436 10527
rect 4560 10629 4594 10631
rect 4560 10597 4594 10629
rect 4560 10527 4594 10559
rect 4560 10525 4594 10527
rect 4710 10629 4744 10631
rect 4710 10597 4744 10629
rect 4710 10527 4744 10559
rect 4710 10525 4744 10527
rect 4868 10629 4902 10631
rect 4868 10597 4902 10629
rect 4868 10527 4902 10559
rect 4868 10525 4902 10527
rect 5700 10630 5734 10632
rect 5700 10598 5734 10630
rect 5700 10528 5734 10560
rect 5700 10526 5734 10528
rect 5858 10630 5892 10632
rect 5858 10598 5892 10630
rect 5858 10528 5892 10560
rect 5858 10526 5892 10528
rect 6008 10630 6042 10632
rect 6008 10598 6042 10630
rect 6008 10528 6042 10560
rect 6008 10526 6042 10528
rect 6166 10630 6200 10632
rect 6166 10598 6200 10630
rect 6166 10528 6200 10560
rect 6166 10526 6200 10528
rect 6360 10630 6394 10632
rect 6360 10598 6394 10630
rect 6360 10528 6394 10560
rect 6360 10526 6394 10528
rect 6518 10630 6552 10632
rect 6518 10598 6552 10630
rect 6518 10528 6552 10560
rect 6518 10526 6552 10528
rect 6668 10630 6702 10632
rect 6668 10598 6702 10630
rect 6668 10528 6702 10560
rect 6668 10526 6702 10528
rect 6826 10630 6860 10632
rect 6826 10598 6860 10630
rect 6826 10528 6860 10560
rect 6826 10526 6860 10528
rect 2857 10377 2891 10411
rect 3670 10401 3704 10435
rect 3984 10392 4018 10426
rect 1410 10263 1444 10297
rect 565 10184 606 10208
rect 712 10184 753 10208
rect 856 10190 897 10213
rect 1568 10263 1602 10297
rect 1698 10263 1732 10297
rect 1856 10263 1890 10297
rect 2030 10263 2064 10297
rect 2188 10263 2222 10297
rect 2372 10263 2406 10297
rect 1010 10190 1051 10214
rect 565 10168 569 10184
rect 569 10168 603 10184
rect 603 10168 606 10184
rect 712 10168 715 10184
rect 715 10168 749 10184
rect 749 10168 753 10184
rect 856 10173 859 10190
rect 859 10173 893 10190
rect 893 10173 897 10190
rect 1010 10174 1013 10190
rect 1013 10174 1047 10190
rect 1047 10174 1051 10190
rect 1373 10086 1387 10120
rect 1387 10086 1407 10120
rect 1445 10086 1455 10120
rect 1455 10086 1479 10120
rect 1517 10086 1523 10120
rect 1523 10086 1551 10120
rect 1589 10086 1591 10120
rect 1591 10086 1623 10120
rect 1661 10086 1693 10120
rect 1693 10086 1695 10120
rect 1733 10086 1761 10120
rect 1761 10086 1767 10120
rect 1805 10086 1829 10120
rect 1829 10086 1839 10120
rect 1877 10086 1897 10120
rect 1897 10086 1911 10120
rect 2530 10263 2564 10297
rect 2369 10061 2403 10095
rect 4306 10386 4340 10420
rect 4637 10404 4671 10438
rect 5628 10402 5662 10436
rect 5942 10392 5976 10426
rect 6264 10386 6298 10420
rect 6596 10404 6630 10438
rect 2776 10263 2810 10297
rect 2934 10263 2968 10297
rect 3120 10263 3154 10297
rect 3278 10263 3312 10297
rect 3742 10273 3776 10307
rect 3900 10273 3934 10307
rect 4050 10273 4084 10307
rect 4208 10273 4242 10307
rect 4402 10275 4436 10309
rect 4560 10275 4594 10309
rect 4710 10275 4744 10309
rect 4868 10275 4902 10309
rect 5700 10274 5734 10308
rect 5858 10274 5892 10308
rect 6008 10274 6042 10308
rect 6166 10274 6200 10308
rect 6360 10276 6394 10310
rect 6518 10276 6552 10310
rect 6668 10276 6702 10310
rect 6826 10276 6860 10310
rect 3741 10097 3753 10131
rect 3753 10097 3775 10131
rect 3813 10097 3821 10131
rect 3821 10097 3847 10131
rect 3885 10097 3889 10131
rect 3889 10097 3919 10131
rect 3957 10097 3991 10131
rect 4029 10097 4059 10131
rect 4059 10097 4063 10131
rect 4101 10097 4127 10131
rect 4127 10097 4135 10131
rect 4173 10097 4195 10131
rect 4195 10097 4207 10131
rect 5700 10098 5712 10132
rect 5712 10098 5734 10132
rect 5772 10098 5780 10132
rect 5780 10098 5806 10132
rect 5844 10098 5848 10132
rect 5848 10098 5878 10132
rect 5916 10098 5950 10132
rect 5988 10098 6018 10132
rect 6018 10098 6022 10132
rect 6060 10098 6086 10132
rect 6086 10098 6094 10132
rect 6132 10098 6154 10132
rect 6154 10098 6166 10132
rect 2642 9945 2696 9999
rect 1383 9560 1395 9594
rect 1395 9560 1417 9594
rect 1455 9560 1463 9594
rect 1463 9560 1489 9594
rect 1527 9560 1531 9594
rect 1531 9560 1561 9594
rect 1599 9560 1633 9594
rect 1671 9560 1701 9594
rect 1701 9560 1705 9594
rect 1743 9560 1769 9594
rect 1769 9560 1777 9594
rect 1815 9560 1837 9594
rect 1837 9560 1849 9594
rect 566 9490 569 9508
rect 569 9490 603 9508
rect 603 9490 607 9508
rect 710 9490 715 9508
rect 715 9490 749 9508
rect 749 9490 751 9508
rect 856 9496 859 9513
rect 859 9496 893 9513
rect 893 9496 897 9513
rect 1009 9496 1013 9513
rect 1013 9496 1047 9513
rect 1047 9496 1050 9513
rect 566 9468 607 9490
rect 710 9468 751 9490
rect 856 9473 897 9496
rect 1009 9473 1050 9496
rect 1410 9391 1444 9393
rect 1410 9359 1444 9391
rect 1410 9289 1444 9321
rect 1410 9287 1444 9289
rect 1568 9391 1602 9393
rect 1568 9359 1602 9391
rect 1568 9289 1602 9321
rect 1568 9287 1602 9289
rect 1698 9391 1732 9393
rect 1698 9359 1732 9391
rect 1698 9289 1732 9321
rect 1698 9287 1732 9289
rect 1856 9391 1890 9393
rect 1856 9359 1890 9391
rect 1856 9289 1890 9321
rect 1856 9287 1890 9289
rect 2030 9391 2064 9393
rect 2030 9359 2064 9391
rect 2030 9289 2064 9321
rect 2030 9287 2064 9289
rect 2188 9391 2222 9393
rect 2188 9359 2222 9391
rect 2188 9289 2222 9321
rect 2188 9287 2222 9289
rect 2372 9391 2406 9393
rect 2372 9359 2406 9391
rect 2372 9289 2406 9321
rect 2372 9287 2406 9289
rect 2530 9391 2564 9393
rect 2530 9359 2564 9391
rect 2776 9391 2810 9393
rect 2530 9289 2564 9321
rect 2530 9287 2564 9289
rect 2647 9307 2681 9341
rect 2776 9359 2810 9391
rect 2776 9289 2810 9321
rect 2776 9287 2810 9289
rect 2934 9391 2968 9393
rect 2934 9359 2968 9391
rect 2934 9289 2968 9321
rect 2934 9287 2968 9289
rect 1269 9153 1303 9187
rect 1773 9153 1807 9187
rect 2273 9151 2307 9185
rect 3797 9559 3807 9593
rect 3807 9559 3831 9593
rect 3869 9559 3875 9593
rect 3875 9559 3903 9593
rect 3941 9559 3943 9593
rect 3943 9559 3975 9593
rect 4013 9559 4045 9593
rect 4045 9559 4047 9593
rect 4085 9559 4113 9593
rect 4113 9559 4119 9593
rect 4157 9559 4181 9593
rect 4181 9559 4191 9593
rect 5756 9558 5766 9592
rect 5766 9558 5790 9592
rect 5828 9558 5834 9592
rect 5834 9558 5862 9592
rect 5900 9558 5902 9592
rect 5902 9558 5934 9592
rect 5972 9558 6004 9592
rect 6004 9558 6006 9592
rect 6044 9558 6072 9592
rect 6072 9558 6078 9592
rect 6116 9558 6140 9592
rect 6140 9558 6150 9592
rect 3120 9391 3154 9393
rect 3120 9359 3154 9391
rect 3120 9289 3154 9321
rect 3120 9287 3154 9289
rect 3278 9391 3312 9393
rect 3278 9359 3312 9391
rect 3278 9289 3312 9321
rect 3278 9287 3312 9289
rect 3742 9401 3776 9403
rect 3742 9369 3776 9401
rect 3742 9299 3776 9331
rect 3742 9297 3776 9299
rect 3900 9401 3934 9403
rect 3900 9369 3934 9401
rect 3900 9299 3934 9331
rect 3900 9297 3934 9299
rect 4050 9401 4084 9403
rect 4050 9369 4084 9401
rect 4050 9299 4084 9331
rect 4050 9297 4084 9299
rect 4208 9401 4242 9403
rect 4208 9369 4242 9401
rect 4208 9299 4242 9331
rect 4208 9297 4242 9299
rect 4402 9401 4436 9403
rect 4402 9369 4436 9401
rect 4402 9299 4436 9331
rect 4402 9297 4436 9299
rect 4560 9401 4594 9403
rect 4560 9369 4594 9401
rect 4560 9299 4594 9331
rect 4560 9297 4594 9299
rect 4710 9401 4744 9403
rect 4710 9369 4744 9401
rect 4710 9299 4744 9331
rect 4710 9297 4744 9299
rect 4868 9401 4902 9403
rect 4868 9369 4902 9401
rect 4868 9299 4902 9331
rect 4868 9297 4902 9299
rect 5700 9402 5734 9404
rect 5700 9370 5734 9402
rect 5700 9300 5734 9332
rect 5700 9298 5734 9300
rect 5858 9402 5892 9404
rect 5858 9370 5892 9402
rect 5858 9300 5892 9332
rect 5858 9298 5892 9300
rect 6008 9402 6042 9404
rect 6008 9370 6042 9402
rect 6008 9300 6042 9332
rect 6008 9298 6042 9300
rect 6166 9402 6200 9404
rect 6166 9370 6200 9402
rect 6166 9300 6200 9332
rect 6166 9298 6200 9300
rect 6360 9402 6394 9404
rect 6360 9370 6394 9402
rect 6360 9300 6394 9332
rect 6360 9298 6394 9300
rect 6518 9402 6552 9404
rect 6518 9370 6552 9402
rect 6518 9300 6552 9332
rect 6518 9298 6552 9300
rect 6668 9402 6702 9404
rect 6668 9370 6702 9402
rect 6668 9300 6702 9332
rect 6668 9298 6702 9300
rect 6826 9402 6860 9404
rect 6826 9370 6860 9402
rect 6826 9300 6860 9332
rect 6826 9298 6860 9300
rect 2857 9149 2891 9183
rect 3670 9173 3704 9207
rect 3984 9164 4018 9198
rect 1410 9035 1444 9069
rect 565 8956 606 8980
rect 712 8956 753 8980
rect 856 8962 897 8985
rect 1568 9035 1602 9069
rect 1698 9035 1732 9069
rect 1856 9035 1890 9069
rect 2030 9035 2064 9069
rect 2188 9035 2222 9069
rect 2372 9035 2406 9069
rect 1010 8962 1051 8986
rect 565 8940 569 8956
rect 569 8940 603 8956
rect 603 8940 606 8956
rect 712 8940 715 8956
rect 715 8940 749 8956
rect 749 8940 753 8956
rect 856 8945 859 8962
rect 859 8945 893 8962
rect 893 8945 897 8962
rect 1010 8946 1013 8962
rect 1013 8946 1047 8962
rect 1047 8946 1051 8962
rect 1373 8858 1387 8892
rect 1387 8858 1407 8892
rect 1445 8858 1455 8892
rect 1455 8858 1479 8892
rect 1517 8858 1523 8892
rect 1523 8858 1551 8892
rect 1589 8858 1591 8892
rect 1591 8858 1623 8892
rect 1661 8858 1693 8892
rect 1693 8858 1695 8892
rect 1733 8858 1761 8892
rect 1761 8858 1767 8892
rect 1805 8858 1829 8892
rect 1829 8858 1839 8892
rect 1877 8858 1897 8892
rect 1897 8858 1911 8892
rect 2530 9035 2564 9069
rect 2369 8833 2403 8867
rect 4306 9158 4340 9192
rect 4637 9176 4671 9210
rect 5628 9174 5662 9208
rect 5942 9164 5976 9198
rect 6264 9158 6298 9192
rect 6596 9176 6630 9210
rect 2776 9035 2810 9069
rect 2934 9035 2968 9069
rect 3120 9035 3154 9069
rect 3278 9035 3312 9069
rect 3742 9045 3776 9079
rect 3900 9045 3934 9079
rect 4050 9045 4084 9079
rect 4208 9045 4242 9079
rect 4402 9047 4436 9081
rect 4560 9047 4594 9081
rect 4710 9047 4744 9081
rect 4868 9047 4902 9081
rect 5700 9046 5734 9080
rect 5858 9046 5892 9080
rect 6008 9046 6042 9080
rect 6166 9046 6200 9080
rect 6360 9048 6394 9082
rect 6518 9048 6552 9082
rect 6668 9048 6702 9082
rect 6826 9048 6860 9082
rect 3741 8869 3753 8903
rect 3753 8869 3775 8903
rect 3813 8869 3821 8903
rect 3821 8869 3847 8903
rect 3885 8869 3889 8903
rect 3889 8869 3919 8903
rect 3957 8869 3991 8903
rect 4029 8869 4059 8903
rect 4059 8869 4063 8903
rect 4101 8869 4127 8903
rect 4127 8869 4135 8903
rect 4173 8869 4195 8903
rect 4195 8869 4207 8903
rect 5700 8870 5712 8904
rect 5712 8870 5734 8904
rect 5772 8870 5780 8904
rect 5780 8870 5806 8904
rect 5844 8870 5848 8904
rect 5848 8870 5878 8904
rect 5916 8870 5950 8904
rect 5988 8870 6018 8904
rect 6018 8870 6022 8904
rect 6060 8870 6086 8904
rect 6086 8870 6094 8904
rect 6132 8870 6154 8904
rect 6154 8870 6166 8904
rect 2642 8717 2696 8771
rect 1383 8332 1395 8366
rect 1395 8332 1417 8366
rect 1455 8332 1463 8366
rect 1463 8332 1489 8366
rect 1527 8332 1531 8366
rect 1531 8332 1561 8366
rect 1599 8332 1633 8366
rect 1671 8332 1701 8366
rect 1701 8332 1705 8366
rect 1743 8332 1769 8366
rect 1769 8332 1777 8366
rect 1815 8332 1837 8366
rect 1837 8332 1849 8366
rect 566 8262 569 8280
rect 569 8262 603 8280
rect 603 8262 607 8280
rect 710 8262 715 8280
rect 715 8262 749 8280
rect 749 8262 751 8280
rect 856 8268 859 8285
rect 859 8268 893 8285
rect 893 8268 897 8285
rect 1009 8268 1013 8285
rect 1013 8268 1047 8285
rect 1047 8268 1050 8285
rect 566 8240 607 8262
rect 710 8240 751 8262
rect 856 8245 897 8268
rect 1009 8245 1050 8268
rect 1410 8163 1444 8165
rect 1410 8131 1444 8163
rect 1410 8061 1444 8093
rect 1410 8059 1444 8061
rect 1568 8163 1602 8165
rect 1568 8131 1602 8163
rect 1568 8061 1602 8093
rect 1568 8059 1602 8061
rect 1698 8163 1732 8165
rect 1698 8131 1732 8163
rect 1698 8061 1732 8093
rect 1698 8059 1732 8061
rect 1856 8163 1890 8165
rect 1856 8131 1890 8163
rect 1856 8061 1890 8093
rect 1856 8059 1890 8061
rect 2030 8163 2064 8165
rect 2030 8131 2064 8163
rect 2030 8061 2064 8093
rect 2030 8059 2064 8061
rect 2188 8163 2222 8165
rect 2188 8131 2222 8163
rect 2188 8061 2222 8093
rect 2188 8059 2222 8061
rect 2372 8163 2406 8165
rect 2372 8131 2406 8163
rect 2372 8061 2406 8093
rect 2372 8059 2406 8061
rect 2530 8163 2564 8165
rect 2530 8131 2564 8163
rect 2776 8163 2810 8165
rect 2530 8061 2564 8093
rect 2530 8059 2564 8061
rect 2647 8079 2681 8113
rect 2776 8131 2810 8163
rect 2776 8061 2810 8093
rect 2776 8059 2810 8061
rect 2934 8163 2968 8165
rect 2934 8131 2968 8163
rect 2934 8061 2968 8093
rect 2934 8059 2968 8061
rect 1269 7925 1303 7959
rect 1773 7925 1807 7959
rect 2273 7923 2307 7957
rect 3797 8331 3807 8365
rect 3807 8331 3831 8365
rect 3869 8331 3875 8365
rect 3875 8331 3903 8365
rect 3941 8331 3943 8365
rect 3943 8331 3975 8365
rect 4013 8331 4045 8365
rect 4045 8331 4047 8365
rect 4085 8331 4113 8365
rect 4113 8331 4119 8365
rect 4157 8331 4181 8365
rect 4181 8331 4191 8365
rect 5756 8330 5766 8364
rect 5766 8330 5790 8364
rect 5828 8330 5834 8364
rect 5834 8330 5862 8364
rect 5900 8330 5902 8364
rect 5902 8330 5934 8364
rect 5972 8330 6004 8364
rect 6004 8330 6006 8364
rect 6044 8330 6072 8364
rect 6072 8330 6078 8364
rect 6116 8330 6140 8364
rect 6140 8330 6150 8364
rect 3120 8163 3154 8165
rect 3120 8131 3154 8163
rect 3120 8061 3154 8093
rect 3120 8059 3154 8061
rect 3278 8163 3312 8165
rect 3278 8131 3312 8163
rect 3278 8061 3312 8093
rect 3278 8059 3312 8061
rect 3742 8173 3776 8175
rect 3742 8141 3776 8173
rect 3742 8071 3776 8103
rect 3742 8069 3776 8071
rect 3900 8173 3934 8175
rect 3900 8141 3934 8173
rect 3900 8071 3934 8103
rect 3900 8069 3934 8071
rect 4050 8173 4084 8175
rect 4050 8141 4084 8173
rect 4050 8071 4084 8103
rect 4050 8069 4084 8071
rect 4208 8173 4242 8175
rect 4208 8141 4242 8173
rect 4208 8071 4242 8103
rect 4208 8069 4242 8071
rect 4402 8173 4436 8175
rect 4402 8141 4436 8173
rect 4402 8071 4436 8103
rect 4402 8069 4436 8071
rect 4560 8173 4594 8175
rect 4560 8141 4594 8173
rect 4560 8071 4594 8103
rect 4560 8069 4594 8071
rect 4710 8173 4744 8175
rect 4710 8141 4744 8173
rect 4710 8071 4744 8103
rect 4710 8069 4744 8071
rect 4868 8173 4902 8175
rect 4868 8141 4902 8173
rect 4868 8071 4902 8103
rect 4868 8069 4902 8071
rect 5700 8174 5734 8176
rect 5700 8142 5734 8174
rect 5700 8072 5734 8104
rect 5700 8070 5734 8072
rect 5858 8174 5892 8176
rect 5858 8142 5892 8174
rect 5858 8072 5892 8104
rect 5858 8070 5892 8072
rect 6008 8174 6042 8176
rect 6008 8142 6042 8174
rect 6008 8072 6042 8104
rect 6008 8070 6042 8072
rect 6166 8174 6200 8176
rect 6166 8142 6200 8174
rect 6166 8072 6200 8104
rect 6166 8070 6200 8072
rect 6360 8174 6394 8176
rect 6360 8142 6394 8174
rect 6360 8072 6394 8104
rect 6360 8070 6394 8072
rect 6518 8174 6552 8176
rect 6518 8142 6552 8174
rect 6518 8072 6552 8104
rect 6518 8070 6552 8072
rect 6668 8174 6702 8176
rect 6668 8142 6702 8174
rect 6668 8072 6702 8104
rect 6668 8070 6702 8072
rect 6826 8174 6860 8176
rect 6826 8142 6860 8174
rect 6826 8072 6860 8104
rect 6826 8070 6860 8072
rect 2857 7921 2891 7955
rect 3670 7945 3704 7979
rect 3984 7936 4018 7970
rect 1410 7807 1444 7841
rect 565 7728 606 7752
rect 712 7728 753 7752
rect 856 7734 897 7757
rect 1568 7807 1602 7841
rect 1698 7807 1732 7841
rect 1856 7807 1890 7841
rect 2030 7807 2064 7841
rect 2188 7807 2222 7841
rect 2372 7807 2406 7841
rect 1010 7734 1051 7758
rect 565 7712 569 7728
rect 569 7712 603 7728
rect 603 7712 606 7728
rect 712 7712 715 7728
rect 715 7712 749 7728
rect 749 7712 753 7728
rect 856 7717 859 7734
rect 859 7717 893 7734
rect 893 7717 897 7734
rect 1010 7718 1013 7734
rect 1013 7718 1047 7734
rect 1047 7718 1051 7734
rect 1373 7630 1387 7664
rect 1387 7630 1407 7664
rect 1445 7630 1455 7664
rect 1455 7630 1479 7664
rect 1517 7630 1523 7664
rect 1523 7630 1551 7664
rect 1589 7630 1591 7664
rect 1591 7630 1623 7664
rect 1661 7630 1693 7664
rect 1693 7630 1695 7664
rect 1733 7630 1761 7664
rect 1761 7630 1767 7664
rect 1805 7630 1829 7664
rect 1829 7630 1839 7664
rect 1877 7630 1897 7664
rect 1897 7630 1911 7664
rect 2530 7807 2564 7841
rect 2369 7605 2403 7639
rect 4306 7930 4340 7964
rect 4637 7948 4671 7982
rect 5628 7946 5662 7980
rect 5942 7936 5976 7970
rect 6264 7930 6298 7964
rect 6596 7948 6630 7982
rect 2776 7807 2810 7841
rect 2934 7807 2968 7841
rect 3120 7807 3154 7841
rect 3278 7807 3312 7841
rect 3742 7817 3776 7851
rect 3900 7817 3934 7851
rect 4050 7817 4084 7851
rect 4208 7817 4242 7851
rect 4402 7819 4436 7853
rect 4560 7819 4594 7853
rect 4710 7819 4744 7853
rect 4868 7819 4902 7853
rect 5700 7818 5734 7852
rect 5858 7818 5892 7852
rect 6008 7818 6042 7852
rect 6166 7818 6200 7852
rect 6360 7820 6394 7854
rect 6518 7820 6552 7854
rect 6668 7820 6702 7854
rect 6826 7820 6860 7854
rect 3741 7641 3753 7675
rect 3753 7641 3775 7675
rect 3813 7641 3821 7675
rect 3821 7641 3847 7675
rect 3885 7641 3889 7675
rect 3889 7641 3919 7675
rect 3957 7641 3991 7675
rect 4029 7641 4059 7675
rect 4059 7641 4063 7675
rect 4101 7641 4127 7675
rect 4127 7641 4135 7675
rect 4173 7641 4195 7675
rect 4195 7641 4207 7675
rect 5700 7642 5712 7676
rect 5712 7642 5734 7676
rect 5772 7642 5780 7676
rect 5780 7642 5806 7676
rect 5844 7642 5848 7676
rect 5848 7642 5878 7676
rect 5916 7642 5950 7676
rect 5988 7642 6018 7676
rect 6018 7642 6022 7676
rect 6060 7642 6086 7676
rect 6086 7642 6094 7676
rect 6132 7642 6154 7676
rect 6154 7642 6166 7676
rect 2642 7489 2696 7543
rect 1383 7104 1395 7138
rect 1395 7104 1417 7138
rect 1455 7104 1463 7138
rect 1463 7104 1489 7138
rect 1527 7104 1531 7138
rect 1531 7104 1561 7138
rect 1599 7104 1633 7138
rect 1671 7104 1701 7138
rect 1701 7104 1705 7138
rect 1743 7104 1769 7138
rect 1769 7104 1777 7138
rect 1815 7104 1837 7138
rect 1837 7104 1849 7138
rect 566 7034 569 7052
rect 569 7034 603 7052
rect 603 7034 607 7052
rect 710 7034 715 7052
rect 715 7034 749 7052
rect 749 7034 751 7052
rect 856 7040 859 7057
rect 859 7040 893 7057
rect 893 7040 897 7057
rect 1009 7040 1013 7057
rect 1013 7040 1047 7057
rect 1047 7040 1050 7057
rect 566 7012 607 7034
rect 710 7012 751 7034
rect 856 7017 897 7040
rect 1009 7017 1050 7040
rect 1410 6935 1444 6937
rect 1410 6903 1444 6935
rect 1410 6833 1444 6865
rect 1410 6831 1444 6833
rect 1568 6935 1602 6937
rect 1568 6903 1602 6935
rect 1568 6833 1602 6865
rect 1568 6831 1602 6833
rect 1698 6935 1732 6937
rect 1698 6903 1732 6935
rect 1698 6833 1732 6865
rect 1698 6831 1732 6833
rect 1856 6935 1890 6937
rect 1856 6903 1890 6935
rect 1856 6833 1890 6865
rect 1856 6831 1890 6833
rect 2030 6935 2064 6937
rect 2030 6903 2064 6935
rect 2030 6833 2064 6865
rect 2030 6831 2064 6833
rect 2188 6935 2222 6937
rect 2188 6903 2222 6935
rect 2188 6833 2222 6865
rect 2188 6831 2222 6833
rect 2372 6935 2406 6937
rect 2372 6903 2406 6935
rect 2372 6833 2406 6865
rect 2372 6831 2406 6833
rect 2530 6935 2564 6937
rect 2530 6903 2564 6935
rect 2776 6935 2810 6937
rect 2530 6833 2564 6865
rect 2530 6831 2564 6833
rect 2647 6851 2681 6885
rect 2776 6903 2810 6935
rect 2776 6833 2810 6865
rect 2776 6831 2810 6833
rect 2934 6935 2968 6937
rect 2934 6903 2968 6935
rect 2934 6833 2968 6865
rect 2934 6831 2968 6833
rect 1269 6697 1303 6731
rect 1773 6697 1807 6731
rect 2273 6695 2307 6729
rect 3797 7103 3807 7137
rect 3807 7103 3831 7137
rect 3869 7103 3875 7137
rect 3875 7103 3903 7137
rect 3941 7103 3943 7137
rect 3943 7103 3975 7137
rect 4013 7103 4045 7137
rect 4045 7103 4047 7137
rect 4085 7103 4113 7137
rect 4113 7103 4119 7137
rect 4157 7103 4181 7137
rect 4181 7103 4191 7137
rect 5756 7102 5766 7136
rect 5766 7102 5790 7136
rect 5828 7102 5834 7136
rect 5834 7102 5862 7136
rect 5900 7102 5902 7136
rect 5902 7102 5934 7136
rect 5972 7102 6004 7136
rect 6004 7102 6006 7136
rect 6044 7102 6072 7136
rect 6072 7102 6078 7136
rect 6116 7102 6140 7136
rect 6140 7102 6150 7136
rect 3120 6935 3154 6937
rect 3120 6903 3154 6935
rect 3120 6833 3154 6865
rect 3120 6831 3154 6833
rect 3278 6935 3312 6937
rect 3278 6903 3312 6935
rect 3278 6833 3312 6865
rect 3278 6831 3312 6833
rect 3742 6945 3776 6947
rect 3742 6913 3776 6945
rect 3742 6843 3776 6875
rect 3742 6841 3776 6843
rect 3900 6945 3934 6947
rect 3900 6913 3934 6945
rect 3900 6843 3934 6875
rect 3900 6841 3934 6843
rect 4050 6945 4084 6947
rect 4050 6913 4084 6945
rect 4050 6843 4084 6875
rect 4050 6841 4084 6843
rect 4208 6945 4242 6947
rect 4208 6913 4242 6945
rect 4208 6843 4242 6875
rect 4208 6841 4242 6843
rect 4402 6945 4436 6947
rect 4402 6913 4436 6945
rect 4402 6843 4436 6875
rect 4402 6841 4436 6843
rect 4560 6945 4594 6947
rect 4560 6913 4594 6945
rect 4560 6843 4594 6875
rect 4560 6841 4594 6843
rect 4710 6945 4744 6947
rect 4710 6913 4744 6945
rect 4710 6843 4744 6875
rect 4710 6841 4744 6843
rect 4868 6945 4902 6947
rect 4868 6913 4902 6945
rect 4868 6843 4902 6875
rect 4868 6841 4902 6843
rect 5700 6946 5734 6948
rect 5700 6914 5734 6946
rect 5700 6844 5734 6876
rect 5700 6842 5734 6844
rect 5858 6946 5892 6948
rect 5858 6914 5892 6946
rect 5858 6844 5892 6876
rect 5858 6842 5892 6844
rect 6008 6946 6042 6948
rect 6008 6914 6042 6946
rect 6008 6844 6042 6876
rect 6008 6842 6042 6844
rect 6166 6946 6200 6948
rect 6166 6914 6200 6946
rect 6166 6844 6200 6876
rect 6166 6842 6200 6844
rect 6360 6946 6394 6948
rect 6360 6914 6394 6946
rect 6360 6844 6394 6876
rect 6360 6842 6394 6844
rect 6518 6946 6552 6948
rect 6518 6914 6552 6946
rect 6518 6844 6552 6876
rect 6518 6842 6552 6844
rect 6668 6946 6702 6948
rect 6668 6914 6702 6946
rect 6668 6844 6702 6876
rect 6668 6842 6702 6844
rect 6826 6946 6860 6948
rect 6826 6914 6860 6946
rect 6826 6844 6860 6876
rect 6826 6842 6860 6844
rect 2857 6693 2891 6727
rect 3670 6717 3704 6751
rect 3984 6708 4018 6742
rect 1410 6579 1444 6613
rect 565 6500 606 6524
rect 712 6500 753 6524
rect 856 6506 897 6529
rect 1568 6579 1602 6613
rect 1698 6579 1732 6613
rect 1856 6579 1890 6613
rect 2030 6579 2064 6613
rect 2188 6579 2222 6613
rect 2372 6579 2406 6613
rect 1010 6506 1051 6530
rect 565 6484 569 6500
rect 569 6484 603 6500
rect 603 6484 606 6500
rect 712 6484 715 6500
rect 715 6484 749 6500
rect 749 6484 753 6500
rect 856 6489 859 6506
rect 859 6489 893 6506
rect 893 6489 897 6506
rect 1010 6490 1013 6506
rect 1013 6490 1047 6506
rect 1047 6490 1051 6506
rect 1373 6402 1387 6436
rect 1387 6402 1407 6436
rect 1445 6402 1455 6436
rect 1455 6402 1479 6436
rect 1517 6402 1523 6436
rect 1523 6402 1551 6436
rect 1589 6402 1591 6436
rect 1591 6402 1623 6436
rect 1661 6402 1693 6436
rect 1693 6402 1695 6436
rect 1733 6402 1761 6436
rect 1761 6402 1767 6436
rect 1805 6402 1829 6436
rect 1829 6402 1839 6436
rect 1877 6402 1897 6436
rect 1897 6402 1911 6436
rect 2530 6579 2564 6613
rect 2369 6377 2403 6411
rect 4306 6702 4340 6736
rect 4637 6720 4671 6754
rect 5628 6718 5662 6752
rect 5942 6708 5976 6742
rect 6264 6702 6298 6736
rect 6596 6720 6630 6754
rect 2776 6579 2810 6613
rect 2934 6579 2968 6613
rect 3120 6579 3154 6613
rect 3278 6579 3312 6613
rect 3742 6589 3776 6623
rect 3900 6589 3934 6623
rect 4050 6589 4084 6623
rect 4208 6589 4242 6623
rect 4402 6591 4436 6625
rect 4560 6591 4594 6625
rect 4710 6591 4744 6625
rect 4868 6591 4902 6625
rect 5700 6590 5734 6624
rect 5858 6590 5892 6624
rect 6008 6590 6042 6624
rect 6166 6590 6200 6624
rect 6360 6592 6394 6626
rect 6518 6592 6552 6626
rect 6668 6592 6702 6626
rect 6826 6592 6860 6626
rect 3741 6413 3753 6447
rect 3753 6413 3775 6447
rect 3813 6413 3821 6447
rect 3821 6413 3847 6447
rect 3885 6413 3889 6447
rect 3889 6413 3919 6447
rect 3957 6413 3991 6447
rect 4029 6413 4059 6447
rect 4059 6413 4063 6447
rect 4101 6413 4127 6447
rect 4127 6413 4135 6447
rect 4173 6413 4195 6447
rect 4195 6413 4207 6447
rect 5700 6414 5712 6448
rect 5712 6414 5734 6448
rect 5772 6414 5780 6448
rect 5780 6414 5806 6448
rect 5844 6414 5848 6448
rect 5848 6414 5878 6448
rect 5916 6414 5950 6448
rect 5988 6414 6018 6448
rect 6018 6414 6022 6448
rect 6060 6414 6086 6448
rect 6086 6414 6094 6448
rect 6132 6414 6154 6448
rect 6154 6414 6166 6448
rect 2642 6261 2696 6315
rect 1383 5876 1395 5910
rect 1395 5876 1417 5910
rect 1455 5876 1463 5910
rect 1463 5876 1489 5910
rect 1527 5876 1531 5910
rect 1531 5876 1561 5910
rect 1599 5876 1633 5910
rect 1671 5876 1701 5910
rect 1701 5876 1705 5910
rect 1743 5876 1769 5910
rect 1769 5876 1777 5910
rect 1815 5876 1837 5910
rect 1837 5876 1849 5910
rect 566 5806 569 5824
rect 569 5806 603 5824
rect 603 5806 607 5824
rect 710 5806 715 5824
rect 715 5806 749 5824
rect 749 5806 751 5824
rect 856 5812 859 5829
rect 859 5812 893 5829
rect 893 5812 897 5829
rect 1009 5812 1013 5829
rect 1013 5812 1047 5829
rect 1047 5812 1050 5829
rect 566 5784 607 5806
rect 710 5784 751 5806
rect 856 5789 897 5812
rect 1009 5789 1050 5812
rect 1410 5707 1444 5709
rect 1410 5675 1444 5707
rect 1410 5605 1444 5637
rect 1410 5603 1444 5605
rect 1568 5707 1602 5709
rect 1568 5675 1602 5707
rect 1568 5605 1602 5637
rect 1568 5603 1602 5605
rect 1698 5707 1732 5709
rect 1698 5675 1732 5707
rect 1698 5605 1732 5637
rect 1698 5603 1732 5605
rect 1856 5707 1890 5709
rect 1856 5675 1890 5707
rect 1856 5605 1890 5637
rect 1856 5603 1890 5605
rect 2030 5707 2064 5709
rect 2030 5675 2064 5707
rect 2030 5605 2064 5637
rect 2030 5603 2064 5605
rect 2188 5707 2222 5709
rect 2188 5675 2222 5707
rect 2188 5605 2222 5637
rect 2188 5603 2222 5605
rect 2372 5707 2406 5709
rect 2372 5675 2406 5707
rect 2372 5605 2406 5637
rect 2372 5603 2406 5605
rect 2530 5707 2564 5709
rect 2530 5675 2564 5707
rect 2776 5707 2810 5709
rect 2530 5605 2564 5637
rect 2530 5603 2564 5605
rect 2647 5623 2681 5657
rect 2776 5675 2810 5707
rect 2776 5605 2810 5637
rect 2776 5603 2810 5605
rect 2934 5707 2968 5709
rect 2934 5675 2968 5707
rect 2934 5605 2968 5637
rect 2934 5603 2968 5605
rect 1269 5469 1303 5503
rect 1773 5469 1807 5503
rect 2273 5467 2307 5501
rect 3797 5875 3807 5909
rect 3807 5875 3831 5909
rect 3869 5875 3875 5909
rect 3875 5875 3903 5909
rect 3941 5875 3943 5909
rect 3943 5875 3975 5909
rect 4013 5875 4045 5909
rect 4045 5875 4047 5909
rect 4085 5875 4113 5909
rect 4113 5875 4119 5909
rect 4157 5875 4181 5909
rect 4181 5875 4191 5909
rect 5756 5874 5766 5908
rect 5766 5874 5790 5908
rect 5828 5874 5834 5908
rect 5834 5874 5862 5908
rect 5900 5874 5902 5908
rect 5902 5874 5934 5908
rect 5972 5874 6004 5908
rect 6004 5874 6006 5908
rect 6044 5874 6072 5908
rect 6072 5874 6078 5908
rect 6116 5874 6140 5908
rect 6140 5874 6150 5908
rect 3120 5707 3154 5709
rect 3120 5675 3154 5707
rect 3120 5605 3154 5637
rect 3120 5603 3154 5605
rect 3278 5707 3312 5709
rect 3278 5675 3312 5707
rect 3278 5605 3312 5637
rect 3278 5603 3312 5605
rect 3742 5717 3776 5719
rect 3742 5685 3776 5717
rect 3742 5615 3776 5647
rect 3742 5613 3776 5615
rect 3900 5717 3934 5719
rect 3900 5685 3934 5717
rect 3900 5615 3934 5647
rect 3900 5613 3934 5615
rect 4050 5717 4084 5719
rect 4050 5685 4084 5717
rect 4050 5615 4084 5647
rect 4050 5613 4084 5615
rect 4208 5717 4242 5719
rect 4208 5685 4242 5717
rect 4208 5615 4242 5647
rect 4208 5613 4242 5615
rect 4402 5717 4436 5719
rect 4402 5685 4436 5717
rect 4402 5615 4436 5647
rect 4402 5613 4436 5615
rect 4560 5717 4594 5719
rect 4560 5685 4594 5717
rect 4560 5615 4594 5647
rect 4560 5613 4594 5615
rect 4710 5717 4744 5719
rect 4710 5685 4744 5717
rect 4710 5615 4744 5647
rect 4710 5613 4744 5615
rect 4868 5717 4902 5719
rect 4868 5685 4902 5717
rect 4868 5615 4902 5647
rect 4868 5613 4902 5615
rect 5700 5718 5734 5720
rect 5700 5686 5734 5718
rect 5700 5616 5734 5648
rect 5700 5614 5734 5616
rect 5858 5718 5892 5720
rect 5858 5686 5892 5718
rect 5858 5616 5892 5648
rect 5858 5614 5892 5616
rect 6008 5718 6042 5720
rect 6008 5686 6042 5718
rect 6008 5616 6042 5648
rect 6008 5614 6042 5616
rect 6166 5718 6200 5720
rect 6166 5686 6200 5718
rect 6166 5616 6200 5648
rect 6166 5614 6200 5616
rect 6360 5718 6394 5720
rect 6360 5686 6394 5718
rect 6360 5616 6394 5648
rect 6360 5614 6394 5616
rect 6518 5718 6552 5720
rect 6518 5686 6552 5718
rect 6518 5616 6552 5648
rect 6518 5614 6552 5616
rect 6668 5718 6702 5720
rect 6668 5686 6702 5718
rect 6668 5616 6702 5648
rect 6668 5614 6702 5616
rect 6826 5718 6860 5720
rect 6826 5686 6860 5718
rect 6826 5616 6860 5648
rect 6826 5614 6860 5616
rect 2857 5465 2891 5499
rect 3670 5489 3704 5523
rect 3984 5480 4018 5514
rect 1410 5351 1444 5385
rect 565 5272 606 5296
rect 712 5272 753 5296
rect 856 5278 897 5301
rect 1568 5351 1602 5385
rect 1698 5351 1732 5385
rect 1856 5351 1890 5385
rect 2030 5351 2064 5385
rect 2188 5351 2222 5385
rect 2372 5351 2406 5385
rect 1010 5278 1051 5302
rect 565 5256 569 5272
rect 569 5256 603 5272
rect 603 5256 606 5272
rect 712 5256 715 5272
rect 715 5256 749 5272
rect 749 5256 753 5272
rect 856 5261 859 5278
rect 859 5261 893 5278
rect 893 5261 897 5278
rect 1010 5262 1013 5278
rect 1013 5262 1047 5278
rect 1047 5262 1051 5278
rect 1373 5174 1387 5208
rect 1387 5174 1407 5208
rect 1445 5174 1455 5208
rect 1455 5174 1479 5208
rect 1517 5174 1523 5208
rect 1523 5174 1551 5208
rect 1589 5174 1591 5208
rect 1591 5174 1623 5208
rect 1661 5174 1693 5208
rect 1693 5174 1695 5208
rect 1733 5174 1761 5208
rect 1761 5174 1767 5208
rect 1805 5174 1829 5208
rect 1829 5174 1839 5208
rect 1877 5174 1897 5208
rect 1897 5174 1911 5208
rect 2530 5351 2564 5385
rect 2369 5149 2403 5183
rect 4306 5474 4340 5508
rect 4637 5492 4671 5526
rect 5628 5490 5662 5524
rect 5942 5480 5976 5514
rect 6264 5474 6298 5508
rect 6596 5492 6630 5526
rect 2776 5351 2810 5385
rect 2934 5351 2968 5385
rect 3120 5351 3154 5385
rect 3278 5351 3312 5385
rect 3742 5361 3776 5395
rect 3900 5361 3934 5395
rect 4050 5361 4084 5395
rect 4208 5361 4242 5395
rect 4402 5363 4436 5397
rect 4560 5363 4594 5397
rect 4710 5363 4744 5397
rect 4868 5363 4902 5397
rect 5700 5362 5734 5396
rect 5858 5362 5892 5396
rect 6008 5362 6042 5396
rect 6166 5362 6200 5396
rect 6360 5364 6394 5398
rect 6518 5364 6552 5398
rect 6668 5364 6702 5398
rect 6826 5364 6860 5398
rect 3741 5185 3753 5219
rect 3753 5185 3775 5219
rect 3813 5185 3821 5219
rect 3821 5185 3847 5219
rect 3885 5185 3889 5219
rect 3889 5185 3919 5219
rect 3957 5185 3991 5219
rect 4029 5185 4059 5219
rect 4059 5185 4063 5219
rect 4101 5185 4127 5219
rect 4127 5185 4135 5219
rect 4173 5185 4195 5219
rect 4195 5185 4207 5219
rect 5700 5186 5712 5220
rect 5712 5186 5734 5220
rect 5772 5186 5780 5220
rect 5780 5186 5806 5220
rect 5844 5186 5848 5220
rect 5848 5186 5878 5220
rect 5916 5186 5950 5220
rect 5988 5186 6018 5220
rect 6018 5186 6022 5220
rect 6060 5186 6086 5220
rect 6086 5186 6094 5220
rect 6132 5186 6154 5220
rect 6154 5186 6166 5220
rect 2642 5033 2696 5087
rect 1383 4648 1395 4682
rect 1395 4648 1417 4682
rect 1455 4648 1463 4682
rect 1463 4648 1489 4682
rect 1527 4648 1531 4682
rect 1531 4648 1561 4682
rect 1599 4648 1633 4682
rect 1671 4648 1701 4682
rect 1701 4648 1705 4682
rect 1743 4648 1769 4682
rect 1769 4648 1777 4682
rect 1815 4648 1837 4682
rect 1837 4648 1849 4682
rect 566 4578 569 4596
rect 569 4578 603 4596
rect 603 4578 607 4596
rect 710 4578 715 4596
rect 715 4578 749 4596
rect 749 4578 751 4596
rect 856 4584 859 4601
rect 859 4584 893 4601
rect 893 4584 897 4601
rect 1009 4584 1013 4601
rect 1013 4584 1047 4601
rect 1047 4584 1050 4601
rect 566 4556 607 4578
rect 710 4556 751 4578
rect 856 4561 897 4584
rect 1009 4561 1050 4584
rect 1410 4479 1444 4481
rect 1410 4447 1444 4479
rect 1410 4377 1444 4409
rect 1410 4375 1444 4377
rect 1568 4479 1602 4481
rect 1568 4447 1602 4479
rect 1568 4377 1602 4409
rect 1568 4375 1602 4377
rect 1698 4479 1732 4481
rect 1698 4447 1732 4479
rect 1698 4377 1732 4409
rect 1698 4375 1732 4377
rect 1856 4479 1890 4481
rect 1856 4447 1890 4479
rect 1856 4377 1890 4409
rect 1856 4375 1890 4377
rect 2030 4479 2064 4481
rect 2030 4447 2064 4479
rect 2030 4377 2064 4409
rect 2030 4375 2064 4377
rect 2188 4479 2222 4481
rect 2188 4447 2222 4479
rect 2188 4377 2222 4409
rect 2188 4375 2222 4377
rect 2372 4479 2406 4481
rect 2372 4447 2406 4479
rect 2372 4377 2406 4409
rect 2372 4375 2406 4377
rect 2530 4479 2564 4481
rect 2530 4447 2564 4479
rect 2776 4479 2810 4481
rect 2530 4377 2564 4409
rect 2530 4375 2564 4377
rect 2647 4395 2681 4429
rect 2776 4447 2810 4479
rect 2776 4377 2810 4409
rect 2776 4375 2810 4377
rect 2934 4479 2968 4481
rect 2934 4447 2968 4479
rect 2934 4377 2968 4409
rect 2934 4375 2968 4377
rect 1269 4241 1303 4275
rect 1773 4241 1807 4275
rect 2273 4239 2307 4273
rect 3797 4647 3807 4681
rect 3807 4647 3831 4681
rect 3869 4647 3875 4681
rect 3875 4647 3903 4681
rect 3941 4647 3943 4681
rect 3943 4647 3975 4681
rect 4013 4647 4045 4681
rect 4045 4647 4047 4681
rect 4085 4647 4113 4681
rect 4113 4647 4119 4681
rect 4157 4647 4181 4681
rect 4181 4647 4191 4681
rect 5756 4646 5766 4680
rect 5766 4646 5790 4680
rect 5828 4646 5834 4680
rect 5834 4646 5862 4680
rect 5900 4646 5902 4680
rect 5902 4646 5934 4680
rect 5972 4646 6004 4680
rect 6004 4646 6006 4680
rect 6044 4646 6072 4680
rect 6072 4646 6078 4680
rect 6116 4646 6140 4680
rect 6140 4646 6150 4680
rect 3120 4479 3154 4481
rect 3120 4447 3154 4479
rect 3120 4377 3154 4409
rect 3120 4375 3154 4377
rect 3278 4479 3312 4481
rect 3278 4447 3312 4479
rect 3278 4377 3312 4409
rect 3278 4375 3312 4377
rect 3742 4489 3776 4491
rect 3742 4457 3776 4489
rect 3742 4387 3776 4419
rect 3742 4385 3776 4387
rect 3900 4489 3934 4491
rect 3900 4457 3934 4489
rect 3900 4387 3934 4419
rect 3900 4385 3934 4387
rect 4050 4489 4084 4491
rect 4050 4457 4084 4489
rect 4050 4387 4084 4419
rect 4050 4385 4084 4387
rect 4208 4489 4242 4491
rect 4208 4457 4242 4489
rect 4208 4387 4242 4419
rect 4208 4385 4242 4387
rect 4402 4489 4436 4491
rect 4402 4457 4436 4489
rect 4402 4387 4436 4419
rect 4402 4385 4436 4387
rect 4560 4489 4594 4491
rect 4560 4457 4594 4489
rect 4560 4387 4594 4419
rect 4560 4385 4594 4387
rect 4710 4489 4744 4491
rect 4710 4457 4744 4489
rect 4710 4387 4744 4419
rect 4710 4385 4744 4387
rect 4868 4489 4902 4491
rect 4868 4457 4902 4489
rect 4868 4387 4902 4419
rect 4868 4385 4902 4387
rect 5700 4490 5734 4492
rect 5700 4458 5734 4490
rect 5700 4388 5734 4420
rect 5700 4386 5734 4388
rect 5858 4490 5892 4492
rect 5858 4458 5892 4490
rect 5858 4388 5892 4420
rect 5858 4386 5892 4388
rect 6008 4490 6042 4492
rect 6008 4458 6042 4490
rect 6008 4388 6042 4420
rect 6008 4386 6042 4388
rect 6166 4490 6200 4492
rect 6166 4458 6200 4490
rect 6166 4388 6200 4420
rect 6166 4386 6200 4388
rect 6360 4490 6394 4492
rect 6360 4458 6394 4490
rect 6360 4388 6394 4420
rect 6360 4386 6394 4388
rect 6518 4490 6552 4492
rect 6518 4458 6552 4490
rect 6518 4388 6552 4420
rect 6518 4386 6552 4388
rect 6668 4490 6702 4492
rect 6668 4458 6702 4490
rect 6668 4388 6702 4420
rect 6668 4386 6702 4388
rect 6826 4490 6860 4492
rect 6826 4458 6860 4490
rect 6826 4388 6860 4420
rect 6826 4386 6860 4388
rect 2857 4237 2891 4271
rect 3670 4261 3704 4295
rect 3984 4252 4018 4286
rect 1410 4123 1444 4157
rect 565 4044 606 4068
rect 712 4044 753 4068
rect 856 4050 897 4073
rect 1568 4123 1602 4157
rect 1698 4123 1732 4157
rect 1856 4123 1890 4157
rect 2030 4123 2064 4157
rect 2188 4123 2222 4157
rect 2372 4123 2406 4157
rect 1010 4050 1051 4074
rect 565 4028 569 4044
rect 569 4028 603 4044
rect 603 4028 606 4044
rect 712 4028 715 4044
rect 715 4028 749 4044
rect 749 4028 753 4044
rect 856 4033 859 4050
rect 859 4033 893 4050
rect 893 4033 897 4050
rect 1010 4034 1013 4050
rect 1013 4034 1047 4050
rect 1047 4034 1051 4050
rect 1373 3946 1387 3980
rect 1387 3946 1407 3980
rect 1445 3946 1455 3980
rect 1455 3946 1479 3980
rect 1517 3946 1523 3980
rect 1523 3946 1551 3980
rect 1589 3946 1591 3980
rect 1591 3946 1623 3980
rect 1661 3946 1693 3980
rect 1693 3946 1695 3980
rect 1733 3946 1761 3980
rect 1761 3946 1767 3980
rect 1805 3946 1829 3980
rect 1829 3946 1839 3980
rect 1877 3946 1897 3980
rect 1897 3946 1911 3980
rect 2530 4123 2564 4157
rect 2369 3921 2403 3955
rect 4306 4246 4340 4280
rect 4637 4264 4671 4298
rect 5628 4262 5662 4296
rect 5942 4252 5976 4286
rect 6264 4246 6298 4280
rect 6596 4264 6630 4298
rect 2776 4123 2810 4157
rect 2934 4123 2968 4157
rect 3120 4123 3154 4157
rect 3278 4123 3312 4157
rect 3742 4133 3776 4167
rect 3900 4133 3934 4167
rect 4050 4133 4084 4167
rect 4208 4133 4242 4167
rect 4402 4135 4436 4169
rect 4560 4135 4594 4169
rect 4710 4135 4744 4169
rect 4868 4135 4902 4169
rect 5700 4134 5734 4168
rect 5858 4134 5892 4168
rect 6008 4134 6042 4168
rect 6166 4134 6200 4168
rect 6360 4136 6394 4170
rect 6518 4136 6552 4170
rect 6668 4136 6702 4170
rect 6826 4136 6860 4170
rect 3741 3957 3753 3991
rect 3753 3957 3775 3991
rect 3813 3957 3821 3991
rect 3821 3957 3847 3991
rect 3885 3957 3889 3991
rect 3889 3957 3919 3991
rect 3957 3957 3991 3991
rect 4029 3957 4059 3991
rect 4059 3957 4063 3991
rect 4101 3957 4127 3991
rect 4127 3957 4135 3991
rect 4173 3957 4195 3991
rect 4195 3957 4207 3991
rect 5700 3958 5712 3992
rect 5712 3958 5734 3992
rect 5772 3958 5780 3992
rect 5780 3958 5806 3992
rect 5844 3958 5848 3992
rect 5848 3958 5878 3992
rect 5916 3958 5950 3992
rect 5988 3958 6018 3992
rect 6018 3958 6022 3992
rect 6060 3958 6086 3992
rect 6086 3958 6094 3992
rect 6132 3958 6154 3992
rect 6154 3958 6166 3992
rect 2642 3805 2696 3859
rect 1383 3420 1395 3454
rect 1395 3420 1417 3454
rect 1455 3420 1463 3454
rect 1463 3420 1489 3454
rect 1527 3420 1531 3454
rect 1531 3420 1561 3454
rect 1599 3420 1633 3454
rect 1671 3420 1701 3454
rect 1701 3420 1705 3454
rect 1743 3420 1769 3454
rect 1769 3420 1777 3454
rect 1815 3420 1837 3454
rect 1837 3420 1849 3454
rect 566 3350 569 3368
rect 569 3350 603 3368
rect 603 3350 607 3368
rect 710 3350 715 3368
rect 715 3350 749 3368
rect 749 3350 751 3368
rect 856 3356 859 3373
rect 859 3356 893 3373
rect 893 3356 897 3373
rect 1009 3356 1013 3373
rect 1013 3356 1047 3373
rect 1047 3356 1050 3373
rect 566 3328 607 3350
rect 710 3328 751 3350
rect 856 3333 897 3356
rect 1009 3333 1050 3356
rect 1410 3251 1444 3253
rect 1410 3219 1444 3251
rect 1410 3149 1444 3181
rect 1410 3147 1444 3149
rect 1568 3251 1602 3253
rect 1568 3219 1602 3251
rect 1568 3149 1602 3181
rect 1568 3147 1602 3149
rect 1698 3251 1732 3253
rect 1698 3219 1732 3251
rect 1698 3149 1732 3181
rect 1698 3147 1732 3149
rect 1856 3251 1890 3253
rect 1856 3219 1890 3251
rect 1856 3149 1890 3181
rect 1856 3147 1890 3149
rect 2030 3251 2064 3253
rect 2030 3219 2064 3251
rect 2030 3149 2064 3181
rect 2030 3147 2064 3149
rect 2188 3251 2222 3253
rect 2188 3219 2222 3251
rect 2188 3149 2222 3181
rect 2188 3147 2222 3149
rect 2372 3251 2406 3253
rect 2372 3219 2406 3251
rect 2372 3149 2406 3181
rect 2372 3147 2406 3149
rect 2530 3251 2564 3253
rect 2530 3219 2564 3251
rect 2776 3251 2810 3253
rect 2530 3149 2564 3181
rect 2530 3147 2564 3149
rect 2647 3167 2681 3201
rect 2776 3219 2810 3251
rect 2776 3149 2810 3181
rect 2776 3147 2810 3149
rect 2934 3251 2968 3253
rect 2934 3219 2968 3251
rect 2934 3149 2968 3181
rect 2934 3147 2968 3149
rect 1269 3013 1303 3047
rect 1773 3013 1807 3047
rect 2273 3011 2307 3045
rect 3797 3419 3807 3453
rect 3807 3419 3831 3453
rect 3869 3419 3875 3453
rect 3875 3419 3903 3453
rect 3941 3419 3943 3453
rect 3943 3419 3975 3453
rect 4013 3419 4045 3453
rect 4045 3419 4047 3453
rect 4085 3419 4113 3453
rect 4113 3419 4119 3453
rect 4157 3419 4181 3453
rect 4181 3419 4191 3453
rect 5756 3418 5766 3452
rect 5766 3418 5790 3452
rect 5828 3418 5834 3452
rect 5834 3418 5862 3452
rect 5900 3418 5902 3452
rect 5902 3418 5934 3452
rect 5972 3418 6004 3452
rect 6004 3418 6006 3452
rect 6044 3418 6072 3452
rect 6072 3418 6078 3452
rect 6116 3418 6140 3452
rect 6140 3418 6150 3452
rect 3120 3251 3154 3253
rect 3120 3219 3154 3251
rect 3120 3149 3154 3181
rect 3120 3147 3154 3149
rect 3278 3251 3312 3253
rect 3278 3219 3312 3251
rect 3278 3149 3312 3181
rect 3278 3147 3312 3149
rect 3742 3261 3776 3263
rect 3742 3229 3776 3261
rect 3742 3159 3776 3191
rect 3742 3157 3776 3159
rect 3900 3261 3934 3263
rect 3900 3229 3934 3261
rect 3900 3159 3934 3191
rect 3900 3157 3934 3159
rect 4050 3261 4084 3263
rect 4050 3229 4084 3261
rect 4050 3159 4084 3191
rect 4050 3157 4084 3159
rect 4208 3261 4242 3263
rect 4208 3229 4242 3261
rect 4208 3159 4242 3191
rect 4208 3157 4242 3159
rect 4402 3261 4436 3263
rect 4402 3229 4436 3261
rect 4402 3159 4436 3191
rect 4402 3157 4436 3159
rect 4560 3261 4594 3263
rect 4560 3229 4594 3261
rect 4560 3159 4594 3191
rect 4560 3157 4594 3159
rect 4710 3261 4744 3263
rect 4710 3229 4744 3261
rect 4710 3159 4744 3191
rect 4710 3157 4744 3159
rect 4868 3261 4902 3263
rect 4868 3229 4902 3261
rect 4868 3159 4902 3191
rect 4868 3157 4902 3159
rect 5700 3262 5734 3264
rect 5700 3230 5734 3262
rect 5700 3160 5734 3192
rect 5700 3158 5734 3160
rect 5858 3262 5892 3264
rect 5858 3230 5892 3262
rect 5858 3160 5892 3192
rect 5858 3158 5892 3160
rect 6008 3262 6042 3264
rect 6008 3230 6042 3262
rect 6008 3160 6042 3192
rect 6008 3158 6042 3160
rect 6166 3262 6200 3264
rect 6166 3230 6200 3262
rect 6166 3160 6200 3192
rect 6166 3158 6200 3160
rect 6360 3262 6394 3264
rect 6360 3230 6394 3262
rect 6360 3160 6394 3192
rect 6360 3158 6394 3160
rect 6518 3262 6552 3264
rect 6518 3230 6552 3262
rect 6518 3160 6552 3192
rect 6518 3158 6552 3160
rect 6668 3262 6702 3264
rect 6668 3230 6702 3262
rect 6668 3160 6702 3192
rect 6668 3158 6702 3160
rect 6826 3262 6860 3264
rect 6826 3230 6860 3262
rect 6826 3160 6860 3192
rect 6826 3158 6860 3160
rect 2857 3009 2891 3043
rect 3670 3033 3704 3067
rect 3984 3024 4018 3058
rect 1410 2895 1444 2929
rect 565 2816 606 2840
rect 712 2816 753 2840
rect 856 2822 897 2845
rect 1568 2895 1602 2929
rect 1698 2895 1732 2929
rect 1856 2895 1890 2929
rect 2030 2895 2064 2929
rect 2188 2895 2222 2929
rect 2372 2895 2406 2929
rect 1010 2822 1051 2846
rect 565 2800 569 2816
rect 569 2800 603 2816
rect 603 2800 606 2816
rect 712 2800 715 2816
rect 715 2800 749 2816
rect 749 2800 753 2816
rect 856 2805 859 2822
rect 859 2805 893 2822
rect 893 2805 897 2822
rect 1010 2806 1013 2822
rect 1013 2806 1047 2822
rect 1047 2806 1051 2822
rect 1373 2718 1387 2752
rect 1387 2718 1407 2752
rect 1445 2718 1455 2752
rect 1455 2718 1479 2752
rect 1517 2718 1523 2752
rect 1523 2718 1551 2752
rect 1589 2718 1591 2752
rect 1591 2718 1623 2752
rect 1661 2718 1693 2752
rect 1693 2718 1695 2752
rect 1733 2718 1761 2752
rect 1761 2718 1767 2752
rect 1805 2718 1829 2752
rect 1829 2718 1839 2752
rect 1877 2718 1897 2752
rect 1897 2718 1911 2752
rect 2530 2895 2564 2929
rect 2369 2693 2403 2727
rect 4306 3018 4340 3052
rect 4637 3036 4671 3070
rect 5628 3034 5662 3068
rect 5942 3024 5976 3058
rect 6264 3018 6298 3052
rect 6596 3036 6630 3070
rect 2776 2895 2810 2929
rect 2934 2895 2968 2929
rect 3120 2895 3154 2929
rect 3278 2895 3312 2929
rect 3742 2905 3776 2939
rect 3900 2905 3934 2939
rect 4050 2905 4084 2939
rect 4208 2905 4242 2939
rect 4402 2907 4436 2941
rect 4560 2907 4594 2941
rect 4710 2907 4744 2941
rect 4868 2907 4902 2941
rect 5700 2906 5734 2940
rect 5858 2906 5892 2940
rect 6008 2906 6042 2940
rect 6166 2906 6200 2940
rect 6360 2908 6394 2942
rect 6518 2908 6552 2942
rect 6668 2908 6702 2942
rect 6826 2908 6860 2942
rect 3741 2729 3753 2763
rect 3753 2729 3775 2763
rect 3813 2729 3821 2763
rect 3821 2729 3847 2763
rect 3885 2729 3889 2763
rect 3889 2729 3919 2763
rect 3957 2729 3991 2763
rect 4029 2729 4059 2763
rect 4059 2729 4063 2763
rect 4101 2729 4127 2763
rect 4127 2729 4135 2763
rect 4173 2729 4195 2763
rect 4195 2729 4207 2763
rect 5700 2730 5712 2764
rect 5712 2730 5734 2764
rect 5772 2730 5780 2764
rect 5780 2730 5806 2764
rect 5844 2730 5848 2764
rect 5848 2730 5878 2764
rect 5916 2730 5950 2764
rect 5988 2730 6018 2764
rect 6018 2730 6022 2764
rect 6060 2730 6086 2764
rect 6086 2730 6094 2764
rect 6132 2730 6154 2764
rect 6154 2730 6166 2764
rect 2642 2577 2696 2631
rect 1383 2192 1395 2226
rect 1395 2192 1417 2226
rect 1455 2192 1463 2226
rect 1463 2192 1489 2226
rect 1527 2192 1531 2226
rect 1531 2192 1561 2226
rect 1599 2192 1633 2226
rect 1671 2192 1701 2226
rect 1701 2192 1705 2226
rect 1743 2192 1769 2226
rect 1769 2192 1777 2226
rect 1815 2192 1837 2226
rect 1837 2192 1849 2226
rect 566 2122 569 2140
rect 569 2122 603 2140
rect 603 2122 607 2140
rect 710 2122 715 2140
rect 715 2122 749 2140
rect 749 2122 751 2140
rect 856 2128 859 2145
rect 859 2128 893 2145
rect 893 2128 897 2145
rect 1009 2128 1013 2145
rect 1013 2128 1047 2145
rect 1047 2128 1050 2145
rect 566 2100 607 2122
rect 710 2100 751 2122
rect 856 2105 897 2128
rect 1009 2105 1050 2128
rect 1410 2023 1444 2025
rect 1410 1991 1444 2023
rect 1410 1921 1444 1953
rect 1410 1919 1444 1921
rect 1568 2023 1602 2025
rect 1568 1991 1602 2023
rect 1568 1921 1602 1953
rect 1568 1919 1602 1921
rect 1698 2023 1732 2025
rect 1698 1991 1732 2023
rect 1698 1921 1732 1953
rect 1698 1919 1732 1921
rect 1856 2023 1890 2025
rect 1856 1991 1890 2023
rect 1856 1921 1890 1953
rect 1856 1919 1890 1921
rect 2030 2023 2064 2025
rect 2030 1991 2064 2023
rect 2030 1921 2064 1953
rect 2030 1919 2064 1921
rect 2188 2023 2222 2025
rect 2188 1991 2222 2023
rect 2188 1921 2222 1953
rect 2188 1919 2222 1921
rect 2372 2023 2406 2025
rect 2372 1991 2406 2023
rect 2372 1921 2406 1953
rect 2372 1919 2406 1921
rect 2530 2023 2564 2025
rect 2530 1991 2564 2023
rect 2776 2023 2810 2025
rect 2530 1921 2564 1953
rect 2530 1919 2564 1921
rect 2647 1939 2681 1973
rect 2776 1991 2810 2023
rect 2776 1921 2810 1953
rect 2776 1919 2810 1921
rect 2934 2023 2968 2025
rect 2934 1991 2968 2023
rect 2934 1921 2968 1953
rect 2934 1919 2968 1921
rect 1269 1785 1303 1819
rect 1773 1785 1807 1819
rect 2273 1783 2307 1817
rect 3797 2191 3807 2225
rect 3807 2191 3831 2225
rect 3869 2191 3875 2225
rect 3875 2191 3903 2225
rect 3941 2191 3943 2225
rect 3943 2191 3975 2225
rect 4013 2191 4045 2225
rect 4045 2191 4047 2225
rect 4085 2191 4113 2225
rect 4113 2191 4119 2225
rect 4157 2191 4181 2225
rect 4181 2191 4191 2225
rect 5756 2190 5766 2224
rect 5766 2190 5790 2224
rect 5828 2190 5834 2224
rect 5834 2190 5862 2224
rect 5900 2190 5902 2224
rect 5902 2190 5934 2224
rect 5972 2190 6004 2224
rect 6004 2190 6006 2224
rect 6044 2190 6072 2224
rect 6072 2190 6078 2224
rect 6116 2190 6140 2224
rect 6140 2190 6150 2224
rect 3120 2023 3154 2025
rect 3120 1991 3154 2023
rect 3120 1921 3154 1953
rect 3120 1919 3154 1921
rect 3278 2023 3312 2025
rect 3278 1991 3312 2023
rect 3278 1921 3312 1953
rect 3278 1919 3312 1921
rect 3742 2033 3776 2035
rect 3742 2001 3776 2033
rect 3742 1931 3776 1963
rect 3742 1929 3776 1931
rect 3900 2033 3934 2035
rect 3900 2001 3934 2033
rect 3900 1931 3934 1963
rect 3900 1929 3934 1931
rect 4050 2033 4084 2035
rect 4050 2001 4084 2033
rect 4050 1931 4084 1963
rect 4050 1929 4084 1931
rect 4208 2033 4242 2035
rect 4208 2001 4242 2033
rect 4208 1931 4242 1963
rect 4208 1929 4242 1931
rect 4402 2033 4436 2035
rect 4402 2001 4436 2033
rect 4402 1931 4436 1963
rect 4402 1929 4436 1931
rect 4560 2033 4594 2035
rect 4560 2001 4594 2033
rect 4560 1931 4594 1963
rect 4560 1929 4594 1931
rect 4710 2033 4744 2035
rect 4710 2001 4744 2033
rect 4710 1931 4744 1963
rect 4710 1929 4744 1931
rect 4868 2033 4902 2035
rect 4868 2001 4902 2033
rect 4868 1931 4902 1963
rect 4868 1929 4902 1931
rect 5700 2034 5734 2036
rect 5700 2002 5734 2034
rect 5700 1932 5734 1964
rect 5700 1930 5734 1932
rect 5858 2034 5892 2036
rect 5858 2002 5892 2034
rect 5858 1932 5892 1964
rect 5858 1930 5892 1932
rect 6008 2034 6042 2036
rect 6008 2002 6042 2034
rect 6008 1932 6042 1964
rect 6008 1930 6042 1932
rect 6166 2034 6200 2036
rect 6166 2002 6200 2034
rect 6166 1932 6200 1964
rect 6166 1930 6200 1932
rect 6360 2034 6394 2036
rect 6360 2002 6394 2034
rect 6360 1932 6394 1964
rect 6360 1930 6394 1932
rect 6518 2034 6552 2036
rect 6518 2002 6552 2034
rect 6518 1932 6552 1964
rect 6518 1930 6552 1932
rect 6668 2034 6702 2036
rect 6668 2002 6702 2034
rect 6668 1932 6702 1964
rect 6668 1930 6702 1932
rect 6826 2034 6860 2036
rect 6826 2002 6860 2034
rect 6826 1932 6860 1964
rect 6826 1930 6860 1932
rect 2857 1781 2891 1815
rect 3670 1805 3704 1839
rect 3984 1796 4018 1830
rect 1410 1667 1444 1701
rect 565 1588 606 1612
rect 712 1588 753 1612
rect 856 1594 897 1617
rect 1568 1667 1602 1701
rect 1698 1667 1732 1701
rect 1856 1667 1890 1701
rect 2030 1667 2064 1701
rect 2188 1667 2222 1701
rect 2372 1667 2406 1701
rect 1010 1594 1051 1618
rect 565 1572 569 1588
rect 569 1572 603 1588
rect 603 1572 606 1588
rect 712 1572 715 1588
rect 715 1572 749 1588
rect 749 1572 753 1588
rect 856 1577 859 1594
rect 859 1577 893 1594
rect 893 1577 897 1594
rect 1010 1578 1013 1594
rect 1013 1578 1047 1594
rect 1047 1578 1051 1594
rect 1373 1490 1387 1524
rect 1387 1490 1407 1524
rect 1445 1490 1455 1524
rect 1455 1490 1479 1524
rect 1517 1490 1523 1524
rect 1523 1490 1551 1524
rect 1589 1490 1591 1524
rect 1591 1490 1623 1524
rect 1661 1490 1693 1524
rect 1693 1490 1695 1524
rect 1733 1490 1761 1524
rect 1761 1490 1767 1524
rect 1805 1490 1829 1524
rect 1829 1490 1839 1524
rect 1877 1490 1897 1524
rect 1897 1490 1911 1524
rect 2530 1667 2564 1701
rect 2369 1465 2403 1499
rect 4306 1790 4340 1824
rect 4637 1808 4671 1842
rect 5628 1806 5662 1840
rect 5942 1796 5976 1830
rect 6264 1790 6298 1824
rect 6596 1808 6630 1842
rect 2776 1667 2810 1701
rect 2934 1667 2968 1701
rect 3120 1667 3154 1701
rect 3278 1667 3312 1701
rect 3742 1677 3776 1711
rect 3900 1677 3934 1711
rect 4050 1677 4084 1711
rect 4208 1677 4242 1711
rect 4402 1679 4436 1713
rect 4560 1679 4594 1713
rect 4710 1679 4744 1713
rect 4868 1679 4902 1713
rect 5700 1678 5734 1712
rect 5858 1678 5892 1712
rect 6008 1678 6042 1712
rect 6166 1678 6200 1712
rect 6360 1680 6394 1714
rect 6518 1680 6552 1714
rect 6668 1680 6702 1714
rect 6826 1680 6860 1714
rect 3741 1501 3753 1535
rect 3753 1501 3775 1535
rect 3813 1501 3821 1535
rect 3821 1501 3847 1535
rect 3885 1501 3889 1535
rect 3889 1501 3919 1535
rect 3957 1501 3991 1535
rect 4029 1501 4059 1535
rect 4059 1501 4063 1535
rect 4101 1501 4127 1535
rect 4127 1501 4135 1535
rect 4173 1501 4195 1535
rect 4195 1501 4207 1535
rect 5700 1502 5712 1536
rect 5712 1502 5734 1536
rect 5772 1502 5780 1536
rect 5780 1502 5806 1536
rect 5844 1502 5848 1536
rect 5848 1502 5878 1536
rect 5916 1502 5950 1536
rect 5988 1502 6018 1536
rect 6018 1502 6022 1536
rect 6060 1502 6086 1536
rect 6086 1502 6094 1536
rect 6132 1502 6154 1536
rect 6154 1502 6166 1536
rect 2642 1349 2696 1403
rect 1383 964 1395 998
rect 1395 964 1417 998
rect 1455 964 1463 998
rect 1463 964 1489 998
rect 1527 964 1531 998
rect 1531 964 1561 998
rect 1599 964 1633 998
rect 1671 964 1701 998
rect 1701 964 1705 998
rect 1743 964 1769 998
rect 1769 964 1777 998
rect 1815 964 1837 998
rect 1837 964 1849 998
rect 566 894 569 912
rect 569 894 603 912
rect 603 894 607 912
rect 710 894 715 912
rect 715 894 749 912
rect 749 894 751 912
rect 856 900 859 917
rect 859 900 893 917
rect 893 900 897 917
rect 1009 900 1013 917
rect 1013 900 1047 917
rect 1047 900 1050 917
rect 566 872 607 894
rect 710 872 751 894
rect 856 877 897 900
rect 1009 877 1050 900
rect 1410 795 1444 797
rect 1410 763 1444 795
rect 1410 693 1444 725
rect 1410 691 1444 693
rect 1568 795 1602 797
rect 1568 763 1602 795
rect 1568 693 1602 725
rect 1568 691 1602 693
rect 1698 795 1732 797
rect 1698 763 1732 795
rect 1698 693 1732 725
rect 1698 691 1732 693
rect 1856 795 1890 797
rect 1856 763 1890 795
rect 1856 693 1890 725
rect 1856 691 1890 693
rect 2030 795 2064 797
rect 2030 763 2064 795
rect 2030 693 2064 725
rect 2030 691 2064 693
rect 2188 795 2222 797
rect 2188 763 2222 795
rect 2188 693 2222 725
rect 2188 691 2222 693
rect 2372 795 2406 797
rect 2372 763 2406 795
rect 2372 693 2406 725
rect 2372 691 2406 693
rect 2530 795 2564 797
rect 2530 763 2564 795
rect 2776 795 2810 797
rect 2530 693 2564 725
rect 2530 691 2564 693
rect 2647 711 2681 745
rect 2776 763 2810 795
rect 2776 693 2810 725
rect 2776 691 2810 693
rect 2934 795 2968 797
rect 2934 763 2968 795
rect 2934 693 2968 725
rect 2934 691 2968 693
rect 1269 557 1303 591
rect 1773 557 1807 591
rect 2273 555 2307 589
rect 3797 963 3807 997
rect 3807 963 3831 997
rect 3869 963 3875 997
rect 3875 963 3903 997
rect 3941 963 3943 997
rect 3943 963 3975 997
rect 4013 963 4045 997
rect 4045 963 4047 997
rect 4085 963 4113 997
rect 4113 963 4119 997
rect 4157 963 4181 997
rect 4181 963 4191 997
rect 3120 795 3154 797
rect 3120 763 3154 795
rect 3120 693 3154 725
rect 3120 691 3154 693
rect 3278 795 3312 797
rect 3278 763 3312 795
rect 3278 693 3312 725
rect 3278 691 3312 693
rect 3742 805 3776 807
rect 3742 773 3776 805
rect 3742 703 3776 735
rect 3742 701 3776 703
rect 3900 805 3934 807
rect 3900 773 3934 805
rect 3900 703 3934 735
rect 3900 701 3934 703
rect 4050 805 4084 807
rect 4050 773 4084 805
rect 4050 703 4084 735
rect 4050 701 4084 703
rect 4208 805 4242 807
rect 4208 773 4242 805
rect 4208 703 4242 735
rect 4208 701 4242 703
rect 4402 805 4436 807
rect 4402 773 4436 805
rect 4402 703 4436 735
rect 4402 701 4436 703
rect 4560 805 4594 807
rect 4560 773 4594 805
rect 4560 703 4594 735
rect 4560 701 4594 703
rect 4710 805 4744 807
rect 4710 773 4744 805
rect 4710 703 4744 735
rect 4710 701 4744 703
rect 4868 805 4902 807
rect 4868 773 4902 805
rect 4868 703 4902 735
rect 4868 701 4902 703
rect 2857 553 2891 587
rect 3670 577 3704 611
rect 3984 568 4018 602
rect 1410 439 1444 473
rect 565 360 606 384
rect 712 360 753 384
rect 856 366 897 389
rect 1568 439 1602 473
rect 1698 439 1732 473
rect 1856 439 1890 473
rect 2030 439 2064 473
rect 2188 439 2222 473
rect 2372 439 2406 473
rect 1010 366 1051 390
rect 565 344 569 360
rect 569 344 603 360
rect 603 344 606 360
rect 712 344 715 360
rect 715 344 749 360
rect 749 344 753 360
rect 856 349 859 366
rect 859 349 893 366
rect 893 349 897 366
rect 1010 350 1013 366
rect 1013 350 1047 366
rect 1047 350 1051 366
rect 1373 262 1387 296
rect 1387 262 1407 296
rect 1445 262 1455 296
rect 1455 262 1479 296
rect 1517 262 1523 296
rect 1523 262 1551 296
rect 1589 262 1591 296
rect 1591 262 1623 296
rect 1661 262 1693 296
rect 1693 262 1695 296
rect 1733 262 1761 296
rect 1761 262 1767 296
rect 1805 262 1829 296
rect 1829 262 1839 296
rect 1877 262 1897 296
rect 1897 262 1911 296
rect 2530 439 2564 473
rect 2369 237 2403 271
rect 4306 562 4340 596
rect 4637 580 4671 614
rect 2776 439 2810 473
rect 2934 439 2968 473
rect 3120 439 3154 473
rect 3278 439 3312 473
rect 3742 449 3776 483
rect 3900 449 3934 483
rect 4050 449 4084 483
rect 4208 449 4242 483
rect 4402 451 4436 485
rect 4560 451 4594 485
rect 4710 451 4744 485
rect 4868 451 4902 485
rect 3741 273 3753 307
rect 3753 273 3775 307
rect 3813 273 3821 307
rect 3821 273 3847 307
rect 3885 273 3889 307
rect 3889 273 3919 307
rect 3957 273 3991 307
rect 4029 273 4059 307
rect 4059 273 4063 307
rect 4101 273 4127 307
rect 4127 273 4135 307
rect 4173 273 4195 307
rect 4195 273 4207 307
rect 2642 121 2696 175
<< metal1 >>
rect 5029 19608 5081 19614
rect 3472 19561 4907 19600
rect 1348 19427 1880 19470
rect 1348 19418 1398 19427
rect 1450 19418 1462 19427
rect 1348 19384 1383 19418
rect 1450 19384 1455 19418
rect 1348 19375 1398 19384
rect 1450 19375 1462 19384
rect 1514 19375 1526 19427
rect 1578 19375 1590 19427
rect 1642 19375 1654 19427
rect 1706 19375 1718 19427
rect 1770 19418 1782 19427
rect 1834 19418 1880 19427
rect 1777 19384 1782 19418
rect 1849 19384 1880 19418
rect 3472 19403 3511 19561
rect 4738 19519 4744 19526
rect 4558 19480 4744 19519
rect 1770 19375 1782 19384
rect 1834 19375 1880 19384
rect 550 19356 622 19360
rect 550 19304 560 19356
rect 612 19304 622 19356
rect 696 19354 768 19360
rect 550 19292 566 19304
rect 607 19292 622 19304
rect 682 19352 768 19354
rect 682 19300 702 19352
rect 754 19300 768 19352
rect 682 19298 710 19300
rect 550 19262 622 19292
rect 696 19292 710 19298
rect 751 19292 768 19300
rect 696 19262 768 19292
rect 840 19337 912 19366
rect 840 19297 856 19337
rect 897 19297 912 19337
rect 840 19268 912 19297
rect 994 19337 1066 19366
rect 994 19297 1009 19337
rect 1050 19297 1066 19337
rect 1348 19330 1880 19375
rect 994 19268 1066 19297
rect 564 19222 608 19262
rect 856 19202 900 19268
rect 378 19194 433 19200
rect 846 19150 852 19202
rect 904 19150 910 19202
rect 378 18909 433 19139
rect 856 19110 900 19150
rect 1008 19110 1052 19268
rect 1407 19264 1448 19330
rect 1693 19264 1735 19330
rect 1941 19327 2687 19372
rect 1404 19217 1450 19264
rect 1404 19183 1410 19217
rect 1444 19183 1450 19217
rect 1404 19145 1450 19183
rect 1404 19111 1410 19145
rect 1444 19111 1450 19145
rect 708 19066 900 19110
rect 372 18854 378 18909
rect 433 18854 439 18909
rect 708 18832 752 19066
rect 998 19058 1004 19110
rect 1056 19058 1062 19110
rect 1404 19064 1450 19111
rect 1562 19217 1608 19264
rect 1562 19183 1568 19217
rect 1602 19183 1608 19217
rect 1562 19145 1608 19183
rect 1562 19111 1568 19145
rect 1602 19111 1608 19145
rect 1562 19064 1608 19111
rect 1692 19217 1738 19264
rect 1692 19183 1698 19217
rect 1732 19183 1738 19217
rect 1692 19145 1738 19183
rect 1692 19111 1698 19145
rect 1732 19111 1738 19145
rect 1692 19064 1738 19111
rect 1850 19261 1896 19264
rect 1941 19261 1986 19327
rect 1850 19217 1986 19261
rect 1850 19183 1856 19217
rect 1890 19216 1986 19217
rect 2024 19217 2070 19264
rect 1890 19183 1896 19216
rect 1850 19145 1896 19183
rect 2024 19183 2030 19217
rect 2064 19183 2070 19217
rect 2024 19148 2070 19183
rect 1998 19146 2070 19148
rect 1850 19111 1856 19145
rect 1890 19111 1896 19145
rect 1850 19064 1896 19111
rect 1928 19145 2070 19146
rect 1928 19121 2030 19145
rect 1928 19104 1935 19121
rect 1929 19069 1935 19104
rect 1987 19111 2030 19121
rect 2064 19111 2070 19145
rect 1987 19104 2070 19111
rect 1987 19069 1993 19104
rect 2024 19064 2070 19104
rect 2182 19220 2228 19264
rect 2366 19220 2412 19264
rect 2182 19217 2412 19220
rect 2182 19183 2188 19217
rect 2222 19183 2372 19217
rect 2406 19183 2412 19217
rect 2182 19145 2412 19183
rect 2182 19111 2188 19145
rect 2222 19111 2372 19145
rect 2406 19111 2412 19145
rect 2182 19094 2412 19111
rect 2182 19064 2228 19094
rect 2366 19064 2412 19094
rect 2524 19217 2570 19264
rect 2524 19183 2530 19217
rect 2564 19183 2570 19217
rect 2642 19193 2687 19327
rect 3118 19364 3511 19403
rect 3724 19426 4264 19470
rect 3724 19374 3776 19426
rect 3828 19417 3840 19426
rect 3892 19417 3904 19426
rect 3956 19417 3968 19426
rect 4020 19417 4032 19426
rect 4084 19417 4096 19426
rect 4148 19417 4160 19426
rect 3831 19383 3840 19417
rect 3903 19383 3904 19417
rect 4084 19383 4085 19417
rect 4148 19383 4157 19417
rect 3828 19374 3840 19383
rect 3892 19374 3904 19383
rect 3956 19374 3968 19383
rect 4020 19374 4032 19383
rect 4084 19374 4096 19383
rect 4148 19374 4160 19383
rect 4212 19374 4264 19426
rect 2774 19320 2816 19321
rect 2758 19312 2816 19320
rect 2758 19260 2769 19312
rect 2821 19260 2827 19312
rect 3118 19264 3157 19364
rect 3724 19330 4264 19374
rect 3741 19274 3787 19330
rect 3736 19273 3787 19274
rect 2758 19217 2816 19260
rect 2524 19145 2570 19183
rect 2524 19111 2530 19145
rect 2564 19111 2570 19145
rect 2524 19104 2570 19111
rect 2613 19165 2715 19193
rect 2613 19131 2647 19165
rect 2681 19131 2715 19165
rect 2524 19064 2574 19104
rect 2613 19103 2715 19131
rect 2758 19183 2776 19217
rect 2810 19183 2816 19217
rect 2758 19145 2816 19183
rect 2758 19111 2776 19145
rect 2810 19111 2816 19145
rect 1008 19004 1052 19058
rect 1245 19023 1328 19042
rect 852 18960 1052 19004
rect 1148 19021 1328 19023
rect 1148 18969 1155 19021
rect 1207 19011 1328 19021
rect 1207 18977 1269 19011
rect 1303 18977 1328 19011
rect 1207 18969 1328 18977
rect 1148 18968 1328 18969
rect 852 18838 896 18960
rect 1245 18947 1328 18968
rect 1568 19030 1602 19064
rect 1568 19020 1820 19030
rect 1568 18968 1758 19020
rect 1810 18968 1820 19020
rect 1568 18958 1820 18968
rect 1568 18926 1608 18958
rect 1853 18926 1892 19064
rect 2185 18926 2224 19064
rect 2255 19027 2325 19033
rect 2255 19018 2331 19027
rect 2255 18966 2270 19018
rect 2322 18966 2331 19018
rect 2255 18957 2331 18966
rect 2255 18951 2325 18957
rect 2368 18926 2407 19064
rect 2530 19030 2574 19064
rect 2758 19064 2816 19111
rect 2928 19217 2974 19264
rect 2928 19183 2934 19217
rect 2968 19204 2974 19217
rect 3114 19217 3160 19264
rect 3114 19204 3120 19217
rect 2968 19183 3120 19204
rect 3154 19183 3160 19217
rect 3272 19217 3318 19264
rect 3272 19207 3278 19217
rect 3312 19207 3318 19217
rect 3736 19227 3782 19273
rect 2928 19145 3160 19183
rect 3262 19155 3268 19207
rect 3320 19155 3326 19207
rect 3736 19193 3742 19227
rect 3776 19193 3782 19227
rect 3736 19155 3782 19193
rect 2928 19111 2934 19145
rect 2968 19111 3120 19145
rect 3154 19111 3160 19145
rect 2928 19094 3160 19111
rect 2928 19064 2974 19094
rect 3114 19064 3160 19094
rect 3272 19145 3318 19155
rect 3272 19111 3278 19145
rect 3312 19111 3318 19145
rect 3272 19064 3318 19111
rect 3736 19121 3742 19155
rect 3776 19121 3782 19155
rect 3736 19074 3782 19121
rect 3894 19227 3940 19274
rect 3894 19193 3900 19227
rect 3934 19193 3940 19227
rect 3894 19155 3940 19193
rect 3894 19121 3900 19155
rect 3934 19121 3940 19155
rect 3894 19074 3940 19121
rect 4044 19227 4090 19330
rect 4558 19274 4597 19480
rect 4738 19474 4744 19480
rect 4796 19474 4802 19526
rect 4868 19274 4907 19561
rect 5081 19567 7015 19597
rect 5029 19550 5081 19556
rect 6862 19519 6868 19526
rect 6516 19480 6868 19519
rect 5682 19426 6222 19470
rect 5682 19374 5734 19426
rect 5786 19416 5798 19426
rect 5850 19416 5862 19426
rect 5914 19416 5926 19426
rect 5978 19416 5990 19426
rect 6042 19416 6054 19426
rect 6106 19416 6118 19426
rect 5790 19382 5798 19416
rect 6042 19382 6044 19416
rect 6106 19382 6116 19416
rect 5786 19374 5798 19382
rect 5850 19374 5862 19382
rect 5914 19374 5926 19382
rect 5978 19374 5990 19382
rect 6042 19374 6054 19382
rect 6106 19374 6118 19382
rect 6170 19374 6222 19426
rect 5682 19330 6222 19374
rect 5700 19274 5746 19330
rect 4044 19193 4050 19227
rect 4084 19193 4090 19227
rect 4044 19155 4090 19193
rect 4044 19121 4050 19155
rect 4084 19121 4090 19155
rect 4044 19074 4090 19121
rect 4202 19227 4248 19274
rect 4202 19193 4208 19227
rect 4242 19193 4248 19227
rect 4396 19227 4442 19274
rect 4396 19201 4402 19227
rect 4202 19155 4248 19193
rect 4202 19121 4208 19155
rect 4242 19121 4248 19155
rect 4285 19199 4402 19201
rect 4285 19147 4292 19199
rect 4344 19193 4402 19199
rect 4436 19193 4442 19227
rect 4344 19155 4442 19193
rect 4344 19147 4402 19155
rect 4285 19146 4402 19147
rect 4202 19074 4248 19121
rect 4396 19121 4402 19146
rect 4436 19121 4442 19155
rect 4396 19074 4442 19121
rect 4554 19227 4600 19274
rect 4554 19193 4560 19227
rect 4594 19194 4600 19227
rect 4704 19227 4750 19274
rect 4704 19194 4710 19227
rect 4594 19193 4710 19194
rect 4744 19193 4750 19227
rect 4554 19155 4750 19193
rect 4554 19121 4560 19155
rect 4594 19128 4710 19155
rect 4594 19121 4600 19128
rect 4554 19074 4600 19121
rect 4704 19121 4710 19128
rect 4744 19121 4750 19155
rect 4704 19074 4750 19121
rect 4862 19227 4908 19274
rect 4862 19193 4868 19227
rect 4902 19193 4908 19227
rect 5694 19228 5740 19274
rect 5027 19198 5057 19207
rect 4862 19155 4908 19193
rect 4862 19121 4868 19155
rect 4902 19121 4908 19155
rect 5010 19146 5016 19198
rect 5068 19146 5074 19198
rect 5694 19194 5700 19228
rect 5734 19194 5740 19228
rect 5694 19156 5740 19194
rect 4862 19074 4908 19121
rect 5026 19105 5057 19146
rect 5694 19122 5700 19156
rect 5734 19122 5740 19156
rect 2758 19030 2802 19064
rect 2530 18986 2656 19030
rect 1242 18906 1248 18910
rect 1138 18862 1248 18906
rect 1138 18838 1182 18862
rect 1242 18858 1248 18862
rect 1300 18858 1306 18910
rect 1404 18893 1450 18926
rect 1404 18859 1410 18893
rect 1444 18859 1450 18893
rect 1404 18855 1450 18859
rect 378 18810 434 18816
rect 550 18810 622 18832
rect 434 18804 622 18810
rect 434 18764 565 18804
rect 606 18764 622 18804
rect 434 18754 622 18764
rect 378 18748 434 18754
rect 550 18734 622 18754
rect 696 18804 768 18832
rect 696 18764 712 18804
rect 753 18764 768 18804
rect 696 18734 768 18764
rect 840 18809 912 18838
rect 840 18769 856 18809
rect 897 18769 912 18809
rect 840 18740 912 18769
rect 994 18810 1182 18838
rect 994 18770 1010 18810
rect 1051 18794 1182 18810
rect 1399 18826 1450 18855
rect 1562 18893 1608 18926
rect 1562 18859 1568 18893
rect 1602 18859 1608 18893
rect 1692 18893 1738 18926
rect 1692 18864 1698 18893
rect 1562 18826 1608 18859
rect 1690 18859 1698 18864
rect 1732 18864 1738 18893
rect 1850 18893 1896 18926
rect 2024 18910 2070 18926
rect 1732 18859 1740 18864
rect 1051 18770 1066 18794
rect 1399 18780 1449 18826
rect 1690 18780 1740 18859
rect 1850 18859 1856 18893
rect 1890 18859 1896 18893
rect 1850 18826 1896 18859
rect 2014 18858 2020 18910
rect 2072 18858 2078 18910
rect 2182 18893 2228 18926
rect 2182 18859 2188 18893
rect 2222 18859 2228 18893
rect 2024 18826 2070 18858
rect 2182 18826 2228 18859
rect 2366 18893 2412 18926
rect 2524 18908 2570 18926
rect 2366 18859 2372 18893
rect 2406 18859 2412 18893
rect 2366 18826 2412 18859
rect 2516 18856 2522 18908
rect 2574 18856 2580 18908
rect 2524 18826 2570 18856
rect 2024 18794 2068 18826
rect 2612 18794 2656 18986
rect 994 18740 1066 18770
rect 1324 18725 1960 18780
rect 2024 18750 2656 18794
rect 2694 18986 2802 19030
rect 2832 19016 2904 19026
rect 2694 18788 2738 18986
rect 2832 18964 2842 19016
rect 2894 18964 2904 19016
rect 2832 18954 2904 18964
rect 2933 18926 2972 19064
rect 3118 18926 3157 19064
rect 3272 19020 3316 19064
rect 3268 19014 3320 19020
rect 3555 18989 3561 19041
rect 3613 19034 3619 19041
rect 3662 19034 3713 19046
rect 3613 19031 3713 19034
rect 3613 18997 3670 19031
rect 3704 18997 3713 19031
rect 3613 18995 3713 18997
rect 3613 18989 3619 18995
rect 3662 18983 3713 18995
rect 3897 19025 3936 19074
rect 3976 19032 4027 19037
rect 3970 19025 3976 19032
rect 3897 18986 3976 19025
rect 3268 18956 3320 18962
rect 3897 18936 3936 18986
rect 3970 18980 3976 18986
rect 4028 18980 4034 19032
rect 4206 19018 4245 19074
rect 4300 19018 4347 19029
rect 4206 19016 4347 19018
rect 4206 18983 4306 19016
rect 3976 18974 4027 18980
rect 4206 18936 4245 18983
rect 4300 18982 4306 18983
rect 4340 18982 4347 19016
rect 4300 18970 4347 18982
rect 2766 18920 2818 18926
rect 2766 18862 2776 18868
rect 2770 18859 2776 18862
rect 2810 18862 2818 18868
rect 2928 18893 2974 18926
rect 2810 18859 2816 18862
rect 2770 18826 2816 18859
rect 2928 18859 2934 18893
rect 2968 18859 2974 18893
rect 2928 18826 2974 18859
rect 3114 18893 3160 18926
rect 3114 18859 3120 18893
rect 3154 18859 3160 18893
rect 3114 18826 3160 18859
rect 3272 18893 3318 18926
rect 3272 18859 3278 18893
rect 3312 18859 3318 18893
rect 3272 18826 3318 18859
rect 3274 18788 3318 18826
rect 2694 18744 3318 18788
rect 3736 18903 3782 18936
rect 3736 18869 3742 18903
rect 3776 18869 3782 18903
rect 3736 18836 3782 18869
rect 3894 18903 3940 18936
rect 3894 18869 3900 18903
rect 3934 18869 3940 18903
rect 4044 18903 4090 18936
rect 4044 18874 4050 18903
rect 3894 18836 3940 18869
rect 4042 18869 4050 18874
rect 4084 18869 4090 18903
rect 4042 18836 4090 18869
rect 4202 18903 4248 18936
rect 4202 18869 4208 18903
rect 4242 18869 4248 18903
rect 4202 18836 4248 18869
rect 3736 18780 3780 18836
rect 4042 18780 4089 18836
rect 1324 18673 1360 18725
rect 1412 18673 1424 18725
rect 1476 18716 1488 18725
rect 1540 18716 1552 18725
rect 1604 18716 1616 18725
rect 1668 18716 1680 18725
rect 1732 18716 1744 18725
rect 1796 18716 1808 18725
rect 1479 18682 1488 18716
rect 1551 18682 1552 18716
rect 1732 18682 1733 18716
rect 1796 18682 1805 18716
rect 1476 18673 1488 18682
rect 1540 18673 1552 18682
rect 1604 18673 1616 18682
rect 1668 18673 1680 18682
rect 1732 18673 1744 18682
rect 1796 18673 1808 18682
rect 1860 18673 1872 18725
rect 1924 18673 1960 18725
rect 3704 18736 4244 18780
rect 3704 18727 3756 18736
rect 3808 18727 3820 18736
rect 1324 18640 1960 18673
rect 2346 18695 2426 18720
rect 2346 18691 3517 18695
rect 2346 18657 2369 18691
rect 2403 18657 3517 18691
rect 2346 18653 3517 18657
rect 2346 18628 2426 18653
rect 2636 18595 2702 18607
rect 272 18541 278 18595
rect 332 18541 2642 18595
rect 2696 18541 2702 18595
rect 2636 18529 2702 18541
rect 3475 18500 3517 18653
rect 3704 18693 3741 18727
rect 3808 18693 3813 18727
rect 3704 18684 3756 18693
rect 3808 18684 3820 18693
rect 3872 18684 3884 18736
rect 3936 18684 3948 18736
rect 4000 18684 4012 18736
rect 4064 18684 4076 18736
rect 4128 18727 4140 18736
rect 4192 18727 4244 18736
rect 4135 18693 4140 18727
rect 4207 18693 4244 18727
rect 4128 18684 4140 18693
rect 4192 18684 4244 18693
rect 3704 18640 4244 18684
rect 3559 18535 3565 18587
rect 3617 18580 3623 18587
rect 4306 18580 4345 18970
rect 4558 18938 4597 19074
rect 4628 19043 4680 19049
rect 4625 18994 4628 19040
rect 4680 18994 4683 19040
rect 4875 18998 4904 19074
rect 4628 18985 4680 18991
rect 4875 18970 4980 18998
rect 4396 18905 4442 18938
rect 4396 18871 4402 18905
rect 4436 18871 4442 18905
rect 4396 18838 4442 18871
rect 4554 18918 4600 18938
rect 4704 18918 4750 18938
rect 4862 18918 4908 18938
rect 4554 18905 4750 18918
rect 4554 18871 4560 18905
rect 4594 18871 4710 18905
rect 4744 18871 4750 18905
rect 4554 18852 4750 18871
rect 4856 18866 4862 18918
rect 4914 18866 4920 18918
rect 4554 18838 4600 18852
rect 4704 18838 4750 18852
rect 4862 18838 4908 18866
rect 4402 18688 4430 18838
rect 4558 18793 4597 18838
rect 4552 18787 4604 18793
rect 4552 18729 4604 18735
rect 4952 18688 4980 18970
rect 5026 18920 5056 19105
rect 5694 19074 5740 19122
rect 5852 19228 5898 19274
rect 5852 19194 5858 19228
rect 5892 19194 5898 19228
rect 5852 19156 5898 19194
rect 5852 19122 5858 19156
rect 5892 19122 5898 19156
rect 5852 19074 5898 19122
rect 6002 19228 6048 19330
rect 6516 19274 6556 19480
rect 6862 19474 6868 19480
rect 6920 19474 6926 19526
rect 6985 19514 7015 19567
rect 6985 19485 7016 19514
rect 6002 19194 6008 19228
rect 6042 19194 6048 19228
rect 6002 19156 6048 19194
rect 6002 19122 6008 19156
rect 6042 19122 6048 19156
rect 6002 19074 6048 19122
rect 6160 19228 6206 19274
rect 6160 19194 6166 19228
rect 6200 19194 6206 19228
rect 6354 19228 6400 19274
rect 6354 19202 6360 19228
rect 6160 19156 6206 19194
rect 6160 19122 6166 19156
rect 6200 19122 6206 19156
rect 6244 19200 6360 19202
rect 6244 19148 6250 19200
rect 6302 19194 6360 19200
rect 6394 19194 6400 19228
rect 6302 19156 6400 19194
rect 6302 19148 6360 19156
rect 6244 19146 6360 19148
rect 6160 19074 6206 19122
rect 6354 19122 6360 19146
rect 6394 19122 6400 19156
rect 6354 19074 6400 19122
rect 6512 19228 6558 19274
rect 6512 19194 6518 19228
rect 6552 19194 6558 19228
rect 6662 19228 6708 19274
rect 6662 19194 6668 19228
rect 6702 19194 6708 19228
rect 6512 19156 6708 19194
rect 6512 19122 6518 19156
rect 6552 19128 6668 19156
rect 6552 19122 6558 19128
rect 6512 19074 6558 19122
rect 6662 19122 6668 19128
rect 6702 19122 6708 19156
rect 6662 19074 6708 19122
rect 6820 19228 6866 19274
rect 6820 19194 6826 19228
rect 6860 19194 6866 19228
rect 6986 19198 7016 19485
rect 6820 19156 6866 19194
rect 6820 19122 6826 19156
rect 6860 19122 6866 19156
rect 6968 19146 6974 19198
rect 7026 19146 7032 19198
rect 6820 19074 6866 19122
rect 6984 19106 7016 19146
rect 5111 18989 5117 19041
rect 5169 19034 5175 19041
rect 5620 19034 5672 19046
rect 5169 19032 5672 19034
rect 5169 18998 5628 19032
rect 5662 18998 5672 19032
rect 5169 18995 5672 18998
rect 5169 18989 5175 18995
rect 5620 18984 5672 18995
rect 5856 19026 5894 19074
rect 5934 19032 5986 19038
rect 5928 19026 5934 19032
rect 5856 18986 5934 19026
rect 5856 18936 5894 18986
rect 5928 18980 5934 18986
rect 5986 18980 5992 19032
rect 6164 19018 6204 19074
rect 6258 19018 6306 19030
rect 6164 19016 6306 19018
rect 6164 18984 6264 19016
rect 5934 18974 5986 18980
rect 6164 18936 6204 18984
rect 6258 18982 6264 18984
rect 6298 18982 6306 19016
rect 6258 18970 6306 18982
rect 5009 18868 5015 18920
rect 5067 18868 5073 18920
rect 5694 18904 5740 18936
rect 5694 18870 5700 18904
rect 5734 18870 5740 18904
rect 4402 18660 4980 18688
rect 3617 18541 4345 18580
rect 3617 18535 3623 18541
rect 5021 18500 5063 18868
rect 5694 18836 5740 18870
rect 5852 18904 5898 18936
rect 5852 18870 5858 18904
rect 5892 18870 5898 18904
rect 6002 18904 6048 18936
rect 6002 18874 6008 18904
rect 5852 18836 5898 18870
rect 6000 18870 6008 18874
rect 6042 18870 6048 18904
rect 5694 18780 5738 18836
rect 6000 18780 6048 18870
rect 6160 18904 6206 18936
rect 6160 18870 6166 18904
rect 6200 18870 6206 18904
rect 6160 18836 6206 18870
rect 5662 18736 6202 18780
rect 5662 18728 5714 18736
rect 5766 18728 5778 18736
rect 5662 18694 5700 18728
rect 5766 18694 5772 18728
rect 5662 18684 5714 18694
rect 5766 18684 5778 18694
rect 5830 18684 5842 18736
rect 5894 18684 5906 18736
rect 5958 18684 5970 18736
rect 6022 18684 6034 18736
rect 6086 18728 6098 18736
rect 6150 18728 6202 18736
rect 6094 18694 6098 18728
rect 6166 18694 6202 18728
rect 6086 18684 6098 18694
rect 6150 18684 6202 18694
rect 5662 18640 6202 18684
rect 5111 18535 5117 18587
rect 5169 18580 5175 18587
rect 6264 18580 6304 18970
rect 6516 18938 6556 19074
rect 6586 19044 6638 19050
rect 6584 18994 6586 19040
rect 6638 18994 6642 19040
rect 6834 18998 6862 19074
rect 6586 18986 6638 18992
rect 6834 18970 6936 18998
rect 6354 18906 6400 18938
rect 6354 18872 6360 18906
rect 6394 18872 6400 18906
rect 6354 18838 6400 18872
rect 6512 18918 6558 18938
rect 6662 18918 6708 18938
rect 6820 18918 6866 18938
rect 6512 18906 6708 18918
rect 6512 18872 6518 18906
rect 6552 18872 6668 18906
rect 6702 18872 6708 18906
rect 6512 18852 6708 18872
rect 6814 18866 6820 18918
rect 6872 18866 6878 18918
rect 6512 18838 6558 18852
rect 6662 18838 6708 18852
rect 6820 18838 6866 18866
rect 6360 18688 6388 18838
rect 6516 18794 6556 18838
rect 6510 18788 6562 18794
rect 6510 18730 6562 18736
rect 6908 18688 6936 18970
rect 6984 18920 7014 19106
rect 6968 18868 6974 18920
rect 7026 18868 7032 18920
rect 6360 18660 6936 18688
rect 6908 18596 6936 18660
rect 5169 18542 6304 18580
rect 6346 18568 6936 18596
rect 5169 18541 5572 18542
rect 5169 18535 5175 18541
rect 3475 18458 5063 18500
rect 5035 18417 5087 18423
rect 3472 18333 4907 18372
rect 6346 18405 6374 18568
rect 6908 18566 6936 18568
rect 6512 18502 6564 18508
rect 6512 18444 6564 18450
rect 5087 18377 6374 18405
rect 6523 18387 6553 18444
rect 5035 18359 5087 18365
rect 6523 18357 7015 18387
rect 1348 18199 1880 18242
rect 1348 18190 1398 18199
rect 1450 18190 1462 18199
rect 1348 18156 1383 18190
rect 1450 18156 1455 18190
rect 1348 18147 1398 18156
rect 1450 18147 1462 18156
rect 1514 18147 1526 18199
rect 1578 18147 1590 18199
rect 1642 18147 1654 18199
rect 1706 18147 1718 18199
rect 1770 18190 1782 18199
rect 1834 18190 1880 18199
rect 1777 18156 1782 18190
rect 1849 18156 1880 18190
rect 3472 18175 3511 18333
rect 4738 18291 4744 18298
rect 4558 18252 4744 18291
rect 1770 18147 1782 18156
rect 1834 18147 1880 18156
rect 550 18128 622 18132
rect 550 18076 560 18128
rect 612 18076 622 18128
rect 696 18126 768 18132
rect 550 18064 566 18076
rect 607 18064 622 18076
rect 682 18124 768 18126
rect 682 18072 702 18124
rect 754 18072 768 18124
rect 682 18070 710 18072
rect 550 18034 622 18064
rect 696 18064 710 18070
rect 751 18064 768 18072
rect 696 18034 768 18064
rect 840 18109 912 18138
rect 840 18069 856 18109
rect 897 18069 912 18109
rect 840 18040 912 18069
rect 994 18109 1066 18138
rect 994 18069 1009 18109
rect 1050 18069 1066 18109
rect 1348 18102 1880 18147
rect 994 18040 1066 18069
rect 564 17994 608 18034
rect 856 17974 900 18040
rect 378 17966 433 17972
rect 846 17922 852 17974
rect 904 17922 910 17974
rect 378 17681 433 17911
rect 856 17882 900 17922
rect 1008 17882 1052 18040
rect 1407 18036 1448 18102
rect 1693 18036 1735 18102
rect 1941 18099 2687 18144
rect 1404 17989 1450 18036
rect 1404 17955 1410 17989
rect 1444 17955 1450 17989
rect 1404 17917 1450 17955
rect 1404 17883 1410 17917
rect 1444 17883 1450 17917
rect 708 17838 900 17882
rect 372 17626 378 17681
rect 433 17626 439 17681
rect 708 17604 752 17838
rect 998 17830 1004 17882
rect 1056 17830 1062 17882
rect 1404 17836 1450 17883
rect 1562 17989 1608 18036
rect 1562 17955 1568 17989
rect 1602 17955 1608 17989
rect 1562 17917 1608 17955
rect 1562 17883 1568 17917
rect 1602 17883 1608 17917
rect 1562 17836 1608 17883
rect 1692 17989 1738 18036
rect 1692 17955 1698 17989
rect 1732 17955 1738 17989
rect 1692 17917 1738 17955
rect 1692 17883 1698 17917
rect 1732 17883 1738 17917
rect 1692 17836 1738 17883
rect 1850 18033 1896 18036
rect 1941 18033 1986 18099
rect 1850 17989 1986 18033
rect 1850 17955 1856 17989
rect 1890 17988 1986 17989
rect 2024 17989 2070 18036
rect 1890 17955 1896 17988
rect 1850 17917 1896 17955
rect 2024 17955 2030 17989
rect 2064 17955 2070 17989
rect 2024 17920 2070 17955
rect 1998 17918 2070 17920
rect 1850 17883 1856 17917
rect 1890 17883 1896 17917
rect 1850 17836 1896 17883
rect 1928 17917 2070 17918
rect 1928 17893 2030 17917
rect 1928 17876 1935 17893
rect 1929 17841 1935 17876
rect 1987 17883 2030 17893
rect 2064 17883 2070 17917
rect 1987 17876 2070 17883
rect 1987 17841 1993 17876
rect 2024 17836 2070 17876
rect 2182 17992 2228 18036
rect 2366 17992 2412 18036
rect 2182 17989 2412 17992
rect 2182 17955 2188 17989
rect 2222 17955 2372 17989
rect 2406 17955 2412 17989
rect 2182 17917 2412 17955
rect 2182 17883 2188 17917
rect 2222 17883 2372 17917
rect 2406 17883 2412 17917
rect 2182 17866 2412 17883
rect 2182 17836 2228 17866
rect 2366 17836 2412 17866
rect 2524 17989 2570 18036
rect 2524 17955 2530 17989
rect 2564 17955 2570 17989
rect 2642 17965 2687 18099
rect 3118 18136 3511 18175
rect 3724 18198 4264 18242
rect 3724 18146 3776 18198
rect 3828 18189 3840 18198
rect 3892 18189 3904 18198
rect 3956 18189 3968 18198
rect 4020 18189 4032 18198
rect 4084 18189 4096 18198
rect 4148 18189 4160 18198
rect 3831 18155 3840 18189
rect 3903 18155 3904 18189
rect 4084 18155 4085 18189
rect 4148 18155 4157 18189
rect 3828 18146 3840 18155
rect 3892 18146 3904 18155
rect 3956 18146 3968 18155
rect 4020 18146 4032 18155
rect 4084 18146 4096 18155
rect 4148 18146 4160 18155
rect 4212 18146 4264 18198
rect 2774 18092 2816 18093
rect 2758 18084 2816 18092
rect 2758 18032 2769 18084
rect 2821 18032 2827 18084
rect 3118 18036 3157 18136
rect 3724 18102 4264 18146
rect 3741 18046 3787 18102
rect 3736 18045 3787 18046
rect 2758 17989 2816 18032
rect 2524 17917 2570 17955
rect 2524 17883 2530 17917
rect 2564 17883 2570 17917
rect 2524 17876 2570 17883
rect 2613 17937 2715 17965
rect 2613 17903 2647 17937
rect 2681 17903 2715 17937
rect 2524 17836 2574 17876
rect 2613 17875 2715 17903
rect 2758 17955 2776 17989
rect 2810 17955 2816 17989
rect 2758 17917 2816 17955
rect 2758 17883 2776 17917
rect 2810 17883 2816 17917
rect 1008 17776 1052 17830
rect 1245 17795 1328 17814
rect 852 17732 1052 17776
rect 1148 17793 1328 17795
rect 1148 17741 1155 17793
rect 1207 17783 1328 17793
rect 1207 17749 1269 17783
rect 1303 17749 1328 17783
rect 1207 17741 1328 17749
rect 1148 17740 1328 17741
rect 852 17610 896 17732
rect 1245 17719 1328 17740
rect 1568 17802 1602 17836
rect 1568 17792 1820 17802
rect 1568 17740 1758 17792
rect 1810 17740 1820 17792
rect 1568 17730 1820 17740
rect 1568 17698 1608 17730
rect 1853 17698 1892 17836
rect 2185 17698 2224 17836
rect 2255 17799 2325 17805
rect 2255 17790 2331 17799
rect 2255 17738 2270 17790
rect 2322 17738 2331 17790
rect 2255 17729 2331 17738
rect 2255 17723 2325 17729
rect 2368 17698 2407 17836
rect 2530 17802 2574 17836
rect 2758 17836 2816 17883
rect 2928 17989 2974 18036
rect 2928 17955 2934 17989
rect 2968 17976 2974 17989
rect 3114 17989 3160 18036
rect 3114 17976 3120 17989
rect 2968 17955 3120 17976
rect 3154 17955 3160 17989
rect 3272 17989 3318 18036
rect 3272 17979 3278 17989
rect 3312 17979 3318 17989
rect 3736 17999 3782 18045
rect 2928 17917 3160 17955
rect 3262 17927 3268 17979
rect 3320 17927 3326 17979
rect 3736 17965 3742 17999
rect 3776 17965 3782 17999
rect 3736 17927 3782 17965
rect 2928 17883 2934 17917
rect 2968 17883 3120 17917
rect 3154 17883 3160 17917
rect 2928 17866 3160 17883
rect 2928 17836 2974 17866
rect 3114 17836 3160 17866
rect 3272 17917 3318 17927
rect 3272 17883 3278 17917
rect 3312 17883 3318 17917
rect 3272 17836 3318 17883
rect 3736 17893 3742 17927
rect 3776 17893 3782 17927
rect 3736 17846 3782 17893
rect 3894 17999 3940 18046
rect 3894 17965 3900 17999
rect 3934 17965 3940 17999
rect 3894 17927 3940 17965
rect 3894 17893 3900 17927
rect 3934 17893 3940 17927
rect 3894 17846 3940 17893
rect 4044 17999 4090 18102
rect 4558 18046 4597 18252
rect 4738 18246 4744 18252
rect 4796 18246 4802 18298
rect 4868 18046 4907 18333
rect 6837 18291 6843 18298
rect 6516 18252 6843 18291
rect 5682 18198 6222 18242
rect 5682 18146 5734 18198
rect 5786 18188 5798 18198
rect 5850 18188 5862 18198
rect 5914 18188 5926 18198
rect 5978 18188 5990 18198
rect 6042 18188 6054 18198
rect 6106 18188 6118 18198
rect 5790 18154 5798 18188
rect 6042 18154 6044 18188
rect 6106 18154 6116 18188
rect 5786 18146 5798 18154
rect 5850 18146 5862 18154
rect 5914 18146 5926 18154
rect 5978 18146 5990 18154
rect 6042 18146 6054 18154
rect 6106 18146 6118 18154
rect 6170 18146 6222 18198
rect 5682 18102 6222 18146
rect 5700 18046 5746 18102
rect 4044 17965 4050 17999
rect 4084 17965 4090 17999
rect 4044 17927 4090 17965
rect 4044 17893 4050 17927
rect 4084 17893 4090 17927
rect 4044 17846 4090 17893
rect 4202 17999 4248 18046
rect 4202 17965 4208 17999
rect 4242 17965 4248 17999
rect 4396 17999 4442 18046
rect 4396 17973 4402 17999
rect 4202 17927 4248 17965
rect 4202 17893 4208 17927
rect 4242 17893 4248 17927
rect 4285 17971 4402 17973
rect 4285 17919 4292 17971
rect 4344 17965 4402 17971
rect 4436 17965 4442 17999
rect 4344 17927 4442 17965
rect 4344 17919 4402 17927
rect 4285 17918 4402 17919
rect 4202 17846 4248 17893
rect 4396 17893 4402 17918
rect 4436 17893 4442 17927
rect 4396 17846 4442 17893
rect 4554 17999 4600 18046
rect 4554 17965 4560 17999
rect 4594 17966 4600 17999
rect 4704 17999 4750 18046
rect 4704 17966 4710 17999
rect 4594 17965 4710 17966
rect 4744 17965 4750 17999
rect 4554 17927 4750 17965
rect 4554 17893 4560 17927
rect 4594 17900 4710 17927
rect 4594 17893 4600 17900
rect 4554 17846 4600 17893
rect 4704 17893 4710 17900
rect 4744 17893 4750 17927
rect 4704 17846 4750 17893
rect 4862 17999 4908 18046
rect 4862 17965 4868 17999
rect 4902 17965 4908 17999
rect 5694 18000 5740 18046
rect 5027 17970 5057 17979
rect 4862 17927 4908 17965
rect 4862 17893 4868 17927
rect 4902 17893 4908 17927
rect 5010 17918 5016 17970
rect 5068 17918 5074 17970
rect 5694 17966 5700 18000
rect 5734 17966 5740 18000
rect 5694 17928 5740 17966
rect 4862 17846 4908 17893
rect 5026 17877 5057 17918
rect 5694 17894 5700 17928
rect 5734 17894 5740 17928
rect 2758 17802 2802 17836
rect 2530 17758 2656 17802
rect 1242 17678 1248 17682
rect 1138 17634 1248 17678
rect 1138 17610 1182 17634
rect 1242 17630 1248 17634
rect 1300 17630 1306 17682
rect 1404 17665 1450 17698
rect 1404 17631 1410 17665
rect 1444 17631 1450 17665
rect 1404 17627 1450 17631
rect 378 17582 434 17588
rect 550 17582 622 17604
rect 434 17576 622 17582
rect 434 17536 565 17576
rect 606 17536 622 17576
rect 434 17526 622 17536
rect 378 17520 434 17526
rect 550 17506 622 17526
rect 696 17576 768 17604
rect 696 17536 712 17576
rect 753 17536 768 17576
rect 696 17506 768 17536
rect 840 17581 912 17610
rect 840 17541 856 17581
rect 897 17541 912 17581
rect 840 17512 912 17541
rect 994 17582 1182 17610
rect 994 17542 1010 17582
rect 1051 17566 1182 17582
rect 1399 17598 1450 17627
rect 1562 17665 1608 17698
rect 1562 17631 1568 17665
rect 1602 17631 1608 17665
rect 1692 17665 1738 17698
rect 1692 17636 1698 17665
rect 1562 17598 1608 17631
rect 1690 17631 1698 17636
rect 1732 17636 1738 17665
rect 1850 17665 1896 17698
rect 2024 17682 2070 17698
rect 1732 17631 1740 17636
rect 1051 17542 1066 17566
rect 1399 17552 1449 17598
rect 1690 17552 1740 17631
rect 1850 17631 1856 17665
rect 1890 17631 1896 17665
rect 1850 17598 1896 17631
rect 2014 17630 2020 17682
rect 2072 17630 2078 17682
rect 2182 17665 2228 17698
rect 2182 17631 2188 17665
rect 2222 17631 2228 17665
rect 2024 17598 2070 17630
rect 2182 17598 2228 17631
rect 2366 17665 2412 17698
rect 2524 17680 2570 17698
rect 2366 17631 2372 17665
rect 2406 17631 2412 17665
rect 2366 17598 2412 17631
rect 2516 17628 2522 17680
rect 2574 17628 2580 17680
rect 2524 17598 2570 17628
rect 2024 17566 2068 17598
rect 2612 17566 2656 17758
rect 994 17512 1066 17542
rect 1324 17497 1960 17552
rect 2024 17522 2656 17566
rect 2694 17758 2802 17802
rect 2832 17788 2904 17798
rect 2694 17560 2738 17758
rect 2832 17736 2842 17788
rect 2894 17736 2904 17788
rect 2832 17726 2904 17736
rect 2933 17698 2972 17836
rect 3118 17698 3157 17836
rect 3272 17792 3316 17836
rect 3268 17786 3320 17792
rect 3555 17761 3561 17813
rect 3613 17806 3619 17813
rect 3662 17806 3713 17818
rect 3613 17803 3713 17806
rect 3613 17769 3670 17803
rect 3704 17769 3713 17803
rect 3613 17767 3713 17769
rect 3613 17761 3619 17767
rect 3662 17755 3713 17767
rect 3897 17797 3936 17846
rect 3976 17804 4027 17809
rect 3970 17797 3976 17804
rect 3897 17758 3976 17797
rect 3268 17728 3320 17734
rect 3897 17708 3936 17758
rect 3970 17752 3976 17758
rect 4028 17752 4034 17804
rect 4206 17790 4245 17846
rect 4300 17790 4347 17801
rect 4206 17788 4347 17790
rect 4206 17755 4306 17788
rect 3976 17746 4027 17752
rect 4206 17708 4245 17755
rect 4300 17754 4306 17755
rect 4340 17754 4347 17788
rect 4300 17742 4347 17754
rect 2766 17692 2818 17698
rect 2766 17634 2776 17640
rect 2770 17631 2776 17634
rect 2810 17634 2818 17640
rect 2928 17665 2974 17698
rect 2810 17631 2816 17634
rect 2770 17598 2816 17631
rect 2928 17631 2934 17665
rect 2968 17631 2974 17665
rect 2928 17598 2974 17631
rect 3114 17665 3160 17698
rect 3114 17631 3120 17665
rect 3154 17631 3160 17665
rect 3114 17598 3160 17631
rect 3272 17665 3318 17698
rect 3272 17631 3278 17665
rect 3312 17631 3318 17665
rect 3272 17598 3318 17631
rect 3274 17560 3318 17598
rect 2694 17516 3318 17560
rect 3736 17675 3782 17708
rect 3736 17641 3742 17675
rect 3776 17641 3782 17675
rect 3736 17608 3782 17641
rect 3894 17675 3940 17708
rect 3894 17641 3900 17675
rect 3934 17641 3940 17675
rect 4044 17675 4090 17708
rect 4044 17646 4050 17675
rect 3894 17608 3940 17641
rect 4042 17641 4050 17646
rect 4084 17641 4090 17675
rect 4042 17608 4090 17641
rect 4202 17675 4248 17708
rect 4202 17641 4208 17675
rect 4242 17641 4248 17675
rect 4202 17608 4248 17641
rect 3736 17552 3780 17608
rect 4042 17552 4089 17608
rect 1324 17445 1360 17497
rect 1412 17445 1424 17497
rect 1476 17488 1488 17497
rect 1540 17488 1552 17497
rect 1604 17488 1616 17497
rect 1668 17488 1680 17497
rect 1732 17488 1744 17497
rect 1796 17488 1808 17497
rect 1479 17454 1488 17488
rect 1551 17454 1552 17488
rect 1732 17454 1733 17488
rect 1796 17454 1805 17488
rect 1476 17445 1488 17454
rect 1540 17445 1552 17454
rect 1604 17445 1616 17454
rect 1668 17445 1680 17454
rect 1732 17445 1744 17454
rect 1796 17445 1808 17454
rect 1860 17445 1872 17497
rect 1924 17445 1960 17497
rect 3704 17508 4244 17552
rect 3704 17499 3756 17508
rect 3808 17499 3820 17508
rect 1324 17412 1960 17445
rect 2346 17467 2426 17492
rect 2346 17463 3517 17467
rect 2346 17429 2369 17463
rect 2403 17429 3517 17463
rect 2346 17425 3517 17429
rect 2346 17400 2426 17425
rect 2636 17367 2702 17379
rect 272 17313 278 17367
rect 332 17313 2642 17367
rect 2696 17313 2702 17367
rect 2636 17301 2702 17313
rect 3475 17272 3517 17425
rect 3704 17465 3741 17499
rect 3808 17465 3813 17499
rect 3704 17456 3756 17465
rect 3808 17456 3820 17465
rect 3872 17456 3884 17508
rect 3936 17456 3948 17508
rect 4000 17456 4012 17508
rect 4064 17456 4076 17508
rect 4128 17499 4140 17508
rect 4192 17499 4244 17508
rect 4135 17465 4140 17499
rect 4207 17465 4244 17499
rect 4128 17456 4140 17465
rect 4192 17456 4244 17465
rect 3704 17412 4244 17456
rect 3559 17307 3565 17359
rect 3617 17352 3623 17359
rect 4306 17352 4345 17742
rect 4558 17710 4597 17846
rect 4628 17815 4680 17821
rect 4625 17766 4628 17812
rect 4680 17766 4683 17812
rect 4875 17770 4904 17846
rect 4628 17757 4680 17763
rect 4875 17742 4980 17770
rect 4396 17677 4442 17710
rect 4396 17643 4402 17677
rect 4436 17643 4442 17677
rect 4396 17610 4442 17643
rect 4554 17690 4600 17710
rect 4704 17690 4750 17710
rect 4862 17690 4908 17710
rect 4554 17677 4750 17690
rect 4554 17643 4560 17677
rect 4594 17643 4710 17677
rect 4744 17643 4750 17677
rect 4554 17624 4750 17643
rect 4856 17638 4862 17690
rect 4914 17638 4920 17690
rect 4554 17610 4600 17624
rect 4704 17610 4750 17624
rect 4862 17610 4908 17638
rect 4402 17460 4430 17610
rect 4558 17565 4597 17610
rect 4552 17559 4604 17565
rect 4552 17501 4604 17507
rect 4952 17460 4980 17742
rect 5026 17692 5056 17877
rect 5694 17846 5740 17894
rect 5852 18000 5898 18046
rect 5852 17966 5858 18000
rect 5892 17966 5898 18000
rect 5852 17928 5898 17966
rect 5852 17894 5858 17928
rect 5892 17894 5898 17928
rect 5852 17846 5898 17894
rect 6002 18000 6048 18102
rect 6516 18046 6556 18252
rect 6837 18246 6843 18252
rect 6895 18246 6901 18298
rect 6985 18286 7015 18357
rect 6985 18257 7016 18286
rect 6002 17966 6008 18000
rect 6042 17966 6048 18000
rect 6002 17928 6048 17966
rect 6002 17894 6008 17928
rect 6042 17894 6048 17928
rect 6002 17846 6048 17894
rect 6160 18000 6206 18046
rect 6160 17966 6166 18000
rect 6200 17966 6206 18000
rect 6354 18000 6400 18046
rect 6354 17974 6360 18000
rect 6160 17928 6206 17966
rect 6160 17894 6166 17928
rect 6200 17894 6206 17928
rect 6244 17972 6360 17974
rect 6244 17920 6250 17972
rect 6302 17966 6360 17972
rect 6394 17966 6400 18000
rect 6302 17928 6400 17966
rect 6302 17920 6360 17928
rect 6244 17918 6360 17920
rect 6160 17846 6206 17894
rect 6354 17894 6360 17918
rect 6394 17894 6400 17928
rect 6354 17846 6400 17894
rect 6512 18000 6558 18046
rect 6512 17966 6518 18000
rect 6552 17966 6558 18000
rect 6662 18000 6708 18046
rect 6662 17966 6668 18000
rect 6702 17966 6708 18000
rect 6512 17928 6708 17966
rect 6512 17894 6518 17928
rect 6552 17900 6668 17928
rect 6552 17894 6558 17900
rect 6512 17846 6558 17894
rect 6662 17894 6668 17900
rect 6702 17894 6708 17928
rect 6662 17846 6708 17894
rect 6820 18000 6866 18046
rect 6820 17966 6826 18000
rect 6860 17966 6866 18000
rect 6986 17970 7016 18257
rect 6820 17928 6866 17966
rect 6820 17894 6826 17928
rect 6860 17894 6866 17928
rect 6968 17918 6974 17970
rect 7026 17918 7032 17970
rect 6820 17846 6866 17894
rect 6984 17878 7016 17918
rect 5191 17761 5197 17813
rect 5249 17806 5255 17813
rect 5620 17806 5672 17818
rect 5249 17804 5672 17806
rect 5249 17770 5628 17804
rect 5662 17770 5672 17804
rect 5249 17767 5672 17770
rect 5249 17761 5255 17767
rect 5620 17756 5672 17767
rect 5856 17798 5894 17846
rect 5934 17804 5986 17810
rect 5928 17798 5934 17804
rect 5856 17758 5934 17798
rect 5856 17708 5894 17758
rect 5928 17752 5934 17758
rect 5986 17752 5992 17804
rect 6164 17790 6204 17846
rect 6258 17790 6306 17802
rect 6164 17788 6306 17790
rect 6164 17756 6264 17788
rect 5934 17746 5986 17752
rect 6164 17708 6204 17756
rect 6258 17754 6264 17756
rect 6298 17754 6306 17788
rect 6258 17742 6306 17754
rect 5009 17640 5015 17692
rect 5067 17640 5073 17692
rect 5694 17676 5740 17708
rect 5694 17642 5700 17676
rect 5734 17642 5740 17676
rect 4402 17432 4980 17460
rect 3617 17313 4345 17352
rect 3617 17307 3623 17313
rect 5021 17272 5063 17640
rect 5694 17608 5740 17642
rect 5852 17676 5898 17708
rect 5852 17642 5858 17676
rect 5892 17642 5898 17676
rect 6002 17676 6048 17708
rect 6002 17646 6008 17676
rect 5852 17608 5898 17642
rect 6000 17642 6008 17646
rect 6042 17642 6048 17676
rect 5694 17552 5738 17608
rect 6000 17552 6048 17642
rect 6160 17676 6206 17708
rect 6160 17642 6166 17676
rect 6200 17642 6206 17676
rect 6160 17608 6206 17642
rect 5662 17508 6202 17552
rect 5662 17500 5714 17508
rect 5766 17500 5778 17508
rect 5662 17466 5700 17500
rect 5766 17466 5772 17500
rect 5662 17456 5714 17466
rect 5766 17456 5778 17466
rect 5830 17456 5842 17508
rect 5894 17456 5906 17508
rect 5958 17456 5970 17508
rect 6022 17456 6034 17508
rect 6086 17500 6098 17508
rect 6150 17500 6202 17508
rect 6094 17466 6098 17500
rect 6166 17466 6202 17500
rect 6086 17456 6098 17466
rect 6150 17456 6202 17466
rect 5662 17412 6202 17456
rect 5191 17307 5197 17359
rect 5249 17352 5255 17359
rect 6264 17352 6304 17742
rect 6516 17710 6556 17846
rect 6586 17816 6638 17822
rect 6584 17766 6586 17812
rect 6638 17766 6642 17812
rect 6834 17770 6862 17846
rect 6586 17758 6638 17764
rect 6834 17742 6936 17770
rect 6354 17678 6400 17710
rect 6354 17644 6360 17678
rect 6394 17644 6400 17678
rect 6354 17610 6400 17644
rect 6512 17690 6558 17710
rect 6662 17690 6708 17710
rect 6820 17690 6866 17710
rect 6512 17678 6708 17690
rect 6512 17644 6518 17678
rect 6552 17644 6668 17678
rect 6702 17644 6708 17678
rect 6512 17624 6708 17644
rect 6814 17638 6820 17690
rect 6872 17638 6878 17690
rect 6512 17610 6558 17624
rect 6662 17610 6708 17624
rect 6820 17610 6866 17638
rect 6360 17460 6388 17610
rect 6516 17566 6556 17610
rect 6510 17560 6562 17566
rect 6510 17502 6562 17508
rect 6908 17460 6936 17742
rect 6984 17692 7014 17878
rect 6968 17640 6974 17692
rect 7026 17640 7032 17692
rect 6360 17432 6936 17460
rect 5249 17314 6304 17352
rect 5249 17313 5587 17314
rect 5249 17307 5255 17313
rect 3475 17230 5063 17272
rect 6908 17260 6936 17432
rect 7107 17272 7159 17278
rect 6908 17232 7107 17260
rect 7107 17214 7159 17220
rect 5029 17152 5081 17158
rect 3472 17105 4907 17144
rect 1348 16971 1880 17014
rect 1348 16962 1398 16971
rect 1450 16962 1462 16971
rect 1348 16928 1383 16962
rect 1450 16928 1455 16962
rect 1348 16919 1398 16928
rect 1450 16919 1462 16928
rect 1514 16919 1526 16971
rect 1578 16919 1590 16971
rect 1642 16919 1654 16971
rect 1706 16919 1718 16971
rect 1770 16962 1782 16971
rect 1834 16962 1880 16971
rect 1777 16928 1782 16962
rect 1849 16928 1880 16962
rect 3472 16947 3511 17105
rect 4738 17063 4744 17070
rect 4558 17024 4744 17063
rect 1770 16919 1782 16928
rect 1834 16919 1880 16928
rect 550 16900 622 16904
rect 550 16848 560 16900
rect 612 16848 622 16900
rect 696 16898 768 16904
rect 550 16836 566 16848
rect 607 16836 622 16848
rect 682 16896 768 16898
rect 682 16844 702 16896
rect 754 16844 768 16896
rect 682 16842 710 16844
rect 550 16806 622 16836
rect 696 16836 710 16842
rect 751 16836 768 16844
rect 696 16806 768 16836
rect 840 16881 912 16910
rect 840 16841 856 16881
rect 897 16841 912 16881
rect 840 16812 912 16841
rect 994 16881 1066 16910
rect 994 16841 1009 16881
rect 1050 16841 1066 16881
rect 1348 16874 1880 16919
rect 994 16812 1066 16841
rect 564 16766 608 16806
rect 856 16746 900 16812
rect 378 16738 433 16744
rect 846 16694 852 16746
rect 904 16694 910 16746
rect 378 16453 433 16683
rect 856 16654 900 16694
rect 1008 16654 1052 16812
rect 1407 16808 1448 16874
rect 1693 16808 1735 16874
rect 1941 16871 2687 16916
rect 1404 16761 1450 16808
rect 1404 16727 1410 16761
rect 1444 16727 1450 16761
rect 1404 16689 1450 16727
rect 1404 16655 1410 16689
rect 1444 16655 1450 16689
rect 708 16610 900 16654
rect 372 16398 378 16453
rect 433 16398 439 16453
rect 708 16376 752 16610
rect 998 16602 1004 16654
rect 1056 16602 1062 16654
rect 1404 16608 1450 16655
rect 1562 16761 1608 16808
rect 1562 16727 1568 16761
rect 1602 16727 1608 16761
rect 1562 16689 1608 16727
rect 1562 16655 1568 16689
rect 1602 16655 1608 16689
rect 1562 16608 1608 16655
rect 1692 16761 1738 16808
rect 1692 16727 1698 16761
rect 1732 16727 1738 16761
rect 1692 16689 1738 16727
rect 1692 16655 1698 16689
rect 1732 16655 1738 16689
rect 1692 16608 1738 16655
rect 1850 16805 1896 16808
rect 1941 16805 1986 16871
rect 1850 16761 1986 16805
rect 1850 16727 1856 16761
rect 1890 16760 1986 16761
rect 2024 16761 2070 16808
rect 1890 16727 1896 16760
rect 1850 16689 1896 16727
rect 2024 16727 2030 16761
rect 2064 16727 2070 16761
rect 2024 16692 2070 16727
rect 1998 16690 2070 16692
rect 1850 16655 1856 16689
rect 1890 16655 1896 16689
rect 1850 16608 1896 16655
rect 1928 16689 2070 16690
rect 1928 16665 2030 16689
rect 1928 16648 1935 16665
rect 1929 16613 1935 16648
rect 1987 16655 2030 16665
rect 2064 16655 2070 16689
rect 1987 16648 2070 16655
rect 1987 16613 1993 16648
rect 2024 16608 2070 16648
rect 2182 16764 2228 16808
rect 2366 16764 2412 16808
rect 2182 16761 2412 16764
rect 2182 16727 2188 16761
rect 2222 16727 2372 16761
rect 2406 16727 2412 16761
rect 2182 16689 2412 16727
rect 2182 16655 2188 16689
rect 2222 16655 2372 16689
rect 2406 16655 2412 16689
rect 2182 16638 2412 16655
rect 2182 16608 2228 16638
rect 2366 16608 2412 16638
rect 2524 16761 2570 16808
rect 2524 16727 2530 16761
rect 2564 16727 2570 16761
rect 2642 16737 2687 16871
rect 3118 16908 3511 16947
rect 3724 16970 4264 17014
rect 3724 16918 3776 16970
rect 3828 16961 3840 16970
rect 3892 16961 3904 16970
rect 3956 16961 3968 16970
rect 4020 16961 4032 16970
rect 4084 16961 4096 16970
rect 4148 16961 4160 16970
rect 3831 16927 3840 16961
rect 3903 16927 3904 16961
rect 4084 16927 4085 16961
rect 4148 16927 4157 16961
rect 3828 16918 3840 16927
rect 3892 16918 3904 16927
rect 3956 16918 3968 16927
rect 4020 16918 4032 16927
rect 4084 16918 4096 16927
rect 4148 16918 4160 16927
rect 4212 16918 4264 16970
rect 2774 16864 2816 16865
rect 2758 16856 2816 16864
rect 2758 16804 2769 16856
rect 2821 16804 2827 16856
rect 3118 16808 3157 16908
rect 3724 16874 4264 16918
rect 3741 16818 3787 16874
rect 3736 16817 3787 16818
rect 2758 16761 2816 16804
rect 2524 16689 2570 16727
rect 2524 16655 2530 16689
rect 2564 16655 2570 16689
rect 2524 16648 2570 16655
rect 2613 16709 2715 16737
rect 2613 16675 2647 16709
rect 2681 16675 2715 16709
rect 2524 16608 2574 16648
rect 2613 16647 2715 16675
rect 2758 16727 2776 16761
rect 2810 16727 2816 16761
rect 2758 16689 2816 16727
rect 2758 16655 2776 16689
rect 2810 16655 2816 16689
rect 1008 16548 1052 16602
rect 1245 16567 1328 16586
rect 852 16504 1052 16548
rect 1148 16565 1328 16567
rect 1148 16513 1155 16565
rect 1207 16555 1328 16565
rect 1207 16521 1269 16555
rect 1303 16521 1328 16555
rect 1207 16513 1328 16521
rect 1148 16512 1328 16513
rect 852 16382 896 16504
rect 1245 16491 1328 16512
rect 1568 16574 1602 16608
rect 1568 16564 1820 16574
rect 1568 16512 1758 16564
rect 1810 16512 1820 16564
rect 1568 16502 1820 16512
rect 1568 16470 1608 16502
rect 1853 16470 1892 16608
rect 2185 16470 2224 16608
rect 2255 16571 2325 16577
rect 2255 16562 2331 16571
rect 2255 16510 2270 16562
rect 2322 16510 2331 16562
rect 2255 16501 2331 16510
rect 2255 16495 2325 16501
rect 2368 16470 2407 16608
rect 2530 16574 2574 16608
rect 2758 16608 2816 16655
rect 2928 16761 2974 16808
rect 2928 16727 2934 16761
rect 2968 16748 2974 16761
rect 3114 16761 3160 16808
rect 3114 16748 3120 16761
rect 2968 16727 3120 16748
rect 3154 16727 3160 16761
rect 3272 16761 3318 16808
rect 3272 16751 3278 16761
rect 3312 16751 3318 16761
rect 3736 16771 3782 16817
rect 2928 16689 3160 16727
rect 3262 16699 3268 16751
rect 3320 16699 3326 16751
rect 3736 16737 3742 16771
rect 3776 16737 3782 16771
rect 3736 16699 3782 16737
rect 2928 16655 2934 16689
rect 2968 16655 3120 16689
rect 3154 16655 3160 16689
rect 2928 16638 3160 16655
rect 2928 16608 2974 16638
rect 3114 16608 3160 16638
rect 3272 16689 3318 16699
rect 3272 16655 3278 16689
rect 3312 16655 3318 16689
rect 3272 16608 3318 16655
rect 3736 16665 3742 16699
rect 3776 16665 3782 16699
rect 3736 16618 3782 16665
rect 3894 16771 3940 16818
rect 3894 16737 3900 16771
rect 3934 16737 3940 16771
rect 3894 16699 3940 16737
rect 3894 16665 3900 16699
rect 3934 16665 3940 16699
rect 3894 16618 3940 16665
rect 4044 16771 4090 16874
rect 4558 16818 4597 17024
rect 4738 17018 4744 17024
rect 4796 17018 4802 17070
rect 4868 16818 4907 17105
rect 5081 17111 7015 17141
rect 5029 17094 5081 17100
rect 6862 17063 6868 17070
rect 6516 17024 6868 17063
rect 5682 16970 6222 17014
rect 5682 16918 5734 16970
rect 5786 16960 5798 16970
rect 5850 16960 5862 16970
rect 5914 16960 5926 16970
rect 5978 16960 5990 16970
rect 6042 16960 6054 16970
rect 6106 16960 6118 16970
rect 5790 16926 5798 16960
rect 6042 16926 6044 16960
rect 6106 16926 6116 16960
rect 5786 16918 5798 16926
rect 5850 16918 5862 16926
rect 5914 16918 5926 16926
rect 5978 16918 5990 16926
rect 6042 16918 6054 16926
rect 6106 16918 6118 16926
rect 6170 16918 6222 16970
rect 5682 16874 6222 16918
rect 5700 16818 5746 16874
rect 4044 16737 4050 16771
rect 4084 16737 4090 16771
rect 4044 16699 4090 16737
rect 4044 16665 4050 16699
rect 4084 16665 4090 16699
rect 4044 16618 4090 16665
rect 4202 16771 4248 16818
rect 4202 16737 4208 16771
rect 4242 16737 4248 16771
rect 4396 16771 4442 16818
rect 4396 16745 4402 16771
rect 4202 16699 4248 16737
rect 4202 16665 4208 16699
rect 4242 16665 4248 16699
rect 4285 16743 4402 16745
rect 4285 16691 4292 16743
rect 4344 16737 4402 16743
rect 4436 16737 4442 16771
rect 4344 16699 4442 16737
rect 4344 16691 4402 16699
rect 4285 16690 4402 16691
rect 4202 16618 4248 16665
rect 4396 16665 4402 16690
rect 4436 16665 4442 16699
rect 4396 16618 4442 16665
rect 4554 16771 4600 16818
rect 4554 16737 4560 16771
rect 4594 16738 4600 16771
rect 4704 16771 4750 16818
rect 4704 16738 4710 16771
rect 4594 16737 4710 16738
rect 4744 16737 4750 16771
rect 4554 16699 4750 16737
rect 4554 16665 4560 16699
rect 4594 16672 4710 16699
rect 4594 16665 4600 16672
rect 4554 16618 4600 16665
rect 4704 16665 4710 16672
rect 4744 16665 4750 16699
rect 4704 16618 4750 16665
rect 4862 16771 4908 16818
rect 4862 16737 4868 16771
rect 4902 16737 4908 16771
rect 5694 16772 5740 16818
rect 5027 16742 5057 16751
rect 4862 16699 4908 16737
rect 4862 16665 4868 16699
rect 4902 16665 4908 16699
rect 5010 16690 5016 16742
rect 5068 16690 5074 16742
rect 5694 16738 5700 16772
rect 5734 16738 5740 16772
rect 5694 16700 5740 16738
rect 4862 16618 4908 16665
rect 5026 16649 5057 16690
rect 5694 16666 5700 16700
rect 5734 16666 5740 16700
rect 2758 16574 2802 16608
rect 2530 16530 2656 16574
rect 1242 16450 1248 16454
rect 1138 16406 1248 16450
rect 1138 16382 1182 16406
rect 1242 16402 1248 16406
rect 1300 16402 1306 16454
rect 1404 16437 1450 16470
rect 1404 16403 1410 16437
rect 1444 16403 1450 16437
rect 1404 16399 1450 16403
rect 378 16354 434 16360
rect 550 16354 622 16376
rect 434 16348 622 16354
rect 434 16308 565 16348
rect 606 16308 622 16348
rect 434 16298 622 16308
rect 378 16292 434 16298
rect 550 16278 622 16298
rect 696 16348 768 16376
rect 696 16308 712 16348
rect 753 16308 768 16348
rect 696 16278 768 16308
rect 840 16353 912 16382
rect 840 16313 856 16353
rect 897 16313 912 16353
rect 840 16284 912 16313
rect 994 16354 1182 16382
rect 994 16314 1010 16354
rect 1051 16338 1182 16354
rect 1399 16370 1450 16399
rect 1562 16437 1608 16470
rect 1562 16403 1568 16437
rect 1602 16403 1608 16437
rect 1692 16437 1738 16470
rect 1692 16408 1698 16437
rect 1562 16370 1608 16403
rect 1690 16403 1698 16408
rect 1732 16408 1738 16437
rect 1850 16437 1896 16470
rect 2024 16454 2070 16470
rect 1732 16403 1740 16408
rect 1051 16314 1066 16338
rect 1399 16324 1449 16370
rect 1690 16324 1740 16403
rect 1850 16403 1856 16437
rect 1890 16403 1896 16437
rect 1850 16370 1896 16403
rect 2014 16402 2020 16454
rect 2072 16402 2078 16454
rect 2182 16437 2228 16470
rect 2182 16403 2188 16437
rect 2222 16403 2228 16437
rect 2024 16370 2070 16402
rect 2182 16370 2228 16403
rect 2366 16437 2412 16470
rect 2524 16452 2570 16470
rect 2366 16403 2372 16437
rect 2406 16403 2412 16437
rect 2366 16370 2412 16403
rect 2516 16400 2522 16452
rect 2574 16400 2580 16452
rect 2524 16370 2570 16400
rect 2024 16338 2068 16370
rect 2612 16338 2656 16530
rect 994 16284 1066 16314
rect 1324 16269 1960 16324
rect 2024 16294 2656 16338
rect 2694 16530 2802 16574
rect 2832 16560 2904 16570
rect 2694 16332 2738 16530
rect 2832 16508 2842 16560
rect 2894 16508 2904 16560
rect 2832 16498 2904 16508
rect 2933 16470 2972 16608
rect 3118 16470 3157 16608
rect 3272 16564 3316 16608
rect 3268 16558 3320 16564
rect 3555 16533 3561 16585
rect 3613 16578 3619 16585
rect 3662 16578 3713 16590
rect 3613 16575 3713 16578
rect 3613 16541 3670 16575
rect 3704 16541 3713 16575
rect 3613 16539 3713 16541
rect 3613 16533 3619 16539
rect 3662 16527 3713 16539
rect 3897 16569 3936 16618
rect 3976 16576 4027 16581
rect 3970 16569 3976 16576
rect 3897 16530 3976 16569
rect 3268 16500 3320 16506
rect 3897 16480 3936 16530
rect 3970 16524 3976 16530
rect 4028 16524 4034 16576
rect 4206 16562 4245 16618
rect 4300 16562 4347 16573
rect 4206 16560 4347 16562
rect 4206 16527 4306 16560
rect 3976 16518 4027 16524
rect 4206 16480 4245 16527
rect 4300 16526 4306 16527
rect 4340 16526 4347 16560
rect 4300 16514 4347 16526
rect 2766 16464 2818 16470
rect 2766 16406 2776 16412
rect 2770 16403 2776 16406
rect 2810 16406 2818 16412
rect 2928 16437 2974 16470
rect 2810 16403 2816 16406
rect 2770 16370 2816 16403
rect 2928 16403 2934 16437
rect 2968 16403 2974 16437
rect 2928 16370 2974 16403
rect 3114 16437 3160 16470
rect 3114 16403 3120 16437
rect 3154 16403 3160 16437
rect 3114 16370 3160 16403
rect 3272 16437 3318 16470
rect 3272 16403 3278 16437
rect 3312 16403 3318 16437
rect 3272 16370 3318 16403
rect 3274 16332 3318 16370
rect 2694 16288 3318 16332
rect 3736 16447 3782 16480
rect 3736 16413 3742 16447
rect 3776 16413 3782 16447
rect 3736 16380 3782 16413
rect 3894 16447 3940 16480
rect 3894 16413 3900 16447
rect 3934 16413 3940 16447
rect 4044 16447 4090 16480
rect 4044 16418 4050 16447
rect 3894 16380 3940 16413
rect 4042 16413 4050 16418
rect 4084 16413 4090 16447
rect 4042 16380 4090 16413
rect 4202 16447 4248 16480
rect 4202 16413 4208 16447
rect 4242 16413 4248 16447
rect 4202 16380 4248 16413
rect 3736 16324 3780 16380
rect 4042 16324 4089 16380
rect 1324 16217 1360 16269
rect 1412 16217 1424 16269
rect 1476 16260 1488 16269
rect 1540 16260 1552 16269
rect 1604 16260 1616 16269
rect 1668 16260 1680 16269
rect 1732 16260 1744 16269
rect 1796 16260 1808 16269
rect 1479 16226 1488 16260
rect 1551 16226 1552 16260
rect 1732 16226 1733 16260
rect 1796 16226 1805 16260
rect 1476 16217 1488 16226
rect 1540 16217 1552 16226
rect 1604 16217 1616 16226
rect 1668 16217 1680 16226
rect 1732 16217 1744 16226
rect 1796 16217 1808 16226
rect 1860 16217 1872 16269
rect 1924 16217 1960 16269
rect 3704 16280 4244 16324
rect 3704 16271 3756 16280
rect 3808 16271 3820 16280
rect 1324 16184 1960 16217
rect 2346 16239 2426 16264
rect 2346 16235 3517 16239
rect 2346 16201 2369 16235
rect 2403 16201 3517 16235
rect 2346 16197 3517 16201
rect 2346 16172 2426 16197
rect 2636 16139 2702 16151
rect 272 16085 278 16139
rect 332 16085 2642 16139
rect 2696 16085 2702 16139
rect 2636 16073 2702 16085
rect 3475 16044 3517 16197
rect 3704 16237 3741 16271
rect 3808 16237 3813 16271
rect 3704 16228 3756 16237
rect 3808 16228 3820 16237
rect 3872 16228 3884 16280
rect 3936 16228 3948 16280
rect 4000 16228 4012 16280
rect 4064 16228 4076 16280
rect 4128 16271 4140 16280
rect 4192 16271 4244 16280
rect 4135 16237 4140 16271
rect 4207 16237 4244 16271
rect 4128 16228 4140 16237
rect 4192 16228 4244 16237
rect 3704 16184 4244 16228
rect 3559 16079 3565 16131
rect 3617 16124 3623 16131
rect 4306 16124 4345 16514
rect 4558 16482 4597 16618
rect 4628 16587 4680 16593
rect 4625 16538 4628 16584
rect 4680 16538 4683 16584
rect 4875 16542 4904 16618
rect 4628 16529 4680 16535
rect 4875 16514 4980 16542
rect 4396 16449 4442 16482
rect 4396 16415 4402 16449
rect 4436 16415 4442 16449
rect 4396 16382 4442 16415
rect 4554 16462 4600 16482
rect 4704 16462 4750 16482
rect 4862 16462 4908 16482
rect 4554 16449 4750 16462
rect 4554 16415 4560 16449
rect 4594 16415 4710 16449
rect 4744 16415 4750 16449
rect 4554 16396 4750 16415
rect 4856 16410 4862 16462
rect 4914 16410 4920 16462
rect 4554 16382 4600 16396
rect 4704 16382 4750 16396
rect 4862 16382 4908 16410
rect 4402 16232 4430 16382
rect 4558 16337 4597 16382
rect 4552 16331 4604 16337
rect 4552 16273 4604 16279
rect 4952 16232 4980 16514
rect 5026 16464 5056 16649
rect 5694 16618 5740 16666
rect 5852 16772 5898 16818
rect 5852 16738 5858 16772
rect 5892 16738 5898 16772
rect 5852 16700 5898 16738
rect 5852 16666 5858 16700
rect 5892 16666 5898 16700
rect 5852 16618 5898 16666
rect 6002 16772 6048 16874
rect 6516 16818 6556 17024
rect 6862 17018 6868 17024
rect 6920 17018 6926 17070
rect 6985 17058 7015 17111
rect 6985 17029 7016 17058
rect 6002 16738 6008 16772
rect 6042 16738 6048 16772
rect 6002 16700 6048 16738
rect 6002 16666 6008 16700
rect 6042 16666 6048 16700
rect 6002 16618 6048 16666
rect 6160 16772 6206 16818
rect 6160 16738 6166 16772
rect 6200 16738 6206 16772
rect 6354 16772 6400 16818
rect 6354 16746 6360 16772
rect 6160 16700 6206 16738
rect 6160 16666 6166 16700
rect 6200 16666 6206 16700
rect 6244 16744 6360 16746
rect 6244 16692 6250 16744
rect 6302 16738 6360 16744
rect 6394 16738 6400 16772
rect 6302 16700 6400 16738
rect 6302 16692 6360 16700
rect 6244 16690 6360 16692
rect 6160 16618 6206 16666
rect 6354 16666 6360 16690
rect 6394 16666 6400 16700
rect 6354 16618 6400 16666
rect 6512 16772 6558 16818
rect 6512 16738 6518 16772
rect 6552 16738 6558 16772
rect 6662 16772 6708 16818
rect 6662 16738 6668 16772
rect 6702 16738 6708 16772
rect 6512 16700 6708 16738
rect 6512 16666 6518 16700
rect 6552 16672 6668 16700
rect 6552 16666 6558 16672
rect 6512 16618 6558 16666
rect 6662 16666 6668 16672
rect 6702 16666 6708 16700
rect 6662 16618 6708 16666
rect 6820 16772 6866 16818
rect 6820 16738 6826 16772
rect 6860 16738 6866 16772
rect 6986 16742 7016 17029
rect 6820 16700 6866 16738
rect 6820 16666 6826 16700
rect 6860 16666 6866 16700
rect 6968 16690 6974 16742
rect 7026 16690 7032 16742
rect 6820 16618 6866 16666
rect 6984 16650 7016 16690
rect 5111 16533 5117 16585
rect 5169 16578 5175 16585
rect 5620 16578 5672 16590
rect 5169 16576 5672 16578
rect 5169 16542 5628 16576
rect 5662 16542 5672 16576
rect 5169 16539 5672 16542
rect 5169 16533 5175 16539
rect 5620 16528 5672 16539
rect 5856 16570 5894 16618
rect 5934 16576 5986 16582
rect 5928 16570 5934 16576
rect 5856 16530 5934 16570
rect 5856 16480 5894 16530
rect 5928 16524 5934 16530
rect 5986 16524 5992 16576
rect 6164 16562 6204 16618
rect 6258 16562 6306 16574
rect 6164 16560 6306 16562
rect 6164 16528 6264 16560
rect 5934 16518 5986 16524
rect 6164 16480 6204 16528
rect 6258 16526 6264 16528
rect 6298 16526 6306 16560
rect 6258 16514 6306 16526
rect 5009 16412 5015 16464
rect 5067 16412 5073 16464
rect 5694 16448 5740 16480
rect 5694 16414 5700 16448
rect 5734 16414 5740 16448
rect 4402 16204 4980 16232
rect 3617 16085 4345 16124
rect 3617 16079 3623 16085
rect 5021 16044 5063 16412
rect 5694 16380 5740 16414
rect 5852 16448 5898 16480
rect 5852 16414 5858 16448
rect 5892 16414 5898 16448
rect 6002 16448 6048 16480
rect 6002 16418 6008 16448
rect 5852 16380 5898 16414
rect 6000 16414 6008 16418
rect 6042 16414 6048 16448
rect 5694 16324 5738 16380
rect 6000 16324 6048 16414
rect 6160 16448 6206 16480
rect 6160 16414 6166 16448
rect 6200 16414 6206 16448
rect 6160 16380 6206 16414
rect 5662 16280 6202 16324
rect 5662 16272 5714 16280
rect 5766 16272 5778 16280
rect 5662 16238 5700 16272
rect 5766 16238 5772 16272
rect 5662 16228 5714 16238
rect 5766 16228 5778 16238
rect 5830 16228 5842 16280
rect 5894 16228 5906 16280
rect 5958 16228 5970 16280
rect 6022 16228 6034 16280
rect 6086 16272 6098 16280
rect 6150 16272 6202 16280
rect 6094 16238 6098 16272
rect 6166 16238 6202 16272
rect 6086 16228 6098 16238
rect 6150 16228 6202 16238
rect 5662 16184 6202 16228
rect 5111 16079 5117 16131
rect 5169 16124 5175 16131
rect 6264 16124 6304 16514
rect 6516 16482 6556 16618
rect 6586 16588 6638 16594
rect 6584 16538 6586 16584
rect 6638 16538 6642 16584
rect 6834 16542 6862 16618
rect 6586 16530 6638 16536
rect 6834 16514 6936 16542
rect 6354 16450 6400 16482
rect 6354 16416 6360 16450
rect 6394 16416 6400 16450
rect 6354 16382 6400 16416
rect 6512 16462 6558 16482
rect 6662 16462 6708 16482
rect 6820 16462 6866 16482
rect 6512 16450 6708 16462
rect 6512 16416 6518 16450
rect 6552 16416 6668 16450
rect 6702 16416 6708 16450
rect 6512 16396 6708 16416
rect 6814 16410 6820 16462
rect 6872 16410 6878 16462
rect 6512 16382 6558 16396
rect 6662 16382 6708 16396
rect 6820 16382 6866 16410
rect 6360 16232 6388 16382
rect 6516 16338 6556 16382
rect 6510 16332 6562 16338
rect 6510 16274 6562 16280
rect 6908 16232 6936 16514
rect 6984 16464 7014 16650
rect 6968 16412 6974 16464
rect 7026 16412 7032 16464
rect 6360 16204 6936 16232
rect 6908 16140 6936 16204
rect 5169 16086 6304 16124
rect 6346 16112 6936 16140
rect 5169 16085 5572 16086
rect 5169 16079 5175 16085
rect 3475 16002 5063 16044
rect 5035 15961 5087 15967
rect 3472 15877 4907 15916
rect 6346 15949 6374 16112
rect 6908 16110 6936 16112
rect 5087 15921 6374 15949
rect 6968 15910 6974 15962
rect 7026 15910 7032 15962
rect 5035 15903 5087 15909
rect 1348 15743 1880 15786
rect 1348 15734 1398 15743
rect 1450 15734 1462 15743
rect 1348 15700 1383 15734
rect 1450 15700 1455 15734
rect 1348 15691 1398 15700
rect 1450 15691 1462 15700
rect 1514 15691 1526 15743
rect 1578 15691 1590 15743
rect 1642 15691 1654 15743
rect 1706 15691 1718 15743
rect 1770 15734 1782 15743
rect 1834 15734 1880 15743
rect 1777 15700 1782 15734
rect 1849 15700 1880 15734
rect 3472 15719 3511 15877
rect 4738 15835 4744 15842
rect 4558 15796 4744 15835
rect 1770 15691 1782 15700
rect 1834 15691 1880 15700
rect 550 15672 622 15676
rect 550 15620 560 15672
rect 612 15620 622 15672
rect 696 15670 768 15676
rect 550 15608 566 15620
rect 607 15608 622 15620
rect 682 15668 768 15670
rect 682 15616 702 15668
rect 754 15616 768 15668
rect 682 15614 710 15616
rect 550 15578 622 15608
rect 696 15608 710 15614
rect 751 15608 768 15616
rect 696 15578 768 15608
rect 840 15653 912 15682
rect 840 15613 856 15653
rect 897 15613 912 15653
rect 840 15584 912 15613
rect 994 15653 1066 15682
rect 994 15613 1009 15653
rect 1050 15613 1066 15653
rect 1348 15646 1880 15691
rect 994 15584 1066 15613
rect 564 15538 608 15578
rect 856 15518 900 15584
rect 378 15510 433 15516
rect 846 15466 852 15518
rect 904 15466 910 15518
rect 378 15225 433 15455
rect 856 15426 900 15466
rect 1008 15426 1052 15584
rect 1407 15580 1448 15646
rect 1693 15580 1735 15646
rect 1941 15643 2687 15688
rect 1404 15533 1450 15580
rect 1404 15499 1410 15533
rect 1444 15499 1450 15533
rect 1404 15461 1450 15499
rect 1404 15427 1410 15461
rect 1444 15427 1450 15461
rect 708 15382 900 15426
rect 372 15170 378 15225
rect 433 15170 439 15225
rect 708 15148 752 15382
rect 998 15374 1004 15426
rect 1056 15374 1062 15426
rect 1404 15380 1450 15427
rect 1562 15533 1608 15580
rect 1562 15499 1568 15533
rect 1602 15499 1608 15533
rect 1562 15461 1608 15499
rect 1562 15427 1568 15461
rect 1602 15427 1608 15461
rect 1562 15380 1608 15427
rect 1692 15533 1738 15580
rect 1692 15499 1698 15533
rect 1732 15499 1738 15533
rect 1692 15461 1738 15499
rect 1692 15427 1698 15461
rect 1732 15427 1738 15461
rect 1692 15380 1738 15427
rect 1850 15577 1896 15580
rect 1941 15577 1986 15643
rect 1850 15533 1986 15577
rect 1850 15499 1856 15533
rect 1890 15532 1986 15533
rect 2024 15533 2070 15580
rect 1890 15499 1896 15532
rect 1850 15461 1896 15499
rect 2024 15499 2030 15533
rect 2064 15499 2070 15533
rect 2024 15464 2070 15499
rect 1998 15462 2070 15464
rect 1850 15427 1856 15461
rect 1890 15427 1896 15461
rect 1850 15380 1896 15427
rect 1928 15461 2070 15462
rect 1928 15437 2030 15461
rect 1928 15420 1935 15437
rect 1929 15385 1935 15420
rect 1987 15427 2030 15437
rect 2064 15427 2070 15461
rect 1987 15420 2070 15427
rect 1987 15385 1993 15420
rect 2024 15380 2070 15420
rect 2182 15536 2228 15580
rect 2366 15536 2412 15580
rect 2182 15533 2412 15536
rect 2182 15499 2188 15533
rect 2222 15499 2372 15533
rect 2406 15499 2412 15533
rect 2182 15461 2412 15499
rect 2182 15427 2188 15461
rect 2222 15427 2372 15461
rect 2406 15427 2412 15461
rect 2182 15410 2412 15427
rect 2182 15380 2228 15410
rect 2366 15380 2412 15410
rect 2524 15533 2570 15580
rect 2524 15499 2530 15533
rect 2564 15499 2570 15533
rect 2642 15509 2687 15643
rect 3118 15680 3511 15719
rect 3724 15742 4264 15786
rect 3724 15690 3776 15742
rect 3828 15733 3840 15742
rect 3892 15733 3904 15742
rect 3956 15733 3968 15742
rect 4020 15733 4032 15742
rect 4084 15733 4096 15742
rect 4148 15733 4160 15742
rect 3831 15699 3840 15733
rect 3903 15699 3904 15733
rect 4084 15699 4085 15733
rect 4148 15699 4157 15733
rect 3828 15690 3840 15699
rect 3892 15690 3904 15699
rect 3956 15690 3968 15699
rect 4020 15690 4032 15699
rect 4084 15690 4096 15699
rect 4148 15690 4160 15699
rect 4212 15690 4264 15742
rect 2774 15636 2816 15637
rect 2758 15628 2816 15636
rect 2758 15576 2769 15628
rect 2821 15576 2827 15628
rect 3118 15580 3157 15680
rect 3724 15646 4264 15690
rect 3741 15590 3787 15646
rect 3736 15589 3787 15590
rect 2758 15533 2816 15576
rect 2524 15461 2570 15499
rect 2524 15427 2530 15461
rect 2564 15427 2570 15461
rect 2524 15420 2570 15427
rect 2613 15481 2715 15509
rect 2613 15447 2647 15481
rect 2681 15447 2715 15481
rect 2524 15380 2574 15420
rect 2613 15419 2715 15447
rect 2758 15499 2776 15533
rect 2810 15499 2816 15533
rect 2758 15461 2816 15499
rect 2758 15427 2776 15461
rect 2810 15427 2816 15461
rect 1008 15320 1052 15374
rect 1245 15339 1328 15358
rect 852 15276 1052 15320
rect 1148 15337 1328 15339
rect 1148 15285 1155 15337
rect 1207 15327 1328 15337
rect 1207 15293 1269 15327
rect 1303 15293 1328 15327
rect 1207 15285 1328 15293
rect 1148 15284 1328 15285
rect 852 15154 896 15276
rect 1245 15263 1328 15284
rect 1568 15346 1602 15380
rect 1568 15336 1820 15346
rect 1568 15284 1758 15336
rect 1810 15284 1820 15336
rect 1568 15274 1820 15284
rect 1568 15242 1608 15274
rect 1853 15242 1892 15380
rect 2185 15242 2224 15380
rect 2255 15343 2325 15349
rect 2255 15334 2331 15343
rect 2255 15282 2270 15334
rect 2322 15282 2331 15334
rect 2255 15273 2331 15282
rect 2255 15267 2325 15273
rect 2368 15242 2407 15380
rect 2530 15346 2574 15380
rect 2758 15380 2816 15427
rect 2928 15533 2974 15580
rect 2928 15499 2934 15533
rect 2968 15520 2974 15533
rect 3114 15533 3160 15580
rect 3114 15520 3120 15533
rect 2968 15499 3120 15520
rect 3154 15499 3160 15533
rect 3272 15533 3318 15580
rect 3272 15523 3278 15533
rect 3312 15523 3318 15533
rect 3736 15543 3782 15589
rect 2928 15461 3160 15499
rect 3262 15471 3268 15523
rect 3320 15471 3326 15523
rect 3736 15509 3742 15543
rect 3776 15509 3782 15543
rect 3736 15471 3782 15509
rect 2928 15427 2934 15461
rect 2968 15427 3120 15461
rect 3154 15427 3160 15461
rect 2928 15410 3160 15427
rect 2928 15380 2974 15410
rect 3114 15380 3160 15410
rect 3272 15461 3318 15471
rect 3272 15427 3278 15461
rect 3312 15427 3318 15461
rect 3272 15380 3318 15427
rect 3736 15437 3742 15471
rect 3776 15437 3782 15471
rect 3736 15390 3782 15437
rect 3894 15543 3940 15590
rect 3894 15509 3900 15543
rect 3934 15509 3940 15543
rect 3894 15471 3940 15509
rect 3894 15437 3900 15471
rect 3934 15437 3940 15471
rect 3894 15390 3940 15437
rect 4044 15543 4090 15646
rect 4558 15590 4597 15796
rect 4738 15790 4744 15796
rect 4796 15790 4802 15842
rect 4868 15590 4907 15877
rect 5682 15742 6222 15786
rect 5682 15690 5734 15742
rect 5786 15732 5798 15742
rect 5850 15732 5862 15742
rect 5914 15732 5926 15742
rect 5978 15732 5990 15742
rect 6042 15732 6054 15742
rect 6106 15732 6118 15742
rect 5790 15698 5798 15732
rect 6042 15698 6044 15732
rect 6106 15698 6116 15732
rect 5786 15690 5798 15698
rect 5850 15690 5862 15698
rect 5914 15690 5926 15698
rect 5978 15690 5990 15698
rect 6042 15690 6054 15698
rect 6106 15690 6118 15698
rect 6170 15690 6222 15742
rect 5682 15646 6222 15690
rect 5700 15590 5746 15646
rect 4044 15509 4050 15543
rect 4084 15509 4090 15543
rect 4044 15471 4090 15509
rect 4044 15437 4050 15471
rect 4084 15437 4090 15471
rect 4044 15390 4090 15437
rect 4202 15543 4248 15590
rect 4202 15509 4208 15543
rect 4242 15509 4248 15543
rect 4396 15543 4442 15590
rect 4396 15517 4402 15543
rect 4202 15471 4248 15509
rect 4202 15437 4208 15471
rect 4242 15437 4248 15471
rect 4285 15515 4402 15517
rect 4285 15463 4292 15515
rect 4344 15509 4402 15515
rect 4436 15509 4442 15543
rect 4344 15471 4442 15509
rect 4344 15463 4402 15471
rect 4285 15462 4402 15463
rect 4202 15390 4248 15437
rect 4396 15437 4402 15462
rect 4436 15437 4442 15471
rect 4396 15390 4442 15437
rect 4554 15543 4600 15590
rect 4554 15509 4560 15543
rect 4594 15510 4600 15543
rect 4704 15543 4750 15590
rect 4704 15510 4710 15543
rect 4594 15509 4710 15510
rect 4744 15509 4750 15543
rect 4554 15471 4750 15509
rect 4554 15437 4560 15471
rect 4594 15444 4710 15471
rect 4594 15437 4600 15444
rect 4554 15390 4600 15437
rect 4704 15437 4710 15444
rect 4744 15437 4750 15471
rect 4704 15390 4750 15437
rect 4862 15543 4908 15590
rect 4862 15509 4868 15543
rect 4902 15509 4908 15543
rect 5694 15544 5740 15590
rect 5027 15514 5057 15523
rect 4862 15471 4908 15509
rect 4862 15437 4868 15471
rect 4902 15437 4908 15471
rect 5010 15462 5016 15514
rect 5068 15462 5074 15514
rect 5694 15510 5700 15544
rect 5734 15510 5740 15544
rect 5694 15472 5740 15510
rect 4862 15390 4908 15437
rect 5026 15421 5057 15462
rect 5694 15438 5700 15472
rect 5734 15438 5740 15472
rect 2758 15346 2802 15380
rect 2530 15302 2656 15346
rect 1242 15222 1248 15226
rect 1138 15178 1248 15222
rect 1138 15154 1182 15178
rect 1242 15174 1248 15178
rect 1300 15174 1306 15226
rect 1404 15209 1450 15242
rect 1404 15175 1410 15209
rect 1444 15175 1450 15209
rect 1404 15171 1450 15175
rect 378 15126 434 15132
rect 550 15126 622 15148
rect 434 15120 622 15126
rect 434 15080 565 15120
rect 606 15080 622 15120
rect 434 15070 622 15080
rect 378 15064 434 15070
rect 550 15050 622 15070
rect 696 15120 768 15148
rect 696 15080 712 15120
rect 753 15080 768 15120
rect 696 15050 768 15080
rect 840 15125 912 15154
rect 840 15085 856 15125
rect 897 15085 912 15125
rect 840 15056 912 15085
rect 994 15126 1182 15154
rect 994 15086 1010 15126
rect 1051 15110 1182 15126
rect 1399 15142 1450 15171
rect 1562 15209 1608 15242
rect 1562 15175 1568 15209
rect 1602 15175 1608 15209
rect 1692 15209 1738 15242
rect 1692 15180 1698 15209
rect 1562 15142 1608 15175
rect 1690 15175 1698 15180
rect 1732 15180 1738 15209
rect 1850 15209 1896 15242
rect 2024 15226 2070 15242
rect 1732 15175 1740 15180
rect 1051 15086 1066 15110
rect 1399 15096 1449 15142
rect 1690 15096 1740 15175
rect 1850 15175 1856 15209
rect 1890 15175 1896 15209
rect 1850 15142 1896 15175
rect 2014 15174 2020 15226
rect 2072 15174 2078 15226
rect 2182 15209 2228 15242
rect 2182 15175 2188 15209
rect 2222 15175 2228 15209
rect 2024 15142 2070 15174
rect 2182 15142 2228 15175
rect 2366 15209 2412 15242
rect 2524 15224 2570 15242
rect 2366 15175 2372 15209
rect 2406 15175 2412 15209
rect 2366 15142 2412 15175
rect 2516 15172 2522 15224
rect 2574 15172 2580 15224
rect 2524 15142 2570 15172
rect 2024 15110 2068 15142
rect 2612 15110 2656 15302
rect 994 15056 1066 15086
rect 1324 15041 1960 15096
rect 2024 15066 2656 15110
rect 2694 15302 2802 15346
rect 2832 15332 2904 15342
rect 2694 15104 2738 15302
rect 2832 15280 2842 15332
rect 2894 15280 2904 15332
rect 2832 15270 2904 15280
rect 2933 15242 2972 15380
rect 3118 15242 3157 15380
rect 3272 15336 3316 15380
rect 3268 15330 3320 15336
rect 3555 15305 3561 15357
rect 3613 15350 3619 15357
rect 3662 15350 3713 15362
rect 3613 15347 3713 15350
rect 3613 15313 3670 15347
rect 3704 15313 3713 15347
rect 3613 15311 3713 15313
rect 3613 15305 3619 15311
rect 3662 15299 3713 15311
rect 3897 15341 3936 15390
rect 3976 15348 4027 15353
rect 3970 15341 3976 15348
rect 3897 15302 3976 15341
rect 3268 15272 3320 15278
rect 3897 15252 3936 15302
rect 3970 15296 3976 15302
rect 4028 15296 4034 15348
rect 4206 15334 4245 15390
rect 4300 15334 4347 15345
rect 4206 15332 4347 15334
rect 4206 15299 4306 15332
rect 3976 15290 4027 15296
rect 4206 15252 4245 15299
rect 4300 15298 4306 15299
rect 4340 15298 4347 15332
rect 4300 15286 4347 15298
rect 2766 15236 2818 15242
rect 2766 15178 2776 15184
rect 2770 15175 2776 15178
rect 2810 15178 2818 15184
rect 2928 15209 2974 15242
rect 2810 15175 2816 15178
rect 2770 15142 2816 15175
rect 2928 15175 2934 15209
rect 2968 15175 2974 15209
rect 2928 15142 2974 15175
rect 3114 15209 3160 15242
rect 3114 15175 3120 15209
rect 3154 15175 3160 15209
rect 3114 15142 3160 15175
rect 3272 15209 3318 15242
rect 3272 15175 3278 15209
rect 3312 15175 3318 15209
rect 3272 15142 3318 15175
rect 3274 15104 3318 15142
rect 2694 15060 3318 15104
rect 3736 15219 3782 15252
rect 3736 15185 3742 15219
rect 3776 15185 3782 15219
rect 3736 15152 3782 15185
rect 3894 15219 3940 15252
rect 3894 15185 3900 15219
rect 3934 15185 3940 15219
rect 4044 15219 4090 15252
rect 4044 15190 4050 15219
rect 3894 15152 3940 15185
rect 4042 15185 4050 15190
rect 4084 15185 4090 15219
rect 4042 15152 4090 15185
rect 4202 15219 4248 15252
rect 4202 15185 4208 15219
rect 4242 15185 4248 15219
rect 4202 15152 4248 15185
rect 3736 15096 3780 15152
rect 4042 15096 4089 15152
rect 1324 14989 1360 15041
rect 1412 14989 1424 15041
rect 1476 15032 1488 15041
rect 1540 15032 1552 15041
rect 1604 15032 1616 15041
rect 1668 15032 1680 15041
rect 1732 15032 1744 15041
rect 1796 15032 1808 15041
rect 1479 14998 1488 15032
rect 1551 14998 1552 15032
rect 1732 14998 1733 15032
rect 1796 14998 1805 15032
rect 1476 14989 1488 14998
rect 1540 14989 1552 14998
rect 1604 14989 1616 14998
rect 1668 14989 1680 14998
rect 1732 14989 1744 14998
rect 1796 14989 1808 14998
rect 1860 14989 1872 15041
rect 1924 14989 1960 15041
rect 3704 15052 4244 15096
rect 3704 15043 3756 15052
rect 3808 15043 3820 15052
rect 1324 14956 1960 14989
rect 2346 15011 2426 15036
rect 2346 15007 3517 15011
rect 2346 14973 2369 15007
rect 2403 14973 3517 15007
rect 2346 14969 3517 14973
rect 2346 14944 2426 14969
rect 2636 14911 2702 14923
rect 272 14857 278 14911
rect 332 14857 2642 14911
rect 2696 14857 2702 14911
rect 2636 14845 2702 14857
rect 3475 14816 3517 14969
rect 3704 15009 3741 15043
rect 3808 15009 3813 15043
rect 3704 15000 3756 15009
rect 3808 15000 3820 15009
rect 3872 15000 3884 15052
rect 3936 15000 3948 15052
rect 4000 15000 4012 15052
rect 4064 15000 4076 15052
rect 4128 15043 4140 15052
rect 4192 15043 4244 15052
rect 4135 15009 4140 15043
rect 4207 15009 4244 15043
rect 4128 15000 4140 15009
rect 4192 15000 4244 15009
rect 3704 14956 4244 15000
rect 3559 14851 3565 14903
rect 3617 14896 3623 14903
rect 4306 14896 4345 15286
rect 4558 15254 4597 15390
rect 4628 15359 4680 15365
rect 4625 15310 4628 15356
rect 4680 15310 4683 15356
rect 4875 15314 4904 15390
rect 4628 15301 4680 15307
rect 4875 15286 4980 15314
rect 4396 15221 4442 15254
rect 4396 15187 4402 15221
rect 4436 15187 4442 15221
rect 4396 15154 4442 15187
rect 4554 15234 4600 15254
rect 4704 15234 4750 15254
rect 4862 15234 4908 15254
rect 4554 15221 4750 15234
rect 4554 15187 4560 15221
rect 4594 15187 4710 15221
rect 4744 15187 4750 15221
rect 4554 15168 4750 15187
rect 4856 15182 4862 15234
rect 4914 15182 4920 15234
rect 4554 15154 4600 15168
rect 4704 15154 4750 15168
rect 4862 15154 4908 15182
rect 4402 15004 4430 15154
rect 4558 15109 4597 15154
rect 4552 15103 4604 15109
rect 4552 15045 4604 15051
rect 4952 15004 4980 15286
rect 5026 15236 5056 15421
rect 5694 15390 5740 15438
rect 5852 15544 5898 15590
rect 5852 15510 5858 15544
rect 5892 15510 5898 15544
rect 5852 15472 5898 15510
rect 5852 15438 5858 15472
rect 5892 15438 5898 15472
rect 5852 15390 5898 15438
rect 6002 15544 6048 15646
rect 6516 15590 6556 15834
rect 6985 15830 7015 15910
rect 6985 15801 7016 15830
rect 6002 15510 6008 15544
rect 6042 15510 6048 15544
rect 6002 15472 6048 15510
rect 6002 15438 6008 15472
rect 6042 15438 6048 15472
rect 6002 15390 6048 15438
rect 6160 15544 6206 15590
rect 6160 15510 6166 15544
rect 6200 15510 6206 15544
rect 6354 15544 6400 15590
rect 6354 15518 6360 15544
rect 6160 15472 6206 15510
rect 6160 15438 6166 15472
rect 6200 15438 6206 15472
rect 6244 15516 6360 15518
rect 6244 15464 6250 15516
rect 6302 15510 6360 15516
rect 6394 15510 6400 15544
rect 6302 15472 6400 15510
rect 6302 15464 6360 15472
rect 6244 15462 6360 15464
rect 6160 15390 6206 15438
rect 6354 15438 6360 15462
rect 6394 15438 6400 15472
rect 6354 15390 6400 15438
rect 6512 15544 6558 15590
rect 6512 15510 6518 15544
rect 6552 15510 6558 15544
rect 6662 15544 6708 15590
rect 6662 15510 6668 15544
rect 6702 15510 6708 15544
rect 6512 15472 6708 15510
rect 6512 15438 6518 15472
rect 6552 15444 6668 15472
rect 6552 15438 6558 15444
rect 6512 15390 6558 15438
rect 6662 15438 6668 15444
rect 6702 15438 6708 15472
rect 6662 15390 6708 15438
rect 6820 15544 6866 15590
rect 6820 15510 6826 15544
rect 6860 15510 6866 15544
rect 6986 15514 7016 15801
rect 6820 15472 6866 15510
rect 6820 15438 6826 15472
rect 6860 15438 6866 15472
rect 6968 15462 6974 15514
rect 7026 15462 7032 15514
rect 6820 15390 6866 15438
rect 6984 15422 7016 15462
rect 5273 15305 5279 15357
rect 5331 15350 5337 15357
rect 5620 15350 5672 15362
rect 5331 15348 5672 15350
rect 5331 15314 5628 15348
rect 5662 15314 5672 15348
rect 5331 15311 5672 15314
rect 5331 15305 5337 15311
rect 5620 15300 5672 15311
rect 5856 15342 5894 15390
rect 5934 15348 5986 15354
rect 5928 15342 5934 15348
rect 5856 15302 5934 15342
rect 5856 15252 5894 15302
rect 5928 15296 5934 15302
rect 5986 15296 5992 15348
rect 6164 15334 6204 15390
rect 6258 15334 6306 15346
rect 6164 15332 6306 15334
rect 6164 15300 6264 15332
rect 5934 15290 5986 15296
rect 6164 15252 6204 15300
rect 6258 15298 6264 15300
rect 6298 15298 6306 15332
rect 6258 15286 6306 15298
rect 5009 15184 5015 15236
rect 5067 15184 5073 15236
rect 5694 15220 5740 15252
rect 5694 15186 5700 15220
rect 5734 15186 5740 15220
rect 4402 14976 4980 15004
rect 3617 14857 4345 14896
rect 3617 14851 3623 14857
rect 5021 14816 5063 15184
rect 5694 15152 5740 15186
rect 5852 15220 5898 15252
rect 5852 15186 5858 15220
rect 5892 15186 5898 15220
rect 6002 15220 6048 15252
rect 6002 15190 6008 15220
rect 5852 15152 5898 15186
rect 6000 15186 6008 15190
rect 6042 15186 6048 15220
rect 5694 15096 5738 15152
rect 6000 15096 6048 15186
rect 6160 15220 6206 15252
rect 6160 15186 6166 15220
rect 6200 15186 6206 15220
rect 6160 15152 6206 15186
rect 5662 15052 6202 15096
rect 5662 15044 5714 15052
rect 5766 15044 5778 15052
rect 5662 15010 5700 15044
rect 5766 15010 5772 15044
rect 5662 15000 5714 15010
rect 5766 15000 5778 15010
rect 5830 15000 5842 15052
rect 5894 15000 5906 15052
rect 5958 15000 5970 15052
rect 6022 15000 6034 15052
rect 6086 15044 6098 15052
rect 6150 15044 6202 15052
rect 6094 15010 6098 15044
rect 6166 15010 6202 15044
rect 6086 15000 6098 15010
rect 6150 15000 6202 15010
rect 5662 14956 6202 15000
rect 5273 14851 5279 14903
rect 5331 14896 5337 14903
rect 6264 14896 6304 15286
rect 6516 15254 6556 15390
rect 6586 15360 6638 15366
rect 6584 15310 6586 15356
rect 6638 15310 6642 15356
rect 6834 15314 6862 15390
rect 6586 15302 6638 15308
rect 6834 15286 6936 15314
rect 6354 15222 6400 15254
rect 6354 15188 6360 15222
rect 6394 15188 6400 15222
rect 6354 15154 6400 15188
rect 6512 15234 6558 15254
rect 6662 15234 6708 15254
rect 6820 15234 6866 15254
rect 6512 15222 6708 15234
rect 6512 15188 6518 15222
rect 6552 15188 6668 15222
rect 6702 15188 6708 15222
rect 6512 15168 6708 15188
rect 6814 15182 6820 15234
rect 6872 15182 6878 15234
rect 6512 15154 6558 15168
rect 6662 15154 6708 15168
rect 6820 15154 6866 15182
rect 6360 15004 6388 15154
rect 6516 15110 6556 15154
rect 6510 15104 6562 15110
rect 6510 15046 6562 15052
rect 6908 15004 6936 15286
rect 6984 15236 7014 15422
rect 6968 15184 6974 15236
rect 7026 15184 7032 15236
rect 6360 14976 6936 15004
rect 5331 14858 6304 14896
rect 5331 14857 5584 14858
rect 5331 14851 5337 14857
rect 3475 14774 5063 14816
rect 6908 14788 6936 14976
rect 6908 14760 7234 14788
rect 5029 14696 5081 14702
rect 3472 14649 4907 14688
rect 1348 14515 1880 14558
rect 1348 14506 1398 14515
rect 1450 14506 1462 14515
rect 1348 14472 1383 14506
rect 1450 14472 1455 14506
rect 1348 14463 1398 14472
rect 1450 14463 1462 14472
rect 1514 14463 1526 14515
rect 1578 14463 1590 14515
rect 1642 14463 1654 14515
rect 1706 14463 1718 14515
rect 1770 14506 1782 14515
rect 1834 14506 1880 14515
rect 1777 14472 1782 14506
rect 1849 14472 1880 14506
rect 3472 14491 3511 14649
rect 4738 14607 4744 14614
rect 4558 14568 4744 14607
rect 1770 14463 1782 14472
rect 1834 14463 1880 14472
rect 550 14444 622 14448
rect 550 14392 560 14444
rect 612 14392 622 14444
rect 696 14442 768 14448
rect 550 14380 566 14392
rect 607 14380 622 14392
rect 682 14440 768 14442
rect 682 14388 702 14440
rect 754 14388 768 14440
rect 682 14386 710 14388
rect 550 14350 622 14380
rect 696 14380 710 14386
rect 751 14380 768 14388
rect 696 14350 768 14380
rect 840 14425 912 14454
rect 840 14385 856 14425
rect 897 14385 912 14425
rect 840 14356 912 14385
rect 994 14425 1066 14454
rect 994 14385 1009 14425
rect 1050 14385 1066 14425
rect 1348 14418 1880 14463
rect 994 14356 1066 14385
rect 564 14310 608 14350
rect 856 14290 900 14356
rect 378 14282 433 14288
rect 846 14238 852 14290
rect 904 14238 910 14290
rect 378 13997 433 14227
rect 856 14198 900 14238
rect 1008 14198 1052 14356
rect 1407 14352 1448 14418
rect 1693 14352 1735 14418
rect 1941 14415 2687 14460
rect 1404 14305 1450 14352
rect 1404 14271 1410 14305
rect 1444 14271 1450 14305
rect 1404 14233 1450 14271
rect 1404 14199 1410 14233
rect 1444 14199 1450 14233
rect 708 14154 900 14198
rect 372 13942 378 13997
rect 433 13942 439 13997
rect 708 13920 752 14154
rect 998 14146 1004 14198
rect 1056 14146 1062 14198
rect 1404 14152 1450 14199
rect 1562 14305 1608 14352
rect 1562 14271 1568 14305
rect 1602 14271 1608 14305
rect 1562 14233 1608 14271
rect 1562 14199 1568 14233
rect 1602 14199 1608 14233
rect 1562 14152 1608 14199
rect 1692 14305 1738 14352
rect 1692 14271 1698 14305
rect 1732 14271 1738 14305
rect 1692 14233 1738 14271
rect 1692 14199 1698 14233
rect 1732 14199 1738 14233
rect 1692 14152 1738 14199
rect 1850 14349 1896 14352
rect 1941 14349 1986 14415
rect 1850 14305 1986 14349
rect 1850 14271 1856 14305
rect 1890 14304 1986 14305
rect 2024 14305 2070 14352
rect 1890 14271 1896 14304
rect 1850 14233 1896 14271
rect 2024 14271 2030 14305
rect 2064 14271 2070 14305
rect 2024 14236 2070 14271
rect 1998 14234 2070 14236
rect 1850 14199 1856 14233
rect 1890 14199 1896 14233
rect 1850 14152 1896 14199
rect 1928 14233 2070 14234
rect 1928 14209 2030 14233
rect 1928 14192 1935 14209
rect 1929 14157 1935 14192
rect 1987 14199 2030 14209
rect 2064 14199 2070 14233
rect 1987 14192 2070 14199
rect 1987 14157 1993 14192
rect 2024 14152 2070 14192
rect 2182 14308 2228 14352
rect 2366 14308 2412 14352
rect 2182 14305 2412 14308
rect 2182 14271 2188 14305
rect 2222 14271 2372 14305
rect 2406 14271 2412 14305
rect 2182 14233 2412 14271
rect 2182 14199 2188 14233
rect 2222 14199 2372 14233
rect 2406 14199 2412 14233
rect 2182 14182 2412 14199
rect 2182 14152 2228 14182
rect 2366 14152 2412 14182
rect 2524 14305 2570 14352
rect 2524 14271 2530 14305
rect 2564 14271 2570 14305
rect 2642 14281 2687 14415
rect 3118 14452 3511 14491
rect 3724 14514 4264 14558
rect 3724 14462 3776 14514
rect 3828 14505 3840 14514
rect 3892 14505 3904 14514
rect 3956 14505 3968 14514
rect 4020 14505 4032 14514
rect 4084 14505 4096 14514
rect 4148 14505 4160 14514
rect 3831 14471 3840 14505
rect 3903 14471 3904 14505
rect 4084 14471 4085 14505
rect 4148 14471 4157 14505
rect 3828 14462 3840 14471
rect 3892 14462 3904 14471
rect 3956 14462 3968 14471
rect 4020 14462 4032 14471
rect 4084 14462 4096 14471
rect 4148 14462 4160 14471
rect 4212 14462 4264 14514
rect 2774 14408 2816 14409
rect 2758 14400 2816 14408
rect 2758 14348 2769 14400
rect 2821 14348 2827 14400
rect 3118 14352 3157 14452
rect 3724 14418 4264 14462
rect 3741 14362 3787 14418
rect 3736 14361 3787 14362
rect 2758 14305 2816 14348
rect 2524 14233 2570 14271
rect 2524 14199 2530 14233
rect 2564 14199 2570 14233
rect 2524 14192 2570 14199
rect 2613 14253 2715 14281
rect 2613 14219 2647 14253
rect 2681 14219 2715 14253
rect 2524 14152 2574 14192
rect 2613 14191 2715 14219
rect 2758 14271 2776 14305
rect 2810 14271 2816 14305
rect 2758 14233 2816 14271
rect 2758 14199 2776 14233
rect 2810 14199 2816 14233
rect 1008 14092 1052 14146
rect 1245 14111 1328 14130
rect 852 14048 1052 14092
rect 1148 14109 1328 14111
rect 1148 14057 1155 14109
rect 1207 14099 1328 14109
rect 1207 14065 1269 14099
rect 1303 14065 1328 14099
rect 1207 14057 1328 14065
rect 1148 14056 1328 14057
rect 852 13926 896 14048
rect 1245 14035 1328 14056
rect 1568 14118 1602 14152
rect 1568 14108 1820 14118
rect 1568 14056 1758 14108
rect 1810 14056 1820 14108
rect 1568 14046 1820 14056
rect 1568 14014 1608 14046
rect 1853 14014 1892 14152
rect 2185 14014 2224 14152
rect 2255 14115 2325 14121
rect 2255 14106 2331 14115
rect 2255 14054 2270 14106
rect 2322 14054 2331 14106
rect 2255 14045 2331 14054
rect 2255 14039 2325 14045
rect 2368 14014 2407 14152
rect 2530 14118 2574 14152
rect 2758 14152 2816 14199
rect 2928 14305 2974 14352
rect 2928 14271 2934 14305
rect 2968 14292 2974 14305
rect 3114 14305 3160 14352
rect 3114 14292 3120 14305
rect 2968 14271 3120 14292
rect 3154 14271 3160 14305
rect 3272 14305 3318 14352
rect 3272 14295 3278 14305
rect 3312 14295 3318 14305
rect 3736 14315 3782 14361
rect 2928 14233 3160 14271
rect 3262 14243 3268 14295
rect 3320 14243 3326 14295
rect 3736 14281 3742 14315
rect 3776 14281 3782 14315
rect 3736 14243 3782 14281
rect 2928 14199 2934 14233
rect 2968 14199 3120 14233
rect 3154 14199 3160 14233
rect 2928 14182 3160 14199
rect 2928 14152 2974 14182
rect 3114 14152 3160 14182
rect 3272 14233 3318 14243
rect 3272 14199 3278 14233
rect 3312 14199 3318 14233
rect 3272 14152 3318 14199
rect 3736 14209 3742 14243
rect 3776 14209 3782 14243
rect 3736 14162 3782 14209
rect 3894 14315 3940 14362
rect 3894 14281 3900 14315
rect 3934 14281 3940 14315
rect 3894 14243 3940 14281
rect 3894 14209 3900 14243
rect 3934 14209 3940 14243
rect 3894 14162 3940 14209
rect 4044 14315 4090 14418
rect 4558 14362 4597 14568
rect 4738 14562 4744 14568
rect 4796 14562 4802 14614
rect 4868 14362 4907 14649
rect 5081 14655 7015 14685
rect 5029 14638 5081 14644
rect 6862 14607 6868 14614
rect 6516 14568 6868 14607
rect 5682 14514 6222 14558
rect 5682 14462 5734 14514
rect 5786 14504 5798 14514
rect 5850 14504 5862 14514
rect 5914 14504 5926 14514
rect 5978 14504 5990 14514
rect 6042 14504 6054 14514
rect 6106 14504 6118 14514
rect 5790 14470 5798 14504
rect 6042 14470 6044 14504
rect 6106 14470 6116 14504
rect 5786 14462 5798 14470
rect 5850 14462 5862 14470
rect 5914 14462 5926 14470
rect 5978 14462 5990 14470
rect 6042 14462 6054 14470
rect 6106 14462 6118 14470
rect 6170 14462 6222 14514
rect 5682 14418 6222 14462
rect 5700 14362 5746 14418
rect 4044 14281 4050 14315
rect 4084 14281 4090 14315
rect 4044 14243 4090 14281
rect 4044 14209 4050 14243
rect 4084 14209 4090 14243
rect 4044 14162 4090 14209
rect 4202 14315 4248 14362
rect 4202 14281 4208 14315
rect 4242 14281 4248 14315
rect 4396 14315 4442 14362
rect 4396 14289 4402 14315
rect 4202 14243 4248 14281
rect 4202 14209 4208 14243
rect 4242 14209 4248 14243
rect 4285 14287 4402 14289
rect 4285 14235 4292 14287
rect 4344 14281 4402 14287
rect 4436 14281 4442 14315
rect 4344 14243 4442 14281
rect 4344 14235 4402 14243
rect 4285 14234 4402 14235
rect 4202 14162 4248 14209
rect 4396 14209 4402 14234
rect 4436 14209 4442 14243
rect 4396 14162 4442 14209
rect 4554 14315 4600 14362
rect 4554 14281 4560 14315
rect 4594 14282 4600 14315
rect 4704 14315 4750 14362
rect 4704 14282 4710 14315
rect 4594 14281 4710 14282
rect 4744 14281 4750 14315
rect 4554 14243 4750 14281
rect 4554 14209 4560 14243
rect 4594 14216 4710 14243
rect 4594 14209 4600 14216
rect 4554 14162 4600 14209
rect 4704 14209 4710 14216
rect 4744 14209 4750 14243
rect 4704 14162 4750 14209
rect 4862 14315 4908 14362
rect 4862 14281 4868 14315
rect 4902 14281 4908 14315
rect 5694 14316 5740 14362
rect 5027 14286 5057 14295
rect 4862 14243 4908 14281
rect 4862 14209 4868 14243
rect 4902 14209 4908 14243
rect 5010 14234 5016 14286
rect 5068 14234 5074 14286
rect 5694 14282 5700 14316
rect 5734 14282 5740 14316
rect 5694 14244 5740 14282
rect 4862 14162 4908 14209
rect 5026 14193 5057 14234
rect 5694 14210 5700 14244
rect 5734 14210 5740 14244
rect 2758 14118 2802 14152
rect 2530 14074 2656 14118
rect 1242 13994 1248 13998
rect 1138 13950 1248 13994
rect 1138 13926 1182 13950
rect 1242 13946 1248 13950
rect 1300 13946 1306 13998
rect 1404 13981 1450 14014
rect 1404 13947 1410 13981
rect 1444 13947 1450 13981
rect 1404 13943 1450 13947
rect 378 13898 434 13904
rect 550 13898 622 13920
rect 434 13892 622 13898
rect 434 13852 565 13892
rect 606 13852 622 13892
rect 434 13842 622 13852
rect 378 13836 434 13842
rect 550 13822 622 13842
rect 696 13892 768 13920
rect 696 13852 712 13892
rect 753 13852 768 13892
rect 696 13822 768 13852
rect 840 13897 912 13926
rect 840 13857 856 13897
rect 897 13857 912 13897
rect 840 13828 912 13857
rect 994 13898 1182 13926
rect 994 13858 1010 13898
rect 1051 13882 1182 13898
rect 1399 13914 1450 13943
rect 1562 13981 1608 14014
rect 1562 13947 1568 13981
rect 1602 13947 1608 13981
rect 1692 13981 1738 14014
rect 1692 13952 1698 13981
rect 1562 13914 1608 13947
rect 1690 13947 1698 13952
rect 1732 13952 1738 13981
rect 1850 13981 1896 14014
rect 2024 13998 2070 14014
rect 1732 13947 1740 13952
rect 1051 13858 1066 13882
rect 1399 13868 1449 13914
rect 1690 13868 1740 13947
rect 1850 13947 1856 13981
rect 1890 13947 1896 13981
rect 1850 13914 1896 13947
rect 2014 13946 2020 13998
rect 2072 13946 2078 13998
rect 2182 13981 2228 14014
rect 2182 13947 2188 13981
rect 2222 13947 2228 13981
rect 2024 13914 2070 13946
rect 2182 13914 2228 13947
rect 2366 13981 2412 14014
rect 2524 13996 2570 14014
rect 2366 13947 2372 13981
rect 2406 13947 2412 13981
rect 2366 13914 2412 13947
rect 2516 13944 2522 13996
rect 2574 13944 2580 13996
rect 2524 13914 2570 13944
rect 2024 13882 2068 13914
rect 2612 13882 2656 14074
rect 994 13828 1066 13858
rect 1324 13813 1960 13868
rect 2024 13838 2656 13882
rect 2694 14074 2802 14118
rect 2832 14104 2904 14114
rect 2694 13876 2738 14074
rect 2832 14052 2842 14104
rect 2894 14052 2904 14104
rect 2832 14042 2904 14052
rect 2933 14014 2972 14152
rect 3118 14014 3157 14152
rect 3272 14108 3316 14152
rect 3268 14102 3320 14108
rect 3555 14077 3561 14129
rect 3613 14122 3619 14129
rect 3662 14122 3713 14134
rect 3613 14119 3713 14122
rect 3613 14085 3670 14119
rect 3704 14085 3713 14119
rect 3613 14083 3713 14085
rect 3613 14077 3619 14083
rect 3662 14071 3713 14083
rect 3897 14113 3936 14162
rect 3976 14120 4027 14125
rect 3970 14113 3976 14120
rect 3897 14074 3976 14113
rect 3268 14044 3320 14050
rect 3897 14024 3936 14074
rect 3970 14068 3976 14074
rect 4028 14068 4034 14120
rect 4206 14106 4245 14162
rect 4300 14106 4347 14117
rect 4206 14104 4347 14106
rect 4206 14071 4306 14104
rect 3976 14062 4027 14068
rect 4206 14024 4245 14071
rect 4300 14070 4306 14071
rect 4340 14070 4347 14104
rect 4300 14058 4347 14070
rect 2766 14008 2818 14014
rect 2766 13950 2776 13956
rect 2770 13947 2776 13950
rect 2810 13950 2818 13956
rect 2928 13981 2974 14014
rect 2810 13947 2816 13950
rect 2770 13914 2816 13947
rect 2928 13947 2934 13981
rect 2968 13947 2974 13981
rect 2928 13914 2974 13947
rect 3114 13981 3160 14014
rect 3114 13947 3120 13981
rect 3154 13947 3160 13981
rect 3114 13914 3160 13947
rect 3272 13981 3318 14014
rect 3272 13947 3278 13981
rect 3312 13947 3318 13981
rect 3272 13914 3318 13947
rect 3274 13876 3318 13914
rect 2694 13832 3318 13876
rect 3736 13991 3782 14024
rect 3736 13957 3742 13991
rect 3776 13957 3782 13991
rect 3736 13924 3782 13957
rect 3894 13991 3940 14024
rect 3894 13957 3900 13991
rect 3934 13957 3940 13991
rect 4044 13991 4090 14024
rect 4044 13962 4050 13991
rect 3894 13924 3940 13957
rect 4042 13957 4050 13962
rect 4084 13957 4090 13991
rect 4042 13924 4090 13957
rect 4202 13991 4248 14024
rect 4202 13957 4208 13991
rect 4242 13957 4248 13991
rect 4202 13924 4248 13957
rect 3736 13868 3780 13924
rect 4042 13868 4089 13924
rect 1324 13761 1360 13813
rect 1412 13761 1424 13813
rect 1476 13804 1488 13813
rect 1540 13804 1552 13813
rect 1604 13804 1616 13813
rect 1668 13804 1680 13813
rect 1732 13804 1744 13813
rect 1796 13804 1808 13813
rect 1479 13770 1488 13804
rect 1551 13770 1552 13804
rect 1732 13770 1733 13804
rect 1796 13770 1805 13804
rect 1476 13761 1488 13770
rect 1540 13761 1552 13770
rect 1604 13761 1616 13770
rect 1668 13761 1680 13770
rect 1732 13761 1744 13770
rect 1796 13761 1808 13770
rect 1860 13761 1872 13813
rect 1924 13761 1960 13813
rect 3704 13824 4244 13868
rect 3704 13815 3756 13824
rect 3808 13815 3820 13824
rect 1324 13728 1960 13761
rect 2346 13783 2426 13808
rect 2346 13779 3517 13783
rect 2346 13745 2369 13779
rect 2403 13745 3517 13779
rect 2346 13741 3517 13745
rect 2346 13716 2426 13741
rect 2636 13683 2702 13695
rect 272 13629 278 13683
rect 332 13629 2642 13683
rect 2696 13629 2702 13683
rect 2636 13617 2702 13629
rect 3475 13588 3517 13741
rect 3704 13781 3741 13815
rect 3808 13781 3813 13815
rect 3704 13772 3756 13781
rect 3808 13772 3820 13781
rect 3872 13772 3884 13824
rect 3936 13772 3948 13824
rect 4000 13772 4012 13824
rect 4064 13772 4076 13824
rect 4128 13815 4140 13824
rect 4192 13815 4244 13824
rect 4135 13781 4140 13815
rect 4207 13781 4244 13815
rect 4128 13772 4140 13781
rect 4192 13772 4244 13781
rect 3704 13728 4244 13772
rect 3559 13623 3565 13675
rect 3617 13668 3623 13675
rect 4306 13668 4345 14058
rect 4558 14026 4597 14162
rect 4628 14131 4680 14137
rect 4625 14082 4628 14128
rect 4680 14082 4683 14128
rect 4875 14086 4904 14162
rect 4628 14073 4680 14079
rect 4875 14058 4980 14086
rect 4396 13993 4442 14026
rect 4396 13959 4402 13993
rect 4436 13959 4442 13993
rect 4396 13926 4442 13959
rect 4554 14006 4600 14026
rect 4704 14006 4750 14026
rect 4862 14006 4908 14026
rect 4554 13993 4750 14006
rect 4554 13959 4560 13993
rect 4594 13959 4710 13993
rect 4744 13959 4750 13993
rect 4554 13940 4750 13959
rect 4856 13954 4862 14006
rect 4914 13954 4920 14006
rect 4554 13926 4600 13940
rect 4704 13926 4750 13940
rect 4862 13926 4908 13954
rect 4402 13776 4430 13926
rect 4558 13881 4597 13926
rect 4552 13875 4604 13881
rect 4552 13817 4604 13823
rect 4952 13776 4980 14058
rect 5026 14008 5056 14193
rect 5694 14162 5740 14210
rect 5852 14316 5898 14362
rect 5852 14282 5858 14316
rect 5892 14282 5898 14316
rect 5852 14244 5898 14282
rect 5852 14210 5858 14244
rect 5892 14210 5898 14244
rect 5852 14162 5898 14210
rect 6002 14316 6048 14418
rect 6516 14362 6556 14568
rect 6862 14562 6868 14568
rect 6920 14562 6926 14614
rect 6985 14602 7015 14655
rect 6985 14573 7016 14602
rect 6002 14282 6008 14316
rect 6042 14282 6048 14316
rect 6002 14244 6048 14282
rect 6002 14210 6008 14244
rect 6042 14210 6048 14244
rect 6002 14162 6048 14210
rect 6160 14316 6206 14362
rect 6160 14282 6166 14316
rect 6200 14282 6206 14316
rect 6354 14316 6400 14362
rect 6354 14290 6360 14316
rect 6160 14244 6206 14282
rect 6160 14210 6166 14244
rect 6200 14210 6206 14244
rect 6244 14288 6360 14290
rect 6244 14236 6250 14288
rect 6302 14282 6360 14288
rect 6394 14282 6400 14316
rect 6302 14244 6400 14282
rect 6302 14236 6360 14244
rect 6244 14234 6360 14236
rect 6160 14162 6206 14210
rect 6354 14210 6360 14234
rect 6394 14210 6400 14244
rect 6354 14162 6400 14210
rect 6512 14316 6558 14362
rect 6512 14282 6518 14316
rect 6552 14282 6558 14316
rect 6662 14316 6708 14362
rect 6662 14282 6668 14316
rect 6702 14282 6708 14316
rect 6512 14244 6708 14282
rect 6512 14210 6518 14244
rect 6552 14216 6668 14244
rect 6552 14210 6558 14216
rect 6512 14162 6558 14210
rect 6662 14210 6668 14216
rect 6702 14210 6708 14244
rect 6662 14162 6708 14210
rect 6820 14316 6866 14362
rect 6820 14282 6826 14316
rect 6860 14282 6866 14316
rect 6986 14286 7016 14573
rect 7206 14502 7234 14760
rect 7194 14496 7246 14502
rect 7194 14438 7246 14444
rect 6820 14244 6866 14282
rect 6820 14210 6826 14244
rect 6860 14210 6866 14244
rect 6968 14234 6974 14286
rect 7026 14234 7032 14286
rect 6820 14162 6866 14210
rect 6984 14194 7016 14234
rect 5111 14077 5117 14129
rect 5169 14122 5175 14129
rect 5620 14122 5672 14134
rect 5169 14120 5672 14122
rect 5169 14086 5628 14120
rect 5662 14086 5672 14120
rect 5169 14083 5672 14086
rect 5169 14077 5175 14083
rect 5620 14072 5672 14083
rect 5856 14114 5894 14162
rect 5934 14120 5986 14126
rect 5928 14114 5934 14120
rect 5856 14074 5934 14114
rect 5856 14024 5894 14074
rect 5928 14068 5934 14074
rect 5986 14068 5992 14120
rect 6164 14106 6204 14162
rect 6258 14106 6306 14118
rect 6164 14104 6306 14106
rect 6164 14072 6264 14104
rect 5934 14062 5986 14068
rect 6164 14024 6204 14072
rect 6258 14070 6264 14072
rect 6298 14070 6306 14104
rect 6258 14058 6306 14070
rect 5009 13956 5015 14008
rect 5067 13956 5073 14008
rect 5694 13992 5740 14024
rect 5694 13958 5700 13992
rect 5734 13958 5740 13992
rect 4402 13748 4980 13776
rect 3617 13629 4345 13668
rect 3617 13623 3623 13629
rect 5021 13588 5063 13956
rect 5694 13924 5740 13958
rect 5852 13992 5898 14024
rect 5852 13958 5858 13992
rect 5892 13958 5898 13992
rect 6002 13992 6048 14024
rect 6002 13962 6008 13992
rect 5852 13924 5898 13958
rect 6000 13958 6008 13962
rect 6042 13958 6048 13992
rect 5694 13868 5738 13924
rect 6000 13868 6048 13958
rect 6160 13992 6206 14024
rect 6160 13958 6166 13992
rect 6200 13958 6206 13992
rect 6160 13924 6206 13958
rect 5662 13824 6202 13868
rect 5662 13816 5714 13824
rect 5766 13816 5778 13824
rect 5662 13782 5700 13816
rect 5766 13782 5772 13816
rect 5662 13772 5714 13782
rect 5766 13772 5778 13782
rect 5830 13772 5842 13824
rect 5894 13772 5906 13824
rect 5958 13772 5970 13824
rect 6022 13772 6034 13824
rect 6086 13816 6098 13824
rect 6150 13816 6202 13824
rect 6094 13782 6098 13816
rect 6166 13782 6202 13816
rect 6086 13772 6098 13782
rect 6150 13772 6202 13782
rect 5662 13728 6202 13772
rect 5111 13623 5117 13675
rect 5169 13668 5175 13675
rect 6264 13668 6304 14058
rect 6516 14026 6556 14162
rect 6586 14132 6638 14138
rect 6584 14082 6586 14128
rect 6638 14082 6642 14128
rect 6834 14086 6862 14162
rect 6586 14074 6638 14080
rect 6834 14058 6936 14086
rect 6354 13994 6400 14026
rect 6354 13960 6360 13994
rect 6394 13960 6400 13994
rect 6354 13926 6400 13960
rect 6512 14006 6558 14026
rect 6662 14006 6708 14026
rect 6820 14006 6866 14026
rect 6512 13994 6708 14006
rect 6512 13960 6518 13994
rect 6552 13960 6668 13994
rect 6702 13960 6708 13994
rect 6512 13940 6708 13960
rect 6814 13954 6820 14006
rect 6872 13954 6878 14006
rect 6512 13926 6558 13940
rect 6662 13926 6708 13940
rect 6820 13926 6866 13954
rect 6360 13776 6388 13926
rect 6516 13882 6556 13926
rect 6510 13876 6562 13882
rect 6510 13818 6562 13824
rect 6908 13776 6936 14058
rect 6984 14008 7014 14194
rect 6968 13956 6974 14008
rect 7026 13956 7032 14008
rect 6360 13748 6936 13776
rect 6908 13684 6936 13748
rect 5169 13630 6304 13668
rect 6346 13656 6936 13684
rect 5169 13629 5572 13630
rect 5169 13623 5175 13629
rect 3475 13546 5063 13588
rect 5035 13505 5087 13511
rect 3472 13421 4907 13460
rect 6346 13493 6374 13656
rect 6908 13654 6936 13656
rect 6512 13590 6564 13596
rect 6512 13532 6564 13538
rect 5087 13465 6374 13493
rect 6523 13475 6553 13532
rect 5035 13447 5087 13453
rect 6523 13445 7015 13475
rect 1348 13287 1880 13330
rect 1348 13278 1398 13287
rect 1450 13278 1462 13287
rect 1348 13244 1383 13278
rect 1450 13244 1455 13278
rect 1348 13235 1398 13244
rect 1450 13235 1462 13244
rect 1514 13235 1526 13287
rect 1578 13235 1590 13287
rect 1642 13235 1654 13287
rect 1706 13235 1718 13287
rect 1770 13278 1782 13287
rect 1834 13278 1880 13287
rect 1777 13244 1782 13278
rect 1849 13244 1880 13278
rect 3472 13263 3511 13421
rect 4738 13379 4744 13386
rect 4558 13340 4744 13379
rect 1770 13235 1782 13244
rect 1834 13235 1880 13244
rect 550 13216 622 13220
rect 550 13164 560 13216
rect 612 13164 622 13216
rect 696 13214 768 13220
rect 550 13152 566 13164
rect 607 13152 622 13164
rect 682 13212 768 13214
rect 682 13160 702 13212
rect 754 13160 768 13212
rect 682 13158 710 13160
rect 550 13122 622 13152
rect 696 13152 710 13158
rect 751 13152 768 13160
rect 696 13122 768 13152
rect 840 13197 912 13226
rect 840 13157 856 13197
rect 897 13157 912 13197
rect 840 13128 912 13157
rect 994 13197 1066 13226
rect 994 13157 1009 13197
rect 1050 13157 1066 13197
rect 1348 13190 1880 13235
rect 994 13128 1066 13157
rect 564 13082 608 13122
rect 856 13062 900 13128
rect 378 13054 433 13060
rect 846 13010 852 13062
rect 904 13010 910 13062
rect 378 12769 433 12999
rect 856 12970 900 13010
rect 1008 12970 1052 13128
rect 1407 13124 1448 13190
rect 1693 13124 1735 13190
rect 1941 13187 2687 13232
rect 1404 13077 1450 13124
rect 1404 13043 1410 13077
rect 1444 13043 1450 13077
rect 1404 13005 1450 13043
rect 1404 12971 1410 13005
rect 1444 12971 1450 13005
rect 708 12926 900 12970
rect 372 12714 378 12769
rect 433 12714 439 12769
rect 708 12692 752 12926
rect 998 12918 1004 12970
rect 1056 12918 1062 12970
rect 1404 12924 1450 12971
rect 1562 13077 1608 13124
rect 1562 13043 1568 13077
rect 1602 13043 1608 13077
rect 1562 13005 1608 13043
rect 1562 12971 1568 13005
rect 1602 12971 1608 13005
rect 1562 12924 1608 12971
rect 1692 13077 1738 13124
rect 1692 13043 1698 13077
rect 1732 13043 1738 13077
rect 1692 13005 1738 13043
rect 1692 12971 1698 13005
rect 1732 12971 1738 13005
rect 1692 12924 1738 12971
rect 1850 13121 1896 13124
rect 1941 13121 1986 13187
rect 1850 13077 1986 13121
rect 1850 13043 1856 13077
rect 1890 13076 1986 13077
rect 2024 13077 2070 13124
rect 1890 13043 1896 13076
rect 1850 13005 1896 13043
rect 2024 13043 2030 13077
rect 2064 13043 2070 13077
rect 2024 13008 2070 13043
rect 1998 13006 2070 13008
rect 1850 12971 1856 13005
rect 1890 12971 1896 13005
rect 1850 12924 1896 12971
rect 1928 13005 2070 13006
rect 1928 12981 2030 13005
rect 1928 12964 1935 12981
rect 1929 12929 1935 12964
rect 1987 12971 2030 12981
rect 2064 12971 2070 13005
rect 1987 12964 2070 12971
rect 1987 12929 1993 12964
rect 2024 12924 2070 12964
rect 2182 13080 2228 13124
rect 2366 13080 2412 13124
rect 2182 13077 2412 13080
rect 2182 13043 2188 13077
rect 2222 13043 2372 13077
rect 2406 13043 2412 13077
rect 2182 13005 2412 13043
rect 2182 12971 2188 13005
rect 2222 12971 2372 13005
rect 2406 12971 2412 13005
rect 2182 12954 2412 12971
rect 2182 12924 2228 12954
rect 2366 12924 2412 12954
rect 2524 13077 2570 13124
rect 2524 13043 2530 13077
rect 2564 13043 2570 13077
rect 2642 13053 2687 13187
rect 3118 13224 3511 13263
rect 3724 13286 4264 13330
rect 3724 13234 3776 13286
rect 3828 13277 3840 13286
rect 3892 13277 3904 13286
rect 3956 13277 3968 13286
rect 4020 13277 4032 13286
rect 4084 13277 4096 13286
rect 4148 13277 4160 13286
rect 3831 13243 3840 13277
rect 3903 13243 3904 13277
rect 4084 13243 4085 13277
rect 4148 13243 4157 13277
rect 3828 13234 3840 13243
rect 3892 13234 3904 13243
rect 3956 13234 3968 13243
rect 4020 13234 4032 13243
rect 4084 13234 4096 13243
rect 4148 13234 4160 13243
rect 4212 13234 4264 13286
rect 2774 13180 2816 13181
rect 2758 13172 2816 13180
rect 2758 13120 2769 13172
rect 2821 13120 2827 13172
rect 3118 13124 3157 13224
rect 3724 13190 4264 13234
rect 3741 13134 3787 13190
rect 3736 13133 3787 13134
rect 2758 13077 2816 13120
rect 2524 13005 2570 13043
rect 2524 12971 2530 13005
rect 2564 12971 2570 13005
rect 2524 12964 2570 12971
rect 2613 13025 2715 13053
rect 2613 12991 2647 13025
rect 2681 12991 2715 13025
rect 2524 12924 2574 12964
rect 2613 12963 2715 12991
rect 2758 13043 2776 13077
rect 2810 13043 2816 13077
rect 2758 13005 2816 13043
rect 2758 12971 2776 13005
rect 2810 12971 2816 13005
rect 1008 12864 1052 12918
rect 1245 12883 1328 12902
rect 852 12820 1052 12864
rect 1148 12881 1328 12883
rect 1148 12829 1155 12881
rect 1207 12871 1328 12881
rect 1207 12837 1269 12871
rect 1303 12837 1328 12871
rect 1207 12829 1328 12837
rect 1148 12828 1328 12829
rect 852 12698 896 12820
rect 1245 12807 1328 12828
rect 1568 12890 1602 12924
rect 1568 12880 1820 12890
rect 1568 12828 1758 12880
rect 1810 12828 1820 12880
rect 1568 12818 1820 12828
rect 1568 12786 1608 12818
rect 1853 12786 1892 12924
rect 2185 12786 2224 12924
rect 2255 12887 2325 12893
rect 2255 12878 2331 12887
rect 2255 12826 2270 12878
rect 2322 12826 2331 12878
rect 2255 12817 2331 12826
rect 2255 12811 2325 12817
rect 2368 12786 2407 12924
rect 2530 12890 2574 12924
rect 2758 12924 2816 12971
rect 2928 13077 2974 13124
rect 2928 13043 2934 13077
rect 2968 13064 2974 13077
rect 3114 13077 3160 13124
rect 3114 13064 3120 13077
rect 2968 13043 3120 13064
rect 3154 13043 3160 13077
rect 3272 13077 3318 13124
rect 3272 13067 3278 13077
rect 3312 13067 3318 13077
rect 3736 13087 3782 13133
rect 2928 13005 3160 13043
rect 3262 13015 3268 13067
rect 3320 13015 3326 13067
rect 3736 13053 3742 13087
rect 3776 13053 3782 13087
rect 3736 13015 3782 13053
rect 2928 12971 2934 13005
rect 2968 12971 3120 13005
rect 3154 12971 3160 13005
rect 2928 12954 3160 12971
rect 2928 12924 2974 12954
rect 3114 12924 3160 12954
rect 3272 13005 3318 13015
rect 3272 12971 3278 13005
rect 3312 12971 3318 13005
rect 3272 12924 3318 12971
rect 3736 12981 3742 13015
rect 3776 12981 3782 13015
rect 3736 12934 3782 12981
rect 3894 13087 3940 13134
rect 3894 13053 3900 13087
rect 3934 13053 3940 13087
rect 3894 13015 3940 13053
rect 3894 12981 3900 13015
rect 3934 12981 3940 13015
rect 3894 12934 3940 12981
rect 4044 13087 4090 13190
rect 4558 13134 4597 13340
rect 4738 13334 4744 13340
rect 4796 13334 4802 13386
rect 4868 13134 4907 13421
rect 6837 13379 6843 13386
rect 6516 13340 6843 13379
rect 5682 13286 6222 13330
rect 5682 13234 5734 13286
rect 5786 13276 5798 13286
rect 5850 13276 5862 13286
rect 5914 13276 5926 13286
rect 5978 13276 5990 13286
rect 6042 13276 6054 13286
rect 6106 13276 6118 13286
rect 5790 13242 5798 13276
rect 6042 13242 6044 13276
rect 6106 13242 6116 13276
rect 5786 13234 5798 13242
rect 5850 13234 5862 13242
rect 5914 13234 5926 13242
rect 5978 13234 5990 13242
rect 6042 13234 6054 13242
rect 6106 13234 6118 13242
rect 6170 13234 6222 13286
rect 5682 13190 6222 13234
rect 5700 13134 5746 13190
rect 4044 13053 4050 13087
rect 4084 13053 4090 13087
rect 4044 13015 4090 13053
rect 4044 12981 4050 13015
rect 4084 12981 4090 13015
rect 4044 12934 4090 12981
rect 4202 13087 4248 13134
rect 4202 13053 4208 13087
rect 4242 13053 4248 13087
rect 4396 13087 4442 13134
rect 4396 13061 4402 13087
rect 4202 13015 4248 13053
rect 4202 12981 4208 13015
rect 4242 12981 4248 13015
rect 4285 13059 4402 13061
rect 4285 13007 4292 13059
rect 4344 13053 4402 13059
rect 4436 13053 4442 13087
rect 4344 13015 4442 13053
rect 4344 13007 4402 13015
rect 4285 13006 4402 13007
rect 4202 12934 4248 12981
rect 4396 12981 4402 13006
rect 4436 12981 4442 13015
rect 4396 12934 4442 12981
rect 4554 13087 4600 13134
rect 4554 13053 4560 13087
rect 4594 13054 4600 13087
rect 4704 13087 4750 13134
rect 4704 13054 4710 13087
rect 4594 13053 4710 13054
rect 4744 13053 4750 13087
rect 4554 13015 4750 13053
rect 4554 12981 4560 13015
rect 4594 12988 4710 13015
rect 4594 12981 4600 12988
rect 4554 12934 4600 12981
rect 4704 12981 4710 12988
rect 4744 12981 4750 13015
rect 4704 12934 4750 12981
rect 4862 13087 4908 13134
rect 4862 13053 4868 13087
rect 4902 13053 4908 13087
rect 5694 13088 5740 13134
rect 5027 13058 5057 13067
rect 4862 13015 4908 13053
rect 4862 12981 4868 13015
rect 4902 12981 4908 13015
rect 5010 13006 5016 13058
rect 5068 13006 5074 13058
rect 5694 13054 5700 13088
rect 5734 13054 5740 13088
rect 5694 13016 5740 13054
rect 4862 12934 4908 12981
rect 5026 12965 5057 13006
rect 5694 12982 5700 13016
rect 5734 12982 5740 13016
rect 2758 12890 2802 12924
rect 2530 12846 2656 12890
rect 1242 12766 1248 12770
rect 1138 12722 1248 12766
rect 1138 12698 1182 12722
rect 1242 12718 1248 12722
rect 1300 12718 1306 12770
rect 1404 12753 1450 12786
rect 1404 12719 1410 12753
rect 1444 12719 1450 12753
rect 1404 12715 1450 12719
rect 378 12670 434 12676
rect 550 12670 622 12692
rect 434 12664 622 12670
rect 434 12624 565 12664
rect 606 12624 622 12664
rect 434 12614 622 12624
rect 378 12608 434 12614
rect 550 12594 622 12614
rect 696 12664 768 12692
rect 696 12624 712 12664
rect 753 12624 768 12664
rect 696 12594 768 12624
rect 840 12669 912 12698
rect 840 12629 856 12669
rect 897 12629 912 12669
rect 840 12600 912 12629
rect 994 12670 1182 12698
rect 994 12630 1010 12670
rect 1051 12654 1182 12670
rect 1399 12686 1450 12715
rect 1562 12753 1608 12786
rect 1562 12719 1568 12753
rect 1602 12719 1608 12753
rect 1692 12753 1738 12786
rect 1692 12724 1698 12753
rect 1562 12686 1608 12719
rect 1690 12719 1698 12724
rect 1732 12724 1738 12753
rect 1850 12753 1896 12786
rect 2024 12770 2070 12786
rect 1732 12719 1740 12724
rect 1051 12630 1066 12654
rect 1399 12640 1449 12686
rect 1690 12640 1740 12719
rect 1850 12719 1856 12753
rect 1890 12719 1896 12753
rect 1850 12686 1896 12719
rect 2014 12718 2020 12770
rect 2072 12718 2078 12770
rect 2182 12753 2228 12786
rect 2182 12719 2188 12753
rect 2222 12719 2228 12753
rect 2024 12686 2070 12718
rect 2182 12686 2228 12719
rect 2366 12753 2412 12786
rect 2524 12768 2570 12786
rect 2366 12719 2372 12753
rect 2406 12719 2412 12753
rect 2366 12686 2412 12719
rect 2516 12716 2522 12768
rect 2574 12716 2580 12768
rect 2524 12686 2570 12716
rect 2024 12654 2068 12686
rect 2612 12654 2656 12846
rect 994 12600 1066 12630
rect 1324 12585 1960 12640
rect 2024 12610 2656 12654
rect 2694 12846 2802 12890
rect 2832 12876 2904 12886
rect 2694 12648 2738 12846
rect 2832 12824 2842 12876
rect 2894 12824 2904 12876
rect 2832 12814 2904 12824
rect 2933 12786 2972 12924
rect 3118 12786 3157 12924
rect 3272 12880 3316 12924
rect 3268 12874 3320 12880
rect 3555 12849 3561 12901
rect 3613 12894 3619 12901
rect 3662 12894 3713 12906
rect 3613 12891 3713 12894
rect 3613 12857 3670 12891
rect 3704 12857 3713 12891
rect 3613 12855 3713 12857
rect 3613 12849 3619 12855
rect 3662 12843 3713 12855
rect 3897 12885 3936 12934
rect 3976 12892 4027 12897
rect 3970 12885 3976 12892
rect 3897 12846 3976 12885
rect 3268 12816 3320 12822
rect 3897 12796 3936 12846
rect 3970 12840 3976 12846
rect 4028 12840 4034 12892
rect 4206 12878 4245 12934
rect 4300 12878 4347 12889
rect 4206 12876 4347 12878
rect 4206 12843 4306 12876
rect 3976 12834 4027 12840
rect 4206 12796 4245 12843
rect 4300 12842 4306 12843
rect 4340 12842 4347 12876
rect 4300 12830 4347 12842
rect 2766 12780 2818 12786
rect 2766 12722 2776 12728
rect 2770 12719 2776 12722
rect 2810 12722 2818 12728
rect 2928 12753 2974 12786
rect 2810 12719 2816 12722
rect 2770 12686 2816 12719
rect 2928 12719 2934 12753
rect 2968 12719 2974 12753
rect 2928 12686 2974 12719
rect 3114 12753 3160 12786
rect 3114 12719 3120 12753
rect 3154 12719 3160 12753
rect 3114 12686 3160 12719
rect 3272 12753 3318 12786
rect 3272 12719 3278 12753
rect 3312 12719 3318 12753
rect 3272 12686 3318 12719
rect 3274 12648 3318 12686
rect 2694 12604 3318 12648
rect 3736 12763 3782 12796
rect 3736 12729 3742 12763
rect 3776 12729 3782 12763
rect 3736 12696 3782 12729
rect 3894 12763 3940 12796
rect 3894 12729 3900 12763
rect 3934 12729 3940 12763
rect 4044 12763 4090 12796
rect 4044 12734 4050 12763
rect 3894 12696 3940 12729
rect 4042 12729 4050 12734
rect 4084 12729 4090 12763
rect 4042 12696 4090 12729
rect 4202 12763 4248 12796
rect 4202 12729 4208 12763
rect 4242 12729 4248 12763
rect 4202 12696 4248 12729
rect 3736 12640 3780 12696
rect 4042 12640 4089 12696
rect 1324 12533 1360 12585
rect 1412 12533 1424 12585
rect 1476 12576 1488 12585
rect 1540 12576 1552 12585
rect 1604 12576 1616 12585
rect 1668 12576 1680 12585
rect 1732 12576 1744 12585
rect 1796 12576 1808 12585
rect 1479 12542 1488 12576
rect 1551 12542 1552 12576
rect 1732 12542 1733 12576
rect 1796 12542 1805 12576
rect 1476 12533 1488 12542
rect 1540 12533 1552 12542
rect 1604 12533 1616 12542
rect 1668 12533 1680 12542
rect 1732 12533 1744 12542
rect 1796 12533 1808 12542
rect 1860 12533 1872 12585
rect 1924 12533 1960 12585
rect 3704 12596 4244 12640
rect 3704 12587 3756 12596
rect 3808 12587 3820 12596
rect 1324 12500 1960 12533
rect 2346 12555 2426 12580
rect 2346 12551 3517 12555
rect 2346 12517 2369 12551
rect 2403 12517 3517 12551
rect 2346 12513 3517 12517
rect 2346 12488 2426 12513
rect 2636 12455 2702 12467
rect 272 12401 278 12455
rect 332 12401 2642 12455
rect 2696 12401 2702 12455
rect 2636 12389 2702 12401
rect 3475 12360 3517 12513
rect 3704 12553 3741 12587
rect 3808 12553 3813 12587
rect 3704 12544 3756 12553
rect 3808 12544 3820 12553
rect 3872 12544 3884 12596
rect 3936 12544 3948 12596
rect 4000 12544 4012 12596
rect 4064 12544 4076 12596
rect 4128 12587 4140 12596
rect 4192 12587 4244 12596
rect 4135 12553 4140 12587
rect 4207 12553 4244 12587
rect 4128 12544 4140 12553
rect 4192 12544 4244 12553
rect 3704 12500 4244 12544
rect 3559 12395 3565 12447
rect 3617 12440 3623 12447
rect 4306 12440 4345 12830
rect 4558 12798 4597 12934
rect 4628 12903 4680 12909
rect 4625 12854 4628 12900
rect 4680 12854 4683 12900
rect 4875 12858 4904 12934
rect 4628 12845 4680 12851
rect 4875 12830 4980 12858
rect 4396 12765 4442 12798
rect 4396 12731 4402 12765
rect 4436 12731 4442 12765
rect 4396 12698 4442 12731
rect 4554 12778 4600 12798
rect 4704 12778 4750 12798
rect 4862 12778 4908 12798
rect 4554 12765 4750 12778
rect 4554 12731 4560 12765
rect 4594 12731 4710 12765
rect 4744 12731 4750 12765
rect 4554 12712 4750 12731
rect 4856 12726 4862 12778
rect 4914 12726 4920 12778
rect 4554 12698 4600 12712
rect 4704 12698 4750 12712
rect 4862 12698 4908 12726
rect 4402 12548 4430 12698
rect 4558 12653 4597 12698
rect 4552 12647 4604 12653
rect 4552 12589 4604 12595
rect 4952 12548 4980 12830
rect 5026 12780 5056 12965
rect 5694 12934 5740 12982
rect 5852 13088 5898 13134
rect 5852 13054 5858 13088
rect 5892 13054 5898 13088
rect 5852 13016 5898 13054
rect 5852 12982 5858 13016
rect 5892 12982 5898 13016
rect 5852 12934 5898 12982
rect 6002 13088 6048 13190
rect 6516 13134 6556 13340
rect 6837 13334 6843 13340
rect 6895 13334 6901 13386
rect 6985 13374 7015 13445
rect 6985 13345 7016 13374
rect 6002 13054 6008 13088
rect 6042 13054 6048 13088
rect 6002 13016 6048 13054
rect 6002 12982 6008 13016
rect 6042 12982 6048 13016
rect 6002 12934 6048 12982
rect 6160 13088 6206 13134
rect 6160 13054 6166 13088
rect 6200 13054 6206 13088
rect 6354 13088 6400 13134
rect 6354 13062 6360 13088
rect 6160 13016 6206 13054
rect 6160 12982 6166 13016
rect 6200 12982 6206 13016
rect 6244 13060 6360 13062
rect 6244 13008 6250 13060
rect 6302 13054 6360 13060
rect 6394 13054 6400 13088
rect 6302 13016 6400 13054
rect 6302 13008 6360 13016
rect 6244 13006 6360 13008
rect 6160 12934 6206 12982
rect 6354 12982 6360 13006
rect 6394 12982 6400 13016
rect 6354 12934 6400 12982
rect 6512 13088 6558 13134
rect 6512 13054 6518 13088
rect 6552 13054 6558 13088
rect 6662 13088 6708 13134
rect 6662 13054 6668 13088
rect 6702 13054 6708 13088
rect 6512 13016 6708 13054
rect 6512 12982 6518 13016
rect 6552 12988 6668 13016
rect 6552 12982 6558 12988
rect 6512 12934 6558 12982
rect 6662 12982 6668 12988
rect 6702 12982 6708 13016
rect 6662 12934 6708 12982
rect 6820 13088 6866 13134
rect 6820 13054 6826 13088
rect 6860 13054 6866 13088
rect 6986 13058 7016 13345
rect 6820 13016 6866 13054
rect 6820 12982 6826 13016
rect 6860 12982 6866 13016
rect 6968 13006 6974 13058
rect 7026 13006 7032 13058
rect 6820 12934 6866 12982
rect 6984 12966 7016 13006
rect 5191 12849 5197 12901
rect 5249 12894 5255 12901
rect 5620 12894 5672 12906
rect 5249 12892 5672 12894
rect 5249 12858 5628 12892
rect 5662 12858 5672 12892
rect 5249 12855 5672 12858
rect 5249 12849 5255 12855
rect 5620 12844 5672 12855
rect 5856 12886 5894 12934
rect 5934 12892 5986 12898
rect 5928 12886 5934 12892
rect 5856 12846 5934 12886
rect 5856 12796 5894 12846
rect 5928 12840 5934 12846
rect 5986 12840 5992 12892
rect 6164 12878 6204 12934
rect 6258 12878 6306 12890
rect 6164 12876 6306 12878
rect 6164 12844 6264 12876
rect 5934 12834 5986 12840
rect 6164 12796 6204 12844
rect 6258 12842 6264 12844
rect 6298 12842 6306 12876
rect 6258 12830 6306 12842
rect 5009 12728 5015 12780
rect 5067 12728 5073 12780
rect 5694 12764 5740 12796
rect 5694 12730 5700 12764
rect 5734 12730 5740 12764
rect 4402 12520 4980 12548
rect 3617 12401 4345 12440
rect 3617 12395 3623 12401
rect 5021 12360 5063 12728
rect 5694 12696 5740 12730
rect 5852 12764 5898 12796
rect 5852 12730 5858 12764
rect 5892 12730 5898 12764
rect 6002 12764 6048 12796
rect 6002 12734 6008 12764
rect 5852 12696 5898 12730
rect 6000 12730 6008 12734
rect 6042 12730 6048 12764
rect 5694 12640 5738 12696
rect 6000 12640 6048 12730
rect 6160 12764 6206 12796
rect 6160 12730 6166 12764
rect 6200 12730 6206 12764
rect 6160 12696 6206 12730
rect 5662 12596 6202 12640
rect 5662 12588 5714 12596
rect 5766 12588 5778 12596
rect 5662 12554 5700 12588
rect 5766 12554 5772 12588
rect 5662 12544 5714 12554
rect 5766 12544 5778 12554
rect 5830 12544 5842 12596
rect 5894 12544 5906 12596
rect 5958 12544 5970 12596
rect 6022 12544 6034 12596
rect 6086 12588 6098 12596
rect 6150 12588 6202 12596
rect 6094 12554 6098 12588
rect 6166 12554 6202 12588
rect 6086 12544 6098 12554
rect 6150 12544 6202 12554
rect 5662 12500 6202 12544
rect 5191 12395 5197 12447
rect 5249 12440 5255 12447
rect 6264 12440 6304 12830
rect 6516 12798 6556 12934
rect 6586 12904 6638 12910
rect 6584 12854 6586 12900
rect 6638 12854 6642 12900
rect 6834 12858 6862 12934
rect 6586 12846 6638 12852
rect 6834 12830 6936 12858
rect 6354 12766 6400 12798
rect 6354 12732 6360 12766
rect 6394 12732 6400 12766
rect 6354 12698 6400 12732
rect 6512 12778 6558 12798
rect 6662 12778 6708 12798
rect 6820 12778 6866 12798
rect 6512 12766 6708 12778
rect 6512 12732 6518 12766
rect 6552 12732 6668 12766
rect 6702 12732 6708 12766
rect 6512 12712 6708 12732
rect 6814 12726 6820 12778
rect 6872 12726 6878 12778
rect 6512 12698 6558 12712
rect 6662 12698 6708 12712
rect 6820 12698 6866 12726
rect 6360 12548 6388 12698
rect 6516 12654 6556 12698
rect 6510 12648 6562 12654
rect 6510 12590 6562 12596
rect 6908 12548 6936 12830
rect 6984 12780 7014 12966
rect 6968 12728 6974 12780
rect 7026 12728 7032 12780
rect 6360 12520 6936 12548
rect 5249 12402 6304 12440
rect 5249 12401 5587 12402
rect 5249 12395 5255 12401
rect 3475 12318 5063 12360
rect 6908 12348 6936 12520
rect 7107 12360 7159 12366
rect 6908 12320 7107 12348
rect 7107 12302 7159 12308
rect 5029 12240 5081 12246
rect 3472 12193 4907 12232
rect 1348 12059 1880 12102
rect 1348 12050 1398 12059
rect 1450 12050 1462 12059
rect 1348 12016 1383 12050
rect 1450 12016 1455 12050
rect 1348 12007 1398 12016
rect 1450 12007 1462 12016
rect 1514 12007 1526 12059
rect 1578 12007 1590 12059
rect 1642 12007 1654 12059
rect 1706 12007 1718 12059
rect 1770 12050 1782 12059
rect 1834 12050 1880 12059
rect 1777 12016 1782 12050
rect 1849 12016 1880 12050
rect 3472 12035 3511 12193
rect 4738 12151 4744 12158
rect 4558 12112 4744 12151
rect 1770 12007 1782 12016
rect 1834 12007 1880 12016
rect 550 11988 622 11992
rect 550 11936 560 11988
rect 612 11936 622 11988
rect 696 11986 768 11992
rect 550 11924 566 11936
rect 607 11924 622 11936
rect 682 11984 768 11986
rect 682 11932 702 11984
rect 754 11932 768 11984
rect 682 11930 710 11932
rect 550 11894 622 11924
rect 696 11924 710 11930
rect 751 11924 768 11932
rect 696 11894 768 11924
rect 840 11969 912 11998
rect 840 11929 856 11969
rect 897 11929 912 11969
rect 840 11900 912 11929
rect 994 11969 1066 11998
rect 994 11929 1009 11969
rect 1050 11929 1066 11969
rect 1348 11962 1880 12007
rect 994 11900 1066 11929
rect 564 11854 608 11894
rect 856 11834 900 11900
rect 378 11826 433 11832
rect 846 11782 852 11834
rect 904 11782 910 11834
rect 378 11541 433 11771
rect 856 11742 900 11782
rect 1008 11742 1052 11900
rect 1407 11896 1448 11962
rect 1693 11896 1735 11962
rect 1941 11959 2687 12004
rect 1404 11849 1450 11896
rect 1404 11815 1410 11849
rect 1444 11815 1450 11849
rect 1404 11777 1450 11815
rect 1404 11743 1410 11777
rect 1444 11743 1450 11777
rect 708 11698 900 11742
rect 372 11486 378 11541
rect 433 11486 439 11541
rect 708 11464 752 11698
rect 998 11690 1004 11742
rect 1056 11690 1062 11742
rect 1404 11696 1450 11743
rect 1562 11849 1608 11896
rect 1562 11815 1568 11849
rect 1602 11815 1608 11849
rect 1562 11777 1608 11815
rect 1562 11743 1568 11777
rect 1602 11743 1608 11777
rect 1562 11696 1608 11743
rect 1692 11849 1738 11896
rect 1692 11815 1698 11849
rect 1732 11815 1738 11849
rect 1692 11777 1738 11815
rect 1692 11743 1698 11777
rect 1732 11743 1738 11777
rect 1692 11696 1738 11743
rect 1850 11893 1896 11896
rect 1941 11893 1986 11959
rect 1850 11849 1986 11893
rect 1850 11815 1856 11849
rect 1890 11848 1986 11849
rect 2024 11849 2070 11896
rect 1890 11815 1896 11848
rect 1850 11777 1896 11815
rect 2024 11815 2030 11849
rect 2064 11815 2070 11849
rect 2024 11780 2070 11815
rect 1998 11778 2070 11780
rect 1850 11743 1856 11777
rect 1890 11743 1896 11777
rect 1850 11696 1896 11743
rect 1928 11777 2070 11778
rect 1928 11753 2030 11777
rect 1928 11736 1935 11753
rect 1929 11701 1935 11736
rect 1987 11743 2030 11753
rect 2064 11743 2070 11777
rect 1987 11736 2070 11743
rect 1987 11701 1993 11736
rect 2024 11696 2070 11736
rect 2182 11852 2228 11896
rect 2366 11852 2412 11896
rect 2182 11849 2412 11852
rect 2182 11815 2188 11849
rect 2222 11815 2372 11849
rect 2406 11815 2412 11849
rect 2182 11777 2412 11815
rect 2182 11743 2188 11777
rect 2222 11743 2372 11777
rect 2406 11743 2412 11777
rect 2182 11726 2412 11743
rect 2182 11696 2228 11726
rect 2366 11696 2412 11726
rect 2524 11849 2570 11896
rect 2524 11815 2530 11849
rect 2564 11815 2570 11849
rect 2642 11825 2687 11959
rect 3118 11996 3511 12035
rect 3724 12058 4264 12102
rect 3724 12006 3776 12058
rect 3828 12049 3840 12058
rect 3892 12049 3904 12058
rect 3956 12049 3968 12058
rect 4020 12049 4032 12058
rect 4084 12049 4096 12058
rect 4148 12049 4160 12058
rect 3831 12015 3840 12049
rect 3903 12015 3904 12049
rect 4084 12015 4085 12049
rect 4148 12015 4157 12049
rect 3828 12006 3840 12015
rect 3892 12006 3904 12015
rect 3956 12006 3968 12015
rect 4020 12006 4032 12015
rect 4084 12006 4096 12015
rect 4148 12006 4160 12015
rect 4212 12006 4264 12058
rect 2774 11952 2816 11953
rect 2758 11944 2816 11952
rect 2758 11892 2769 11944
rect 2821 11892 2827 11944
rect 3118 11896 3157 11996
rect 3724 11962 4264 12006
rect 3741 11906 3787 11962
rect 3736 11905 3787 11906
rect 2758 11849 2816 11892
rect 2524 11777 2570 11815
rect 2524 11743 2530 11777
rect 2564 11743 2570 11777
rect 2524 11736 2570 11743
rect 2613 11797 2715 11825
rect 2613 11763 2647 11797
rect 2681 11763 2715 11797
rect 2524 11696 2574 11736
rect 2613 11735 2715 11763
rect 2758 11815 2776 11849
rect 2810 11815 2816 11849
rect 2758 11777 2816 11815
rect 2758 11743 2776 11777
rect 2810 11743 2816 11777
rect 1008 11636 1052 11690
rect 1245 11655 1328 11674
rect 852 11592 1052 11636
rect 1148 11653 1328 11655
rect 1148 11601 1155 11653
rect 1207 11643 1328 11653
rect 1207 11609 1269 11643
rect 1303 11609 1328 11643
rect 1207 11601 1328 11609
rect 1148 11600 1328 11601
rect 852 11470 896 11592
rect 1245 11579 1328 11600
rect 1568 11662 1602 11696
rect 1568 11652 1820 11662
rect 1568 11600 1758 11652
rect 1810 11600 1820 11652
rect 1568 11590 1820 11600
rect 1568 11558 1608 11590
rect 1853 11558 1892 11696
rect 2185 11558 2224 11696
rect 2255 11659 2325 11665
rect 2255 11650 2331 11659
rect 2255 11598 2270 11650
rect 2322 11598 2331 11650
rect 2255 11589 2331 11598
rect 2255 11583 2325 11589
rect 2368 11558 2407 11696
rect 2530 11662 2574 11696
rect 2758 11696 2816 11743
rect 2928 11849 2974 11896
rect 2928 11815 2934 11849
rect 2968 11836 2974 11849
rect 3114 11849 3160 11896
rect 3114 11836 3120 11849
rect 2968 11815 3120 11836
rect 3154 11815 3160 11849
rect 3272 11849 3318 11896
rect 3272 11839 3278 11849
rect 3312 11839 3318 11849
rect 3736 11859 3782 11905
rect 2928 11777 3160 11815
rect 3262 11787 3268 11839
rect 3320 11787 3326 11839
rect 3736 11825 3742 11859
rect 3776 11825 3782 11859
rect 3736 11787 3782 11825
rect 2928 11743 2934 11777
rect 2968 11743 3120 11777
rect 3154 11743 3160 11777
rect 2928 11726 3160 11743
rect 2928 11696 2974 11726
rect 3114 11696 3160 11726
rect 3272 11777 3318 11787
rect 3272 11743 3278 11777
rect 3312 11743 3318 11777
rect 3272 11696 3318 11743
rect 3736 11753 3742 11787
rect 3776 11753 3782 11787
rect 3736 11706 3782 11753
rect 3894 11859 3940 11906
rect 3894 11825 3900 11859
rect 3934 11825 3940 11859
rect 3894 11787 3940 11825
rect 3894 11753 3900 11787
rect 3934 11753 3940 11787
rect 3894 11706 3940 11753
rect 4044 11859 4090 11962
rect 4558 11906 4597 12112
rect 4738 12106 4744 12112
rect 4796 12106 4802 12158
rect 4868 11906 4907 12193
rect 5081 12199 7015 12229
rect 5029 12182 5081 12188
rect 6862 12151 6868 12158
rect 6516 12112 6868 12151
rect 5682 12058 6222 12102
rect 5682 12006 5734 12058
rect 5786 12048 5798 12058
rect 5850 12048 5862 12058
rect 5914 12048 5926 12058
rect 5978 12048 5990 12058
rect 6042 12048 6054 12058
rect 6106 12048 6118 12058
rect 5790 12014 5798 12048
rect 6042 12014 6044 12048
rect 6106 12014 6116 12048
rect 5786 12006 5798 12014
rect 5850 12006 5862 12014
rect 5914 12006 5926 12014
rect 5978 12006 5990 12014
rect 6042 12006 6054 12014
rect 6106 12006 6118 12014
rect 6170 12006 6222 12058
rect 5682 11962 6222 12006
rect 5700 11906 5746 11962
rect 4044 11825 4050 11859
rect 4084 11825 4090 11859
rect 4044 11787 4090 11825
rect 4044 11753 4050 11787
rect 4084 11753 4090 11787
rect 4044 11706 4090 11753
rect 4202 11859 4248 11906
rect 4202 11825 4208 11859
rect 4242 11825 4248 11859
rect 4396 11859 4442 11906
rect 4396 11833 4402 11859
rect 4202 11787 4248 11825
rect 4202 11753 4208 11787
rect 4242 11753 4248 11787
rect 4285 11831 4402 11833
rect 4285 11779 4292 11831
rect 4344 11825 4402 11831
rect 4436 11825 4442 11859
rect 4344 11787 4442 11825
rect 4344 11779 4402 11787
rect 4285 11778 4402 11779
rect 4202 11706 4248 11753
rect 4396 11753 4402 11778
rect 4436 11753 4442 11787
rect 4396 11706 4442 11753
rect 4554 11859 4600 11906
rect 4554 11825 4560 11859
rect 4594 11826 4600 11859
rect 4704 11859 4750 11906
rect 4704 11826 4710 11859
rect 4594 11825 4710 11826
rect 4744 11825 4750 11859
rect 4554 11787 4750 11825
rect 4554 11753 4560 11787
rect 4594 11760 4710 11787
rect 4594 11753 4600 11760
rect 4554 11706 4600 11753
rect 4704 11753 4710 11760
rect 4744 11753 4750 11787
rect 4704 11706 4750 11753
rect 4862 11859 4908 11906
rect 4862 11825 4868 11859
rect 4902 11825 4908 11859
rect 5694 11860 5740 11906
rect 5027 11830 5057 11839
rect 4862 11787 4908 11825
rect 4862 11753 4868 11787
rect 4902 11753 4908 11787
rect 5010 11778 5016 11830
rect 5068 11778 5074 11830
rect 5694 11826 5700 11860
rect 5734 11826 5740 11860
rect 5694 11788 5740 11826
rect 4862 11706 4908 11753
rect 5026 11737 5057 11778
rect 5694 11754 5700 11788
rect 5734 11754 5740 11788
rect 2758 11662 2802 11696
rect 2530 11618 2656 11662
rect 1242 11538 1248 11542
rect 1138 11494 1248 11538
rect 1138 11470 1182 11494
rect 1242 11490 1248 11494
rect 1300 11490 1306 11542
rect 1404 11525 1450 11558
rect 1404 11491 1410 11525
rect 1444 11491 1450 11525
rect 1404 11487 1450 11491
rect 378 11442 434 11448
rect 550 11442 622 11464
rect 434 11436 622 11442
rect 434 11396 565 11436
rect 606 11396 622 11436
rect 434 11386 622 11396
rect 378 11380 434 11386
rect 550 11366 622 11386
rect 696 11436 768 11464
rect 696 11396 712 11436
rect 753 11396 768 11436
rect 696 11366 768 11396
rect 840 11441 912 11470
rect 840 11401 856 11441
rect 897 11401 912 11441
rect 840 11372 912 11401
rect 994 11442 1182 11470
rect 994 11402 1010 11442
rect 1051 11426 1182 11442
rect 1399 11458 1450 11487
rect 1562 11525 1608 11558
rect 1562 11491 1568 11525
rect 1602 11491 1608 11525
rect 1692 11525 1738 11558
rect 1692 11496 1698 11525
rect 1562 11458 1608 11491
rect 1690 11491 1698 11496
rect 1732 11496 1738 11525
rect 1850 11525 1896 11558
rect 2024 11542 2070 11558
rect 1732 11491 1740 11496
rect 1051 11402 1066 11426
rect 1399 11412 1449 11458
rect 1690 11412 1740 11491
rect 1850 11491 1856 11525
rect 1890 11491 1896 11525
rect 1850 11458 1896 11491
rect 2014 11490 2020 11542
rect 2072 11490 2078 11542
rect 2182 11525 2228 11558
rect 2182 11491 2188 11525
rect 2222 11491 2228 11525
rect 2024 11458 2070 11490
rect 2182 11458 2228 11491
rect 2366 11525 2412 11558
rect 2524 11540 2570 11558
rect 2366 11491 2372 11525
rect 2406 11491 2412 11525
rect 2366 11458 2412 11491
rect 2516 11488 2522 11540
rect 2574 11488 2580 11540
rect 2524 11458 2570 11488
rect 2024 11426 2068 11458
rect 2612 11426 2656 11618
rect 994 11372 1066 11402
rect 1324 11357 1960 11412
rect 2024 11382 2656 11426
rect 2694 11618 2802 11662
rect 2832 11648 2904 11658
rect 2694 11420 2738 11618
rect 2832 11596 2842 11648
rect 2894 11596 2904 11648
rect 2832 11586 2904 11596
rect 2933 11558 2972 11696
rect 3118 11558 3157 11696
rect 3272 11652 3316 11696
rect 3268 11646 3320 11652
rect 3555 11621 3561 11673
rect 3613 11666 3619 11673
rect 3662 11666 3713 11678
rect 3613 11663 3713 11666
rect 3613 11629 3670 11663
rect 3704 11629 3713 11663
rect 3613 11627 3713 11629
rect 3613 11621 3619 11627
rect 3662 11615 3713 11627
rect 3897 11657 3936 11706
rect 3976 11664 4027 11669
rect 3970 11657 3976 11664
rect 3897 11618 3976 11657
rect 3268 11588 3320 11594
rect 3897 11568 3936 11618
rect 3970 11612 3976 11618
rect 4028 11612 4034 11664
rect 4206 11650 4245 11706
rect 4300 11650 4347 11661
rect 4206 11648 4347 11650
rect 4206 11615 4306 11648
rect 3976 11606 4027 11612
rect 4206 11568 4245 11615
rect 4300 11614 4306 11615
rect 4340 11614 4347 11648
rect 4300 11602 4347 11614
rect 2766 11552 2818 11558
rect 2766 11494 2776 11500
rect 2770 11491 2776 11494
rect 2810 11494 2818 11500
rect 2928 11525 2974 11558
rect 2810 11491 2816 11494
rect 2770 11458 2816 11491
rect 2928 11491 2934 11525
rect 2968 11491 2974 11525
rect 2928 11458 2974 11491
rect 3114 11525 3160 11558
rect 3114 11491 3120 11525
rect 3154 11491 3160 11525
rect 3114 11458 3160 11491
rect 3272 11525 3318 11558
rect 3272 11491 3278 11525
rect 3312 11491 3318 11525
rect 3272 11458 3318 11491
rect 3274 11420 3318 11458
rect 2694 11376 3318 11420
rect 3736 11535 3782 11568
rect 3736 11501 3742 11535
rect 3776 11501 3782 11535
rect 3736 11468 3782 11501
rect 3894 11535 3940 11568
rect 3894 11501 3900 11535
rect 3934 11501 3940 11535
rect 4044 11535 4090 11568
rect 4044 11506 4050 11535
rect 3894 11468 3940 11501
rect 4042 11501 4050 11506
rect 4084 11501 4090 11535
rect 4042 11468 4090 11501
rect 4202 11535 4248 11568
rect 4202 11501 4208 11535
rect 4242 11501 4248 11535
rect 4202 11468 4248 11501
rect 3736 11412 3780 11468
rect 4042 11412 4089 11468
rect 1324 11305 1360 11357
rect 1412 11305 1424 11357
rect 1476 11348 1488 11357
rect 1540 11348 1552 11357
rect 1604 11348 1616 11357
rect 1668 11348 1680 11357
rect 1732 11348 1744 11357
rect 1796 11348 1808 11357
rect 1479 11314 1488 11348
rect 1551 11314 1552 11348
rect 1732 11314 1733 11348
rect 1796 11314 1805 11348
rect 1476 11305 1488 11314
rect 1540 11305 1552 11314
rect 1604 11305 1616 11314
rect 1668 11305 1680 11314
rect 1732 11305 1744 11314
rect 1796 11305 1808 11314
rect 1860 11305 1872 11357
rect 1924 11305 1960 11357
rect 3704 11368 4244 11412
rect 3704 11359 3756 11368
rect 3808 11359 3820 11368
rect 1324 11272 1960 11305
rect 2346 11327 2426 11352
rect 2346 11323 3517 11327
rect 2346 11289 2369 11323
rect 2403 11289 3517 11323
rect 2346 11285 3517 11289
rect 2346 11260 2426 11285
rect 2636 11227 2702 11239
rect 272 11173 278 11227
rect 332 11173 2642 11227
rect 2696 11173 2702 11227
rect 2636 11161 2702 11173
rect 3475 11132 3517 11285
rect 3704 11325 3741 11359
rect 3808 11325 3813 11359
rect 3704 11316 3756 11325
rect 3808 11316 3820 11325
rect 3872 11316 3884 11368
rect 3936 11316 3948 11368
rect 4000 11316 4012 11368
rect 4064 11316 4076 11368
rect 4128 11359 4140 11368
rect 4192 11359 4244 11368
rect 4135 11325 4140 11359
rect 4207 11325 4244 11359
rect 4128 11316 4140 11325
rect 4192 11316 4244 11325
rect 3704 11272 4244 11316
rect 3559 11167 3565 11219
rect 3617 11212 3623 11219
rect 4306 11212 4345 11602
rect 4558 11570 4597 11706
rect 4628 11675 4680 11681
rect 4625 11626 4628 11672
rect 4680 11626 4683 11672
rect 4875 11630 4904 11706
rect 4628 11617 4680 11623
rect 4875 11602 4980 11630
rect 4396 11537 4442 11570
rect 4396 11503 4402 11537
rect 4436 11503 4442 11537
rect 4396 11470 4442 11503
rect 4554 11550 4600 11570
rect 4704 11550 4750 11570
rect 4862 11550 4908 11570
rect 4554 11537 4750 11550
rect 4554 11503 4560 11537
rect 4594 11503 4710 11537
rect 4744 11503 4750 11537
rect 4554 11484 4750 11503
rect 4856 11498 4862 11550
rect 4914 11498 4920 11550
rect 4554 11470 4600 11484
rect 4704 11470 4750 11484
rect 4862 11470 4908 11498
rect 4402 11320 4430 11470
rect 4558 11425 4597 11470
rect 4552 11419 4604 11425
rect 4552 11361 4604 11367
rect 4952 11320 4980 11602
rect 5026 11552 5056 11737
rect 5694 11706 5740 11754
rect 5852 11860 5898 11906
rect 5852 11826 5858 11860
rect 5892 11826 5898 11860
rect 5852 11788 5898 11826
rect 5852 11754 5858 11788
rect 5892 11754 5898 11788
rect 5852 11706 5898 11754
rect 6002 11860 6048 11962
rect 6516 11906 6556 12112
rect 6862 12106 6868 12112
rect 6920 12106 6926 12158
rect 6985 12146 7015 12199
rect 6985 12117 7016 12146
rect 6002 11826 6008 11860
rect 6042 11826 6048 11860
rect 6002 11788 6048 11826
rect 6002 11754 6008 11788
rect 6042 11754 6048 11788
rect 6002 11706 6048 11754
rect 6160 11860 6206 11906
rect 6160 11826 6166 11860
rect 6200 11826 6206 11860
rect 6354 11860 6400 11906
rect 6354 11834 6360 11860
rect 6160 11788 6206 11826
rect 6160 11754 6166 11788
rect 6200 11754 6206 11788
rect 6244 11832 6360 11834
rect 6244 11780 6250 11832
rect 6302 11826 6360 11832
rect 6394 11826 6400 11860
rect 6302 11788 6400 11826
rect 6302 11780 6360 11788
rect 6244 11778 6360 11780
rect 6160 11706 6206 11754
rect 6354 11754 6360 11778
rect 6394 11754 6400 11788
rect 6354 11706 6400 11754
rect 6512 11860 6558 11906
rect 6512 11826 6518 11860
rect 6552 11826 6558 11860
rect 6662 11860 6708 11906
rect 6662 11826 6668 11860
rect 6702 11826 6708 11860
rect 6512 11788 6708 11826
rect 6512 11754 6518 11788
rect 6552 11760 6668 11788
rect 6552 11754 6558 11760
rect 6512 11706 6558 11754
rect 6662 11754 6668 11760
rect 6702 11754 6708 11788
rect 6662 11706 6708 11754
rect 6820 11860 6866 11906
rect 6820 11826 6826 11860
rect 6860 11826 6866 11860
rect 6986 11830 7016 12117
rect 6820 11788 6866 11826
rect 6820 11754 6826 11788
rect 6860 11754 6866 11788
rect 6968 11778 6974 11830
rect 7026 11778 7032 11830
rect 6820 11706 6866 11754
rect 6984 11738 7016 11778
rect 5111 11621 5117 11673
rect 5169 11666 5175 11673
rect 5620 11666 5672 11678
rect 5169 11664 5672 11666
rect 5169 11630 5628 11664
rect 5662 11630 5672 11664
rect 5169 11627 5672 11630
rect 5169 11621 5175 11627
rect 5620 11616 5672 11627
rect 5856 11658 5894 11706
rect 5934 11664 5986 11670
rect 5928 11658 5934 11664
rect 5856 11618 5934 11658
rect 5856 11568 5894 11618
rect 5928 11612 5934 11618
rect 5986 11612 5992 11664
rect 6164 11650 6204 11706
rect 6258 11650 6306 11662
rect 6164 11648 6306 11650
rect 6164 11616 6264 11648
rect 5934 11606 5986 11612
rect 6164 11568 6204 11616
rect 6258 11614 6264 11616
rect 6298 11614 6306 11648
rect 6258 11602 6306 11614
rect 5009 11500 5015 11552
rect 5067 11500 5073 11552
rect 5694 11536 5740 11568
rect 5694 11502 5700 11536
rect 5734 11502 5740 11536
rect 4402 11292 4980 11320
rect 3617 11173 4345 11212
rect 3617 11167 3623 11173
rect 5021 11132 5063 11500
rect 5694 11468 5740 11502
rect 5852 11536 5898 11568
rect 5852 11502 5858 11536
rect 5892 11502 5898 11536
rect 6002 11536 6048 11568
rect 6002 11506 6008 11536
rect 5852 11468 5898 11502
rect 6000 11502 6008 11506
rect 6042 11502 6048 11536
rect 5694 11412 5738 11468
rect 6000 11412 6048 11502
rect 6160 11536 6206 11568
rect 6160 11502 6166 11536
rect 6200 11502 6206 11536
rect 6160 11468 6206 11502
rect 5662 11368 6202 11412
rect 5662 11360 5714 11368
rect 5766 11360 5778 11368
rect 5662 11326 5700 11360
rect 5766 11326 5772 11360
rect 5662 11316 5714 11326
rect 5766 11316 5778 11326
rect 5830 11316 5842 11368
rect 5894 11316 5906 11368
rect 5958 11316 5970 11368
rect 6022 11316 6034 11368
rect 6086 11360 6098 11368
rect 6150 11360 6202 11368
rect 6094 11326 6098 11360
rect 6166 11326 6202 11360
rect 6086 11316 6098 11326
rect 6150 11316 6202 11326
rect 5662 11272 6202 11316
rect 5111 11167 5117 11219
rect 5169 11212 5175 11219
rect 6264 11212 6304 11602
rect 6516 11570 6556 11706
rect 6586 11676 6638 11682
rect 6584 11626 6586 11672
rect 6638 11626 6642 11672
rect 6834 11630 6862 11706
rect 6586 11618 6638 11624
rect 6834 11602 6936 11630
rect 6354 11538 6400 11570
rect 6354 11504 6360 11538
rect 6394 11504 6400 11538
rect 6354 11470 6400 11504
rect 6512 11550 6558 11570
rect 6662 11550 6708 11570
rect 6820 11550 6866 11570
rect 6512 11538 6708 11550
rect 6512 11504 6518 11538
rect 6552 11504 6668 11538
rect 6702 11504 6708 11538
rect 6512 11484 6708 11504
rect 6814 11498 6820 11550
rect 6872 11498 6878 11550
rect 6512 11470 6558 11484
rect 6662 11470 6708 11484
rect 6820 11470 6866 11498
rect 6360 11320 6388 11470
rect 6516 11426 6556 11470
rect 6510 11420 6562 11426
rect 6510 11362 6562 11368
rect 6908 11320 6936 11602
rect 6984 11552 7014 11738
rect 6968 11500 6974 11552
rect 7026 11500 7032 11552
rect 6360 11292 6936 11320
rect 6908 11228 6936 11292
rect 5169 11174 6304 11212
rect 6346 11200 6936 11228
rect 5169 11173 5572 11174
rect 5169 11167 5175 11173
rect 3475 11090 5063 11132
rect 5035 11049 5087 11055
rect 3472 10965 4907 11004
rect 6346 11037 6374 11200
rect 6908 11198 6936 11200
rect 5087 11009 6374 11037
rect 5035 10991 5087 10997
rect 6968 10970 6974 11022
rect 7026 10970 7032 11022
rect 1348 10831 1880 10874
rect 1348 10822 1398 10831
rect 1450 10822 1462 10831
rect 1348 10788 1383 10822
rect 1450 10788 1455 10822
rect 1348 10779 1398 10788
rect 1450 10779 1462 10788
rect 1514 10779 1526 10831
rect 1578 10779 1590 10831
rect 1642 10779 1654 10831
rect 1706 10779 1718 10831
rect 1770 10822 1782 10831
rect 1834 10822 1880 10831
rect 1777 10788 1782 10822
rect 1849 10788 1880 10822
rect 3472 10807 3511 10965
rect 4738 10923 4744 10930
rect 4558 10884 4744 10923
rect 1770 10779 1782 10788
rect 1834 10779 1880 10788
rect 550 10760 622 10764
rect 550 10708 560 10760
rect 612 10708 622 10760
rect 696 10758 768 10764
rect 550 10696 566 10708
rect 607 10696 622 10708
rect 682 10756 768 10758
rect 682 10704 702 10756
rect 754 10704 768 10756
rect 682 10702 710 10704
rect 550 10666 622 10696
rect 696 10696 710 10702
rect 751 10696 768 10704
rect 696 10666 768 10696
rect 840 10741 912 10770
rect 840 10701 856 10741
rect 897 10701 912 10741
rect 840 10672 912 10701
rect 994 10741 1066 10770
rect 994 10701 1009 10741
rect 1050 10701 1066 10741
rect 1348 10734 1880 10779
rect 994 10672 1066 10701
rect 564 10626 608 10666
rect 856 10606 900 10672
rect 378 10598 433 10604
rect 846 10554 852 10606
rect 904 10554 910 10606
rect 378 10313 433 10543
rect 856 10514 900 10554
rect 1008 10514 1052 10672
rect 1407 10668 1448 10734
rect 1693 10668 1735 10734
rect 1941 10731 2687 10776
rect 1404 10621 1450 10668
rect 1404 10587 1410 10621
rect 1444 10587 1450 10621
rect 1404 10549 1450 10587
rect 1404 10515 1410 10549
rect 1444 10515 1450 10549
rect 708 10470 900 10514
rect 372 10258 378 10313
rect 433 10258 439 10313
rect 708 10236 752 10470
rect 998 10462 1004 10514
rect 1056 10462 1062 10514
rect 1404 10468 1450 10515
rect 1562 10621 1608 10668
rect 1562 10587 1568 10621
rect 1602 10587 1608 10621
rect 1562 10549 1608 10587
rect 1562 10515 1568 10549
rect 1602 10515 1608 10549
rect 1562 10468 1608 10515
rect 1692 10621 1738 10668
rect 1692 10587 1698 10621
rect 1732 10587 1738 10621
rect 1692 10549 1738 10587
rect 1692 10515 1698 10549
rect 1732 10515 1738 10549
rect 1692 10468 1738 10515
rect 1850 10665 1896 10668
rect 1941 10665 1986 10731
rect 1850 10621 1986 10665
rect 1850 10587 1856 10621
rect 1890 10620 1986 10621
rect 2024 10621 2070 10668
rect 1890 10587 1896 10620
rect 1850 10549 1896 10587
rect 2024 10587 2030 10621
rect 2064 10587 2070 10621
rect 2024 10552 2070 10587
rect 1998 10550 2070 10552
rect 1850 10515 1856 10549
rect 1890 10515 1896 10549
rect 1850 10468 1896 10515
rect 1928 10549 2070 10550
rect 1928 10525 2030 10549
rect 1928 10508 1935 10525
rect 1929 10473 1935 10508
rect 1987 10515 2030 10525
rect 2064 10515 2070 10549
rect 1987 10508 2070 10515
rect 1987 10473 1993 10508
rect 2024 10468 2070 10508
rect 2182 10624 2228 10668
rect 2366 10624 2412 10668
rect 2182 10621 2412 10624
rect 2182 10587 2188 10621
rect 2222 10587 2372 10621
rect 2406 10587 2412 10621
rect 2182 10549 2412 10587
rect 2182 10515 2188 10549
rect 2222 10515 2372 10549
rect 2406 10515 2412 10549
rect 2182 10498 2412 10515
rect 2182 10468 2228 10498
rect 2366 10468 2412 10498
rect 2524 10621 2570 10668
rect 2524 10587 2530 10621
rect 2564 10587 2570 10621
rect 2642 10597 2687 10731
rect 3118 10768 3511 10807
rect 3724 10830 4264 10874
rect 3724 10778 3776 10830
rect 3828 10821 3840 10830
rect 3892 10821 3904 10830
rect 3956 10821 3968 10830
rect 4020 10821 4032 10830
rect 4084 10821 4096 10830
rect 4148 10821 4160 10830
rect 3831 10787 3840 10821
rect 3903 10787 3904 10821
rect 4084 10787 4085 10821
rect 4148 10787 4157 10821
rect 3828 10778 3840 10787
rect 3892 10778 3904 10787
rect 3956 10778 3968 10787
rect 4020 10778 4032 10787
rect 4084 10778 4096 10787
rect 4148 10778 4160 10787
rect 4212 10778 4264 10830
rect 2774 10724 2816 10725
rect 2758 10716 2816 10724
rect 2758 10664 2769 10716
rect 2821 10664 2827 10716
rect 3118 10668 3157 10768
rect 3724 10734 4264 10778
rect 3741 10678 3787 10734
rect 3736 10677 3787 10678
rect 2758 10621 2816 10664
rect 2524 10549 2570 10587
rect 2524 10515 2530 10549
rect 2564 10515 2570 10549
rect 2524 10508 2570 10515
rect 2613 10569 2715 10597
rect 2613 10535 2647 10569
rect 2681 10535 2715 10569
rect 2524 10468 2574 10508
rect 2613 10507 2715 10535
rect 2758 10587 2776 10621
rect 2810 10587 2816 10621
rect 2758 10549 2816 10587
rect 2758 10515 2776 10549
rect 2810 10515 2816 10549
rect 1008 10408 1052 10462
rect 1245 10427 1328 10446
rect 852 10364 1052 10408
rect 1148 10425 1328 10427
rect 1148 10373 1155 10425
rect 1207 10415 1328 10425
rect 1207 10381 1269 10415
rect 1303 10381 1328 10415
rect 1207 10373 1328 10381
rect 1148 10372 1328 10373
rect 852 10242 896 10364
rect 1245 10351 1328 10372
rect 1568 10434 1602 10468
rect 1568 10424 1820 10434
rect 1568 10372 1758 10424
rect 1810 10372 1820 10424
rect 1568 10362 1820 10372
rect 1568 10330 1608 10362
rect 1853 10330 1892 10468
rect 2185 10330 2224 10468
rect 2255 10431 2325 10437
rect 2255 10422 2331 10431
rect 2255 10370 2270 10422
rect 2322 10370 2331 10422
rect 2255 10361 2331 10370
rect 2255 10355 2325 10361
rect 2368 10330 2407 10468
rect 2530 10434 2574 10468
rect 2758 10468 2816 10515
rect 2928 10621 2974 10668
rect 2928 10587 2934 10621
rect 2968 10608 2974 10621
rect 3114 10621 3160 10668
rect 3114 10608 3120 10621
rect 2968 10587 3120 10608
rect 3154 10587 3160 10621
rect 3272 10621 3318 10668
rect 3272 10611 3278 10621
rect 3312 10611 3318 10621
rect 3736 10631 3782 10677
rect 2928 10549 3160 10587
rect 3262 10559 3268 10611
rect 3320 10559 3326 10611
rect 3736 10597 3742 10631
rect 3776 10597 3782 10631
rect 3736 10559 3782 10597
rect 2928 10515 2934 10549
rect 2968 10515 3120 10549
rect 3154 10515 3160 10549
rect 2928 10498 3160 10515
rect 2928 10468 2974 10498
rect 3114 10468 3160 10498
rect 3272 10549 3318 10559
rect 3272 10515 3278 10549
rect 3312 10515 3318 10549
rect 3272 10468 3318 10515
rect 3736 10525 3742 10559
rect 3776 10525 3782 10559
rect 3736 10478 3782 10525
rect 3894 10631 3940 10678
rect 3894 10597 3900 10631
rect 3934 10597 3940 10631
rect 3894 10559 3940 10597
rect 3894 10525 3900 10559
rect 3934 10525 3940 10559
rect 3894 10478 3940 10525
rect 4044 10631 4090 10734
rect 4558 10678 4597 10884
rect 4738 10878 4744 10884
rect 4796 10878 4802 10930
rect 4868 10678 4907 10965
rect 6829 10923 6835 10930
rect 6516 10884 6835 10923
rect 5682 10830 6222 10874
rect 5682 10778 5734 10830
rect 5786 10820 5798 10830
rect 5850 10820 5862 10830
rect 5914 10820 5926 10830
rect 5978 10820 5990 10830
rect 6042 10820 6054 10830
rect 6106 10820 6118 10830
rect 5790 10786 5798 10820
rect 6042 10786 6044 10820
rect 6106 10786 6116 10820
rect 5786 10778 5798 10786
rect 5850 10778 5862 10786
rect 5914 10778 5926 10786
rect 5978 10778 5990 10786
rect 6042 10778 6054 10786
rect 6106 10778 6118 10786
rect 6170 10778 6222 10830
rect 5682 10734 6222 10778
rect 5700 10678 5746 10734
rect 4044 10597 4050 10631
rect 4084 10597 4090 10631
rect 4044 10559 4090 10597
rect 4044 10525 4050 10559
rect 4084 10525 4090 10559
rect 4044 10478 4090 10525
rect 4202 10631 4248 10678
rect 4202 10597 4208 10631
rect 4242 10597 4248 10631
rect 4396 10631 4442 10678
rect 4396 10605 4402 10631
rect 4202 10559 4248 10597
rect 4202 10525 4208 10559
rect 4242 10525 4248 10559
rect 4285 10603 4402 10605
rect 4285 10551 4292 10603
rect 4344 10597 4402 10603
rect 4436 10597 4442 10631
rect 4344 10559 4442 10597
rect 4344 10551 4402 10559
rect 4285 10550 4402 10551
rect 4202 10478 4248 10525
rect 4396 10525 4402 10550
rect 4436 10525 4442 10559
rect 4396 10478 4442 10525
rect 4554 10631 4600 10678
rect 4554 10597 4560 10631
rect 4594 10598 4600 10631
rect 4704 10631 4750 10678
rect 4704 10598 4710 10631
rect 4594 10597 4710 10598
rect 4744 10597 4750 10631
rect 4554 10559 4750 10597
rect 4554 10525 4560 10559
rect 4594 10532 4710 10559
rect 4594 10525 4600 10532
rect 4554 10478 4600 10525
rect 4704 10525 4710 10532
rect 4744 10525 4750 10559
rect 4704 10478 4750 10525
rect 4862 10631 4908 10678
rect 4862 10597 4868 10631
rect 4902 10597 4908 10631
rect 5694 10632 5740 10678
rect 5027 10602 5057 10611
rect 4862 10559 4908 10597
rect 4862 10525 4868 10559
rect 4902 10525 4908 10559
rect 5010 10550 5016 10602
rect 5068 10550 5074 10602
rect 5694 10598 5700 10632
rect 5734 10598 5740 10632
rect 5694 10560 5740 10598
rect 4862 10478 4908 10525
rect 5026 10509 5057 10550
rect 5694 10526 5700 10560
rect 5734 10526 5740 10560
rect 2758 10434 2802 10468
rect 2530 10390 2656 10434
rect 1242 10310 1248 10314
rect 1138 10266 1248 10310
rect 1138 10242 1182 10266
rect 1242 10262 1248 10266
rect 1300 10262 1306 10314
rect 1404 10297 1450 10330
rect 1404 10263 1410 10297
rect 1444 10263 1450 10297
rect 1404 10259 1450 10263
rect 378 10214 434 10220
rect 550 10214 622 10236
rect 434 10208 622 10214
rect 434 10168 565 10208
rect 606 10168 622 10208
rect 434 10158 622 10168
rect 378 10152 434 10158
rect 550 10138 622 10158
rect 696 10208 768 10236
rect 696 10168 712 10208
rect 753 10168 768 10208
rect 696 10138 768 10168
rect 840 10213 912 10242
rect 840 10173 856 10213
rect 897 10173 912 10213
rect 840 10144 912 10173
rect 994 10214 1182 10242
rect 994 10174 1010 10214
rect 1051 10198 1182 10214
rect 1399 10230 1450 10259
rect 1562 10297 1608 10330
rect 1562 10263 1568 10297
rect 1602 10263 1608 10297
rect 1692 10297 1738 10330
rect 1692 10268 1698 10297
rect 1562 10230 1608 10263
rect 1690 10263 1698 10268
rect 1732 10268 1738 10297
rect 1850 10297 1896 10330
rect 2024 10314 2070 10330
rect 1732 10263 1740 10268
rect 1051 10174 1066 10198
rect 1399 10184 1449 10230
rect 1690 10184 1740 10263
rect 1850 10263 1856 10297
rect 1890 10263 1896 10297
rect 1850 10230 1896 10263
rect 2014 10262 2020 10314
rect 2072 10262 2078 10314
rect 2182 10297 2228 10330
rect 2182 10263 2188 10297
rect 2222 10263 2228 10297
rect 2024 10230 2070 10262
rect 2182 10230 2228 10263
rect 2366 10297 2412 10330
rect 2524 10312 2570 10330
rect 2366 10263 2372 10297
rect 2406 10263 2412 10297
rect 2366 10230 2412 10263
rect 2516 10260 2522 10312
rect 2574 10260 2580 10312
rect 2524 10230 2570 10260
rect 2024 10198 2068 10230
rect 2612 10198 2656 10390
rect 994 10144 1066 10174
rect 1324 10129 1960 10184
rect 2024 10154 2656 10198
rect 2694 10390 2802 10434
rect 2832 10420 2904 10430
rect 2694 10192 2738 10390
rect 2832 10368 2842 10420
rect 2894 10368 2904 10420
rect 2832 10358 2904 10368
rect 2933 10330 2972 10468
rect 3118 10330 3157 10468
rect 3272 10424 3316 10468
rect 3268 10418 3320 10424
rect 3555 10393 3561 10445
rect 3613 10438 3619 10445
rect 3662 10438 3713 10450
rect 3613 10435 3713 10438
rect 3613 10401 3670 10435
rect 3704 10401 3713 10435
rect 3613 10399 3713 10401
rect 3613 10393 3619 10399
rect 3662 10387 3713 10399
rect 3897 10429 3936 10478
rect 3976 10436 4027 10441
rect 3970 10429 3976 10436
rect 3897 10390 3976 10429
rect 3268 10360 3320 10366
rect 3897 10340 3936 10390
rect 3970 10384 3976 10390
rect 4028 10384 4034 10436
rect 4206 10422 4245 10478
rect 4300 10422 4347 10433
rect 4206 10420 4347 10422
rect 4206 10387 4306 10420
rect 3976 10378 4027 10384
rect 4206 10340 4245 10387
rect 4300 10386 4306 10387
rect 4340 10386 4347 10420
rect 4300 10374 4347 10386
rect 2766 10324 2818 10330
rect 2766 10266 2776 10272
rect 2770 10263 2776 10266
rect 2810 10266 2818 10272
rect 2928 10297 2974 10330
rect 2810 10263 2816 10266
rect 2770 10230 2816 10263
rect 2928 10263 2934 10297
rect 2968 10263 2974 10297
rect 2928 10230 2974 10263
rect 3114 10297 3160 10330
rect 3114 10263 3120 10297
rect 3154 10263 3160 10297
rect 3114 10230 3160 10263
rect 3272 10297 3318 10330
rect 3272 10263 3278 10297
rect 3312 10263 3318 10297
rect 3272 10230 3318 10263
rect 3274 10192 3318 10230
rect 2694 10148 3318 10192
rect 3736 10307 3782 10340
rect 3736 10273 3742 10307
rect 3776 10273 3782 10307
rect 3736 10240 3782 10273
rect 3894 10307 3940 10340
rect 3894 10273 3900 10307
rect 3934 10273 3940 10307
rect 4044 10307 4090 10340
rect 4044 10278 4050 10307
rect 3894 10240 3940 10273
rect 4042 10273 4050 10278
rect 4084 10273 4090 10307
rect 4042 10240 4090 10273
rect 4202 10307 4248 10340
rect 4202 10273 4208 10307
rect 4242 10273 4248 10307
rect 4202 10240 4248 10273
rect 3736 10184 3780 10240
rect 4042 10184 4089 10240
rect 1324 10077 1360 10129
rect 1412 10077 1424 10129
rect 1476 10120 1488 10129
rect 1540 10120 1552 10129
rect 1604 10120 1616 10129
rect 1668 10120 1680 10129
rect 1732 10120 1744 10129
rect 1796 10120 1808 10129
rect 1479 10086 1488 10120
rect 1551 10086 1552 10120
rect 1732 10086 1733 10120
rect 1796 10086 1805 10120
rect 1476 10077 1488 10086
rect 1540 10077 1552 10086
rect 1604 10077 1616 10086
rect 1668 10077 1680 10086
rect 1732 10077 1744 10086
rect 1796 10077 1808 10086
rect 1860 10077 1872 10129
rect 1924 10077 1960 10129
rect 3704 10140 4244 10184
rect 3704 10131 3756 10140
rect 3808 10131 3820 10140
rect 1324 10044 1960 10077
rect 2346 10099 2426 10124
rect 2346 10095 3517 10099
rect 2346 10061 2369 10095
rect 2403 10061 3517 10095
rect 2346 10057 3517 10061
rect 2346 10032 2426 10057
rect 2636 9999 2702 10011
rect 272 9945 278 9999
rect 332 9945 2642 9999
rect 2696 9945 2702 9999
rect 2636 9933 2702 9945
rect 3475 9904 3517 10057
rect 3704 10097 3741 10131
rect 3808 10097 3813 10131
rect 3704 10088 3756 10097
rect 3808 10088 3820 10097
rect 3872 10088 3884 10140
rect 3936 10088 3948 10140
rect 4000 10088 4012 10140
rect 4064 10088 4076 10140
rect 4128 10131 4140 10140
rect 4192 10131 4244 10140
rect 4135 10097 4140 10131
rect 4207 10097 4244 10131
rect 4128 10088 4140 10097
rect 4192 10088 4244 10097
rect 3704 10044 4244 10088
rect 3559 9939 3565 9991
rect 3617 9984 3623 9991
rect 4306 9984 4345 10374
rect 4558 10342 4597 10478
rect 4628 10447 4680 10453
rect 4625 10398 4628 10444
rect 4680 10398 4683 10444
rect 4875 10402 4904 10478
rect 4628 10389 4680 10395
rect 4875 10374 4980 10402
rect 4396 10309 4442 10342
rect 4396 10275 4402 10309
rect 4436 10275 4442 10309
rect 4396 10242 4442 10275
rect 4554 10322 4600 10342
rect 4704 10322 4750 10342
rect 4862 10322 4908 10342
rect 4554 10309 4750 10322
rect 4554 10275 4560 10309
rect 4594 10275 4710 10309
rect 4744 10275 4750 10309
rect 4554 10256 4750 10275
rect 4856 10270 4862 10322
rect 4914 10270 4920 10322
rect 4554 10242 4600 10256
rect 4704 10242 4750 10256
rect 4862 10242 4908 10270
rect 4402 10092 4430 10242
rect 4558 10197 4597 10242
rect 4552 10191 4604 10197
rect 4552 10133 4604 10139
rect 4952 10092 4980 10374
rect 5026 10324 5056 10509
rect 5694 10478 5740 10526
rect 5852 10632 5898 10678
rect 5852 10598 5858 10632
rect 5892 10598 5898 10632
rect 5852 10560 5898 10598
rect 5852 10526 5858 10560
rect 5892 10526 5898 10560
rect 5852 10478 5898 10526
rect 6002 10632 6048 10734
rect 6516 10678 6556 10884
rect 6829 10878 6835 10884
rect 6887 10878 6893 10930
rect 6985 10918 7015 10970
rect 6985 10889 7016 10918
rect 6002 10598 6008 10632
rect 6042 10598 6048 10632
rect 6002 10560 6048 10598
rect 6002 10526 6008 10560
rect 6042 10526 6048 10560
rect 6002 10478 6048 10526
rect 6160 10632 6206 10678
rect 6160 10598 6166 10632
rect 6200 10598 6206 10632
rect 6354 10632 6400 10678
rect 6354 10606 6360 10632
rect 6160 10560 6206 10598
rect 6160 10526 6166 10560
rect 6200 10526 6206 10560
rect 6244 10604 6360 10606
rect 6244 10552 6250 10604
rect 6302 10598 6360 10604
rect 6394 10598 6400 10632
rect 6302 10560 6400 10598
rect 6302 10552 6360 10560
rect 6244 10550 6360 10552
rect 6160 10478 6206 10526
rect 6354 10526 6360 10550
rect 6394 10526 6400 10560
rect 6354 10478 6400 10526
rect 6512 10632 6558 10678
rect 6512 10598 6518 10632
rect 6552 10598 6558 10632
rect 6662 10632 6708 10678
rect 6662 10598 6668 10632
rect 6702 10598 6708 10632
rect 6512 10560 6708 10598
rect 6512 10526 6518 10560
rect 6552 10532 6668 10560
rect 6552 10526 6558 10532
rect 6512 10478 6558 10526
rect 6662 10526 6668 10532
rect 6702 10526 6708 10560
rect 6662 10478 6708 10526
rect 6820 10632 6866 10678
rect 6820 10598 6826 10632
rect 6860 10598 6866 10632
rect 6986 10602 7016 10889
rect 6820 10560 6866 10598
rect 6820 10526 6826 10560
rect 6860 10526 6866 10560
rect 6968 10550 6974 10602
rect 7026 10550 7032 10602
rect 6820 10478 6866 10526
rect 6984 10510 7016 10550
rect 5350 10393 5356 10445
rect 5408 10438 5414 10445
rect 5620 10438 5672 10450
rect 5408 10436 5672 10438
rect 5408 10402 5628 10436
rect 5662 10402 5672 10436
rect 5408 10399 5672 10402
rect 5408 10393 5414 10399
rect 5620 10388 5672 10399
rect 5856 10430 5894 10478
rect 5934 10436 5986 10442
rect 5928 10430 5934 10436
rect 5856 10390 5934 10430
rect 5856 10340 5894 10390
rect 5928 10384 5934 10390
rect 5986 10384 5992 10436
rect 6164 10422 6204 10478
rect 6258 10422 6306 10434
rect 6164 10420 6306 10422
rect 6164 10388 6264 10420
rect 5934 10378 5986 10384
rect 6164 10340 6204 10388
rect 6258 10386 6264 10388
rect 6298 10386 6306 10420
rect 6258 10374 6306 10386
rect 5009 10272 5015 10324
rect 5067 10272 5073 10324
rect 5694 10308 5740 10340
rect 5694 10274 5700 10308
rect 5734 10274 5740 10308
rect 4402 10064 4980 10092
rect 3617 9945 4345 9984
rect 3617 9939 3623 9945
rect 5021 9904 5063 10272
rect 5694 10240 5740 10274
rect 5852 10308 5898 10340
rect 5852 10274 5858 10308
rect 5892 10274 5898 10308
rect 6002 10308 6048 10340
rect 6002 10278 6008 10308
rect 5852 10240 5898 10274
rect 6000 10274 6008 10278
rect 6042 10274 6048 10308
rect 5694 10184 5738 10240
rect 6000 10184 6048 10274
rect 6160 10308 6206 10340
rect 6160 10274 6166 10308
rect 6200 10274 6206 10308
rect 6160 10240 6206 10274
rect 5662 10140 6202 10184
rect 5662 10132 5714 10140
rect 5766 10132 5778 10140
rect 5662 10098 5700 10132
rect 5766 10098 5772 10132
rect 5662 10088 5714 10098
rect 5766 10088 5778 10098
rect 5830 10088 5842 10140
rect 5894 10088 5906 10140
rect 5958 10088 5970 10140
rect 6022 10088 6034 10140
rect 6086 10132 6098 10140
rect 6150 10132 6202 10140
rect 6094 10098 6098 10132
rect 6166 10098 6202 10132
rect 6086 10088 6098 10098
rect 6150 10088 6202 10098
rect 5662 10044 6202 10088
rect 5348 9939 5354 9991
rect 5406 9984 5412 9991
rect 6264 9984 6304 10374
rect 6516 10342 6556 10478
rect 6586 10448 6638 10454
rect 6584 10398 6586 10444
rect 6638 10398 6642 10444
rect 6834 10402 6862 10478
rect 6586 10390 6638 10396
rect 6834 10374 6936 10402
rect 6354 10310 6400 10342
rect 6354 10276 6360 10310
rect 6394 10276 6400 10310
rect 6354 10242 6400 10276
rect 6512 10322 6558 10342
rect 6662 10322 6708 10342
rect 6820 10322 6866 10342
rect 6512 10310 6708 10322
rect 6512 10276 6518 10310
rect 6552 10276 6668 10310
rect 6702 10276 6708 10310
rect 6512 10256 6708 10276
rect 6814 10270 6820 10322
rect 6872 10270 6878 10322
rect 6512 10242 6558 10256
rect 6662 10242 6708 10256
rect 6820 10242 6866 10270
rect 6360 10092 6388 10242
rect 6516 10198 6556 10242
rect 6510 10192 6562 10198
rect 6510 10134 6562 10140
rect 6908 10092 6936 10374
rect 6984 10324 7014 10510
rect 6968 10272 6974 10324
rect 7026 10272 7032 10324
rect 6360 10064 6936 10092
rect 5406 9946 6304 9984
rect 6908 9998 6936 10064
rect 7079 9998 7085 10010
rect 6908 9970 7085 9998
rect 7079 9958 7085 9970
rect 7137 9958 7143 10010
rect 5406 9945 5603 9946
rect 5406 9939 5412 9945
rect 3475 9862 5063 9904
rect 5029 9784 5081 9790
rect 3472 9737 4907 9776
rect 1348 9603 1880 9646
rect 1348 9594 1398 9603
rect 1450 9594 1462 9603
rect 1348 9560 1383 9594
rect 1450 9560 1455 9594
rect 1348 9551 1398 9560
rect 1450 9551 1462 9560
rect 1514 9551 1526 9603
rect 1578 9551 1590 9603
rect 1642 9551 1654 9603
rect 1706 9551 1718 9603
rect 1770 9594 1782 9603
rect 1834 9594 1880 9603
rect 1777 9560 1782 9594
rect 1849 9560 1880 9594
rect 3472 9579 3511 9737
rect 4738 9695 4744 9702
rect 4558 9656 4744 9695
rect 1770 9551 1782 9560
rect 1834 9551 1880 9560
rect 550 9532 622 9536
rect 550 9480 560 9532
rect 612 9480 622 9532
rect 696 9530 768 9536
rect 550 9468 566 9480
rect 607 9468 622 9480
rect 682 9528 768 9530
rect 682 9476 702 9528
rect 754 9476 768 9528
rect 682 9474 710 9476
rect 550 9438 622 9468
rect 696 9468 710 9474
rect 751 9468 768 9476
rect 696 9438 768 9468
rect 840 9513 912 9542
rect 840 9473 856 9513
rect 897 9473 912 9513
rect 840 9444 912 9473
rect 994 9513 1066 9542
rect 994 9473 1009 9513
rect 1050 9473 1066 9513
rect 1348 9506 1880 9551
rect 994 9444 1066 9473
rect 564 9398 608 9438
rect 856 9378 900 9444
rect 378 9370 433 9376
rect 846 9326 852 9378
rect 904 9326 910 9378
rect 378 9085 433 9315
rect 856 9286 900 9326
rect 1008 9286 1052 9444
rect 1407 9440 1448 9506
rect 1693 9440 1735 9506
rect 1941 9503 2687 9548
rect 1404 9393 1450 9440
rect 1404 9359 1410 9393
rect 1444 9359 1450 9393
rect 1404 9321 1450 9359
rect 1404 9287 1410 9321
rect 1444 9287 1450 9321
rect 708 9242 900 9286
rect 372 9030 378 9085
rect 433 9030 439 9085
rect 708 9008 752 9242
rect 998 9234 1004 9286
rect 1056 9234 1062 9286
rect 1404 9240 1450 9287
rect 1562 9393 1608 9440
rect 1562 9359 1568 9393
rect 1602 9359 1608 9393
rect 1562 9321 1608 9359
rect 1562 9287 1568 9321
rect 1602 9287 1608 9321
rect 1562 9240 1608 9287
rect 1692 9393 1738 9440
rect 1692 9359 1698 9393
rect 1732 9359 1738 9393
rect 1692 9321 1738 9359
rect 1692 9287 1698 9321
rect 1732 9287 1738 9321
rect 1692 9240 1738 9287
rect 1850 9437 1896 9440
rect 1941 9437 1986 9503
rect 1850 9393 1986 9437
rect 1850 9359 1856 9393
rect 1890 9392 1986 9393
rect 2024 9393 2070 9440
rect 1890 9359 1896 9392
rect 1850 9321 1896 9359
rect 2024 9359 2030 9393
rect 2064 9359 2070 9393
rect 2024 9324 2070 9359
rect 1998 9322 2070 9324
rect 1850 9287 1856 9321
rect 1890 9287 1896 9321
rect 1850 9240 1896 9287
rect 1928 9321 2070 9322
rect 1928 9297 2030 9321
rect 1928 9280 1935 9297
rect 1929 9245 1935 9280
rect 1987 9287 2030 9297
rect 2064 9287 2070 9321
rect 1987 9280 2070 9287
rect 1987 9245 1993 9280
rect 2024 9240 2070 9280
rect 2182 9396 2228 9440
rect 2366 9396 2412 9440
rect 2182 9393 2412 9396
rect 2182 9359 2188 9393
rect 2222 9359 2372 9393
rect 2406 9359 2412 9393
rect 2182 9321 2412 9359
rect 2182 9287 2188 9321
rect 2222 9287 2372 9321
rect 2406 9287 2412 9321
rect 2182 9270 2412 9287
rect 2182 9240 2228 9270
rect 2366 9240 2412 9270
rect 2524 9393 2570 9440
rect 2524 9359 2530 9393
rect 2564 9359 2570 9393
rect 2642 9369 2687 9503
rect 3118 9540 3511 9579
rect 3724 9602 4264 9646
rect 3724 9550 3776 9602
rect 3828 9593 3840 9602
rect 3892 9593 3904 9602
rect 3956 9593 3968 9602
rect 4020 9593 4032 9602
rect 4084 9593 4096 9602
rect 4148 9593 4160 9602
rect 3831 9559 3840 9593
rect 3903 9559 3904 9593
rect 4084 9559 4085 9593
rect 4148 9559 4157 9593
rect 3828 9550 3840 9559
rect 3892 9550 3904 9559
rect 3956 9550 3968 9559
rect 4020 9550 4032 9559
rect 4084 9550 4096 9559
rect 4148 9550 4160 9559
rect 4212 9550 4264 9602
rect 2774 9496 2816 9497
rect 2758 9488 2816 9496
rect 2758 9436 2769 9488
rect 2821 9436 2827 9488
rect 3118 9440 3157 9540
rect 3724 9506 4264 9550
rect 3741 9450 3787 9506
rect 3736 9449 3787 9450
rect 2758 9393 2816 9436
rect 2524 9321 2570 9359
rect 2524 9287 2530 9321
rect 2564 9287 2570 9321
rect 2524 9280 2570 9287
rect 2613 9341 2715 9369
rect 2613 9307 2647 9341
rect 2681 9307 2715 9341
rect 2524 9240 2574 9280
rect 2613 9279 2715 9307
rect 2758 9359 2776 9393
rect 2810 9359 2816 9393
rect 2758 9321 2816 9359
rect 2758 9287 2776 9321
rect 2810 9287 2816 9321
rect 1008 9180 1052 9234
rect 1245 9199 1328 9218
rect 852 9136 1052 9180
rect 1148 9197 1328 9199
rect 1148 9145 1155 9197
rect 1207 9187 1328 9197
rect 1207 9153 1269 9187
rect 1303 9153 1328 9187
rect 1207 9145 1328 9153
rect 1148 9144 1328 9145
rect 852 9014 896 9136
rect 1245 9123 1328 9144
rect 1568 9206 1602 9240
rect 1568 9196 1820 9206
rect 1568 9144 1758 9196
rect 1810 9144 1820 9196
rect 1568 9134 1820 9144
rect 1568 9102 1608 9134
rect 1853 9102 1892 9240
rect 2185 9102 2224 9240
rect 2255 9203 2325 9209
rect 2255 9194 2331 9203
rect 2255 9142 2270 9194
rect 2322 9142 2331 9194
rect 2255 9133 2331 9142
rect 2255 9127 2325 9133
rect 2368 9102 2407 9240
rect 2530 9206 2574 9240
rect 2758 9240 2816 9287
rect 2928 9393 2974 9440
rect 2928 9359 2934 9393
rect 2968 9380 2974 9393
rect 3114 9393 3160 9440
rect 3114 9380 3120 9393
rect 2968 9359 3120 9380
rect 3154 9359 3160 9393
rect 3272 9393 3318 9440
rect 3272 9383 3278 9393
rect 3312 9383 3318 9393
rect 3736 9403 3782 9449
rect 2928 9321 3160 9359
rect 3262 9331 3268 9383
rect 3320 9331 3326 9383
rect 3736 9369 3742 9403
rect 3776 9369 3782 9403
rect 3736 9331 3782 9369
rect 2928 9287 2934 9321
rect 2968 9287 3120 9321
rect 3154 9287 3160 9321
rect 2928 9270 3160 9287
rect 2928 9240 2974 9270
rect 3114 9240 3160 9270
rect 3272 9321 3318 9331
rect 3272 9287 3278 9321
rect 3312 9287 3318 9321
rect 3272 9240 3318 9287
rect 3736 9297 3742 9331
rect 3776 9297 3782 9331
rect 3736 9250 3782 9297
rect 3894 9403 3940 9450
rect 3894 9369 3900 9403
rect 3934 9369 3940 9403
rect 3894 9331 3940 9369
rect 3894 9297 3900 9331
rect 3934 9297 3940 9331
rect 3894 9250 3940 9297
rect 4044 9403 4090 9506
rect 4558 9450 4597 9656
rect 4738 9650 4744 9656
rect 4796 9650 4802 9702
rect 4868 9450 4907 9737
rect 5081 9743 7015 9773
rect 5029 9726 5081 9732
rect 6862 9695 6868 9702
rect 6516 9656 6868 9695
rect 5682 9602 6222 9646
rect 5682 9550 5734 9602
rect 5786 9592 5798 9602
rect 5850 9592 5862 9602
rect 5914 9592 5926 9602
rect 5978 9592 5990 9602
rect 6042 9592 6054 9602
rect 6106 9592 6118 9602
rect 5790 9558 5798 9592
rect 6042 9558 6044 9592
rect 6106 9558 6116 9592
rect 5786 9550 5798 9558
rect 5850 9550 5862 9558
rect 5914 9550 5926 9558
rect 5978 9550 5990 9558
rect 6042 9550 6054 9558
rect 6106 9550 6118 9558
rect 6170 9550 6222 9602
rect 5682 9506 6222 9550
rect 5700 9450 5746 9506
rect 4044 9369 4050 9403
rect 4084 9369 4090 9403
rect 4044 9331 4090 9369
rect 4044 9297 4050 9331
rect 4084 9297 4090 9331
rect 4044 9250 4090 9297
rect 4202 9403 4248 9450
rect 4202 9369 4208 9403
rect 4242 9369 4248 9403
rect 4396 9403 4442 9450
rect 4396 9377 4402 9403
rect 4202 9331 4248 9369
rect 4202 9297 4208 9331
rect 4242 9297 4248 9331
rect 4285 9375 4402 9377
rect 4285 9323 4292 9375
rect 4344 9369 4402 9375
rect 4436 9369 4442 9403
rect 4344 9331 4442 9369
rect 4344 9323 4402 9331
rect 4285 9322 4402 9323
rect 4202 9250 4248 9297
rect 4396 9297 4402 9322
rect 4436 9297 4442 9331
rect 4396 9250 4442 9297
rect 4554 9403 4600 9450
rect 4554 9369 4560 9403
rect 4594 9370 4600 9403
rect 4704 9403 4750 9450
rect 4704 9370 4710 9403
rect 4594 9369 4710 9370
rect 4744 9369 4750 9403
rect 4554 9331 4750 9369
rect 4554 9297 4560 9331
rect 4594 9304 4710 9331
rect 4594 9297 4600 9304
rect 4554 9250 4600 9297
rect 4704 9297 4710 9304
rect 4744 9297 4750 9331
rect 4704 9250 4750 9297
rect 4862 9403 4908 9450
rect 4862 9369 4868 9403
rect 4902 9369 4908 9403
rect 5694 9404 5740 9450
rect 5027 9374 5057 9383
rect 4862 9331 4908 9369
rect 4862 9297 4868 9331
rect 4902 9297 4908 9331
rect 5010 9322 5016 9374
rect 5068 9322 5074 9374
rect 5694 9370 5700 9404
rect 5734 9370 5740 9404
rect 5694 9332 5740 9370
rect 4862 9250 4908 9297
rect 5026 9281 5057 9322
rect 5694 9298 5700 9332
rect 5734 9298 5740 9332
rect 2758 9206 2802 9240
rect 2530 9162 2656 9206
rect 1242 9082 1248 9086
rect 1138 9038 1248 9082
rect 1138 9014 1182 9038
rect 1242 9034 1248 9038
rect 1300 9034 1306 9086
rect 1404 9069 1450 9102
rect 1404 9035 1410 9069
rect 1444 9035 1450 9069
rect 1404 9031 1450 9035
rect 378 8986 434 8992
rect 550 8986 622 9008
rect 434 8980 622 8986
rect 434 8940 565 8980
rect 606 8940 622 8980
rect 434 8930 622 8940
rect 378 8924 434 8930
rect 550 8910 622 8930
rect 696 8980 768 9008
rect 696 8940 712 8980
rect 753 8940 768 8980
rect 696 8910 768 8940
rect 840 8985 912 9014
rect 840 8945 856 8985
rect 897 8945 912 8985
rect 840 8916 912 8945
rect 994 8986 1182 9014
rect 994 8946 1010 8986
rect 1051 8970 1182 8986
rect 1399 9002 1450 9031
rect 1562 9069 1608 9102
rect 1562 9035 1568 9069
rect 1602 9035 1608 9069
rect 1692 9069 1738 9102
rect 1692 9040 1698 9069
rect 1562 9002 1608 9035
rect 1690 9035 1698 9040
rect 1732 9040 1738 9069
rect 1850 9069 1896 9102
rect 2024 9086 2070 9102
rect 1732 9035 1740 9040
rect 1051 8946 1066 8970
rect 1399 8956 1449 9002
rect 1690 8956 1740 9035
rect 1850 9035 1856 9069
rect 1890 9035 1896 9069
rect 1850 9002 1896 9035
rect 2014 9034 2020 9086
rect 2072 9034 2078 9086
rect 2182 9069 2228 9102
rect 2182 9035 2188 9069
rect 2222 9035 2228 9069
rect 2024 9002 2070 9034
rect 2182 9002 2228 9035
rect 2366 9069 2412 9102
rect 2524 9084 2570 9102
rect 2366 9035 2372 9069
rect 2406 9035 2412 9069
rect 2366 9002 2412 9035
rect 2516 9032 2522 9084
rect 2574 9032 2580 9084
rect 2524 9002 2570 9032
rect 2024 8970 2068 9002
rect 2612 8970 2656 9162
rect 994 8916 1066 8946
rect 1324 8901 1960 8956
rect 2024 8926 2656 8970
rect 2694 9162 2802 9206
rect 2832 9192 2904 9202
rect 2694 8964 2738 9162
rect 2832 9140 2842 9192
rect 2894 9140 2904 9192
rect 2832 9130 2904 9140
rect 2933 9102 2972 9240
rect 3118 9102 3157 9240
rect 3272 9196 3316 9240
rect 3268 9190 3320 9196
rect 3555 9165 3561 9217
rect 3613 9210 3619 9217
rect 3662 9210 3713 9222
rect 3613 9207 3713 9210
rect 3613 9173 3670 9207
rect 3704 9173 3713 9207
rect 3613 9171 3713 9173
rect 3613 9165 3619 9171
rect 3662 9159 3713 9171
rect 3897 9201 3936 9250
rect 3976 9208 4027 9213
rect 3970 9201 3976 9208
rect 3897 9162 3976 9201
rect 3268 9132 3320 9138
rect 3897 9112 3936 9162
rect 3970 9156 3976 9162
rect 4028 9156 4034 9208
rect 4206 9194 4245 9250
rect 4300 9194 4347 9205
rect 4206 9192 4347 9194
rect 4206 9159 4306 9192
rect 3976 9150 4027 9156
rect 4206 9112 4245 9159
rect 4300 9158 4306 9159
rect 4340 9158 4347 9192
rect 4300 9146 4347 9158
rect 2766 9096 2818 9102
rect 2766 9038 2776 9044
rect 2770 9035 2776 9038
rect 2810 9038 2818 9044
rect 2928 9069 2974 9102
rect 2810 9035 2816 9038
rect 2770 9002 2816 9035
rect 2928 9035 2934 9069
rect 2968 9035 2974 9069
rect 2928 9002 2974 9035
rect 3114 9069 3160 9102
rect 3114 9035 3120 9069
rect 3154 9035 3160 9069
rect 3114 9002 3160 9035
rect 3272 9069 3318 9102
rect 3272 9035 3278 9069
rect 3312 9035 3318 9069
rect 3272 9002 3318 9035
rect 3274 8964 3318 9002
rect 2694 8920 3318 8964
rect 3736 9079 3782 9112
rect 3736 9045 3742 9079
rect 3776 9045 3782 9079
rect 3736 9012 3782 9045
rect 3894 9079 3940 9112
rect 3894 9045 3900 9079
rect 3934 9045 3940 9079
rect 4044 9079 4090 9112
rect 4044 9050 4050 9079
rect 3894 9012 3940 9045
rect 4042 9045 4050 9050
rect 4084 9045 4090 9079
rect 4042 9012 4090 9045
rect 4202 9079 4248 9112
rect 4202 9045 4208 9079
rect 4242 9045 4248 9079
rect 4202 9012 4248 9045
rect 3736 8956 3780 9012
rect 4042 8956 4089 9012
rect 1324 8849 1360 8901
rect 1412 8849 1424 8901
rect 1476 8892 1488 8901
rect 1540 8892 1552 8901
rect 1604 8892 1616 8901
rect 1668 8892 1680 8901
rect 1732 8892 1744 8901
rect 1796 8892 1808 8901
rect 1479 8858 1488 8892
rect 1551 8858 1552 8892
rect 1732 8858 1733 8892
rect 1796 8858 1805 8892
rect 1476 8849 1488 8858
rect 1540 8849 1552 8858
rect 1604 8849 1616 8858
rect 1668 8849 1680 8858
rect 1732 8849 1744 8858
rect 1796 8849 1808 8858
rect 1860 8849 1872 8901
rect 1924 8849 1960 8901
rect 3704 8912 4244 8956
rect 3704 8903 3756 8912
rect 3808 8903 3820 8912
rect 1324 8816 1960 8849
rect 2346 8871 2426 8896
rect 2346 8867 3517 8871
rect 2346 8833 2369 8867
rect 2403 8833 3517 8867
rect 2346 8829 3517 8833
rect 2346 8804 2426 8829
rect 2636 8771 2702 8783
rect 272 8717 278 8771
rect 332 8717 2642 8771
rect 2696 8717 2702 8771
rect 2636 8705 2702 8717
rect 3475 8676 3517 8829
rect 3704 8869 3741 8903
rect 3808 8869 3813 8903
rect 3704 8860 3756 8869
rect 3808 8860 3820 8869
rect 3872 8860 3884 8912
rect 3936 8860 3948 8912
rect 4000 8860 4012 8912
rect 4064 8860 4076 8912
rect 4128 8903 4140 8912
rect 4192 8903 4244 8912
rect 4135 8869 4140 8903
rect 4207 8869 4244 8903
rect 4128 8860 4140 8869
rect 4192 8860 4244 8869
rect 3704 8816 4244 8860
rect 3559 8711 3565 8763
rect 3617 8756 3623 8763
rect 4306 8756 4345 9146
rect 4558 9114 4597 9250
rect 4628 9219 4680 9225
rect 4625 9170 4628 9216
rect 4680 9170 4683 9216
rect 4875 9174 4904 9250
rect 4628 9161 4680 9167
rect 4875 9146 4980 9174
rect 4396 9081 4442 9114
rect 4396 9047 4402 9081
rect 4436 9047 4442 9081
rect 4396 9014 4442 9047
rect 4554 9094 4600 9114
rect 4704 9094 4750 9114
rect 4862 9094 4908 9114
rect 4554 9081 4750 9094
rect 4554 9047 4560 9081
rect 4594 9047 4710 9081
rect 4744 9047 4750 9081
rect 4554 9028 4750 9047
rect 4856 9042 4862 9094
rect 4914 9042 4920 9094
rect 4554 9014 4600 9028
rect 4704 9014 4750 9028
rect 4862 9014 4908 9042
rect 4402 8864 4430 9014
rect 4558 8969 4597 9014
rect 4552 8963 4604 8969
rect 4552 8905 4604 8911
rect 4952 8864 4980 9146
rect 5026 9096 5056 9281
rect 5694 9250 5740 9298
rect 5852 9404 5898 9450
rect 5852 9370 5858 9404
rect 5892 9370 5898 9404
rect 5852 9332 5898 9370
rect 5852 9298 5858 9332
rect 5892 9298 5898 9332
rect 5852 9250 5898 9298
rect 6002 9404 6048 9506
rect 6516 9450 6556 9656
rect 6862 9650 6868 9656
rect 6920 9650 6926 9702
rect 6985 9690 7015 9743
rect 6985 9661 7016 9690
rect 6002 9370 6008 9404
rect 6042 9370 6048 9404
rect 6002 9332 6048 9370
rect 6002 9298 6008 9332
rect 6042 9298 6048 9332
rect 6002 9250 6048 9298
rect 6160 9404 6206 9450
rect 6160 9370 6166 9404
rect 6200 9370 6206 9404
rect 6354 9404 6400 9450
rect 6354 9378 6360 9404
rect 6160 9332 6206 9370
rect 6160 9298 6166 9332
rect 6200 9298 6206 9332
rect 6244 9376 6360 9378
rect 6244 9324 6250 9376
rect 6302 9370 6360 9376
rect 6394 9370 6400 9404
rect 6302 9332 6400 9370
rect 6302 9324 6360 9332
rect 6244 9322 6360 9324
rect 6160 9250 6206 9298
rect 6354 9298 6360 9322
rect 6394 9298 6400 9332
rect 6354 9250 6400 9298
rect 6512 9404 6558 9450
rect 6512 9370 6518 9404
rect 6552 9370 6558 9404
rect 6662 9404 6708 9450
rect 6662 9370 6668 9404
rect 6702 9370 6708 9404
rect 6512 9332 6708 9370
rect 6512 9298 6518 9332
rect 6552 9304 6668 9332
rect 6552 9298 6558 9304
rect 6512 9250 6558 9298
rect 6662 9298 6668 9304
rect 6702 9298 6708 9332
rect 6662 9250 6708 9298
rect 6820 9404 6866 9450
rect 6820 9370 6826 9404
rect 6860 9370 6866 9404
rect 6986 9374 7016 9661
rect 6820 9332 6866 9370
rect 6820 9298 6826 9332
rect 6860 9298 6866 9332
rect 6968 9322 6974 9374
rect 7026 9322 7032 9374
rect 6820 9250 6866 9298
rect 6984 9282 7016 9322
rect 5111 9165 5117 9217
rect 5169 9210 5175 9217
rect 5620 9210 5672 9222
rect 5169 9208 5672 9210
rect 5169 9174 5628 9208
rect 5662 9174 5672 9208
rect 5169 9171 5672 9174
rect 5169 9165 5175 9171
rect 5620 9160 5672 9171
rect 5856 9202 5894 9250
rect 5934 9208 5986 9214
rect 5928 9202 5934 9208
rect 5856 9162 5934 9202
rect 5856 9112 5894 9162
rect 5928 9156 5934 9162
rect 5986 9156 5992 9208
rect 6164 9194 6204 9250
rect 6258 9194 6306 9206
rect 6164 9192 6306 9194
rect 6164 9160 6264 9192
rect 5934 9150 5986 9156
rect 6164 9112 6204 9160
rect 6258 9158 6264 9160
rect 6298 9158 6306 9192
rect 6258 9146 6306 9158
rect 5009 9044 5015 9096
rect 5067 9044 5073 9096
rect 5694 9080 5740 9112
rect 5694 9046 5700 9080
rect 5734 9046 5740 9080
rect 4402 8836 4980 8864
rect 3617 8717 4345 8756
rect 3617 8711 3623 8717
rect 5021 8676 5063 9044
rect 5694 9012 5740 9046
rect 5852 9080 5898 9112
rect 5852 9046 5858 9080
rect 5892 9046 5898 9080
rect 6002 9080 6048 9112
rect 6002 9050 6008 9080
rect 5852 9012 5898 9046
rect 6000 9046 6008 9050
rect 6042 9046 6048 9080
rect 5694 8956 5738 9012
rect 6000 8956 6048 9046
rect 6160 9080 6206 9112
rect 6160 9046 6166 9080
rect 6200 9046 6206 9080
rect 6160 9012 6206 9046
rect 5662 8912 6202 8956
rect 5662 8904 5714 8912
rect 5766 8904 5778 8912
rect 5662 8870 5700 8904
rect 5766 8870 5772 8904
rect 5662 8860 5714 8870
rect 5766 8860 5778 8870
rect 5830 8860 5842 8912
rect 5894 8860 5906 8912
rect 5958 8860 5970 8912
rect 6022 8860 6034 8912
rect 6086 8904 6098 8912
rect 6150 8904 6202 8912
rect 6094 8870 6098 8904
rect 6166 8870 6202 8904
rect 6086 8860 6098 8870
rect 6150 8860 6202 8870
rect 5662 8816 6202 8860
rect 5111 8711 5117 8763
rect 5169 8756 5175 8763
rect 6264 8756 6304 9146
rect 6516 9114 6556 9250
rect 6586 9220 6638 9226
rect 6584 9170 6586 9216
rect 6638 9170 6642 9216
rect 6834 9174 6862 9250
rect 6586 9162 6638 9168
rect 6834 9146 6936 9174
rect 6354 9082 6400 9114
rect 6354 9048 6360 9082
rect 6394 9048 6400 9082
rect 6354 9014 6400 9048
rect 6512 9094 6558 9114
rect 6662 9094 6708 9114
rect 6820 9094 6866 9114
rect 6512 9082 6708 9094
rect 6512 9048 6518 9082
rect 6552 9048 6668 9082
rect 6702 9048 6708 9082
rect 6512 9028 6708 9048
rect 6814 9042 6820 9094
rect 6872 9042 6878 9094
rect 6512 9014 6558 9028
rect 6662 9014 6708 9028
rect 6820 9014 6866 9042
rect 6360 8864 6388 9014
rect 6516 8970 6556 9014
rect 6510 8964 6562 8970
rect 6510 8906 6562 8912
rect 6908 8864 6936 9146
rect 6984 9096 7014 9282
rect 6968 9044 6974 9096
rect 7026 9044 7032 9096
rect 6360 8836 6936 8864
rect 6908 8772 6936 8836
rect 5169 8718 6304 8756
rect 6346 8744 6936 8772
rect 5169 8717 5572 8718
rect 5169 8711 5175 8717
rect 3475 8634 5063 8676
rect 5035 8593 5087 8599
rect 3472 8509 4907 8548
rect 6346 8581 6374 8744
rect 6908 8742 6936 8744
rect 6512 8678 6564 8684
rect 6512 8620 6564 8626
rect 5087 8553 6374 8581
rect 6523 8563 6553 8620
rect 5035 8535 5087 8541
rect 6523 8533 7015 8563
rect 1348 8375 1880 8418
rect 1348 8366 1398 8375
rect 1450 8366 1462 8375
rect 1348 8332 1383 8366
rect 1450 8332 1455 8366
rect 1348 8323 1398 8332
rect 1450 8323 1462 8332
rect 1514 8323 1526 8375
rect 1578 8323 1590 8375
rect 1642 8323 1654 8375
rect 1706 8323 1718 8375
rect 1770 8366 1782 8375
rect 1834 8366 1880 8375
rect 1777 8332 1782 8366
rect 1849 8332 1880 8366
rect 3472 8351 3511 8509
rect 4738 8467 4744 8474
rect 4558 8428 4744 8467
rect 1770 8323 1782 8332
rect 1834 8323 1880 8332
rect 550 8304 622 8308
rect 550 8252 560 8304
rect 612 8252 622 8304
rect 696 8302 768 8308
rect 550 8240 566 8252
rect 607 8240 622 8252
rect 682 8300 768 8302
rect 682 8248 702 8300
rect 754 8248 768 8300
rect 682 8246 710 8248
rect 550 8210 622 8240
rect 696 8240 710 8246
rect 751 8240 768 8248
rect 696 8210 768 8240
rect 840 8285 912 8314
rect 840 8245 856 8285
rect 897 8245 912 8285
rect 840 8216 912 8245
rect 994 8285 1066 8314
rect 994 8245 1009 8285
rect 1050 8245 1066 8285
rect 1348 8278 1880 8323
rect 994 8216 1066 8245
rect 564 8170 608 8210
rect 856 8150 900 8216
rect 378 8142 433 8148
rect 846 8098 852 8150
rect 904 8098 910 8150
rect 378 7857 433 8087
rect 856 8058 900 8098
rect 1008 8058 1052 8216
rect 1407 8212 1448 8278
rect 1693 8212 1735 8278
rect 1941 8275 2687 8320
rect 1404 8165 1450 8212
rect 1404 8131 1410 8165
rect 1444 8131 1450 8165
rect 1404 8093 1450 8131
rect 1404 8059 1410 8093
rect 1444 8059 1450 8093
rect 708 8014 900 8058
rect 372 7802 378 7857
rect 433 7802 439 7857
rect 708 7780 752 8014
rect 998 8006 1004 8058
rect 1056 8006 1062 8058
rect 1404 8012 1450 8059
rect 1562 8165 1608 8212
rect 1562 8131 1568 8165
rect 1602 8131 1608 8165
rect 1562 8093 1608 8131
rect 1562 8059 1568 8093
rect 1602 8059 1608 8093
rect 1562 8012 1608 8059
rect 1692 8165 1738 8212
rect 1692 8131 1698 8165
rect 1732 8131 1738 8165
rect 1692 8093 1738 8131
rect 1692 8059 1698 8093
rect 1732 8059 1738 8093
rect 1692 8012 1738 8059
rect 1850 8209 1896 8212
rect 1941 8209 1986 8275
rect 1850 8165 1986 8209
rect 1850 8131 1856 8165
rect 1890 8164 1986 8165
rect 2024 8165 2070 8212
rect 1890 8131 1896 8164
rect 1850 8093 1896 8131
rect 2024 8131 2030 8165
rect 2064 8131 2070 8165
rect 2024 8096 2070 8131
rect 1998 8094 2070 8096
rect 1850 8059 1856 8093
rect 1890 8059 1896 8093
rect 1850 8012 1896 8059
rect 1928 8093 2070 8094
rect 1928 8069 2030 8093
rect 1928 8052 1935 8069
rect 1929 8017 1935 8052
rect 1987 8059 2030 8069
rect 2064 8059 2070 8093
rect 1987 8052 2070 8059
rect 1987 8017 1993 8052
rect 2024 8012 2070 8052
rect 2182 8168 2228 8212
rect 2366 8168 2412 8212
rect 2182 8165 2412 8168
rect 2182 8131 2188 8165
rect 2222 8131 2372 8165
rect 2406 8131 2412 8165
rect 2182 8093 2412 8131
rect 2182 8059 2188 8093
rect 2222 8059 2372 8093
rect 2406 8059 2412 8093
rect 2182 8042 2412 8059
rect 2182 8012 2228 8042
rect 2366 8012 2412 8042
rect 2524 8165 2570 8212
rect 2524 8131 2530 8165
rect 2564 8131 2570 8165
rect 2642 8141 2687 8275
rect 3118 8312 3511 8351
rect 3724 8374 4264 8418
rect 3724 8322 3776 8374
rect 3828 8365 3840 8374
rect 3892 8365 3904 8374
rect 3956 8365 3968 8374
rect 4020 8365 4032 8374
rect 4084 8365 4096 8374
rect 4148 8365 4160 8374
rect 3831 8331 3840 8365
rect 3903 8331 3904 8365
rect 4084 8331 4085 8365
rect 4148 8331 4157 8365
rect 3828 8322 3840 8331
rect 3892 8322 3904 8331
rect 3956 8322 3968 8331
rect 4020 8322 4032 8331
rect 4084 8322 4096 8331
rect 4148 8322 4160 8331
rect 4212 8322 4264 8374
rect 2774 8268 2816 8269
rect 2758 8260 2816 8268
rect 2758 8208 2769 8260
rect 2821 8208 2827 8260
rect 3118 8212 3157 8312
rect 3724 8278 4264 8322
rect 3741 8222 3787 8278
rect 3736 8221 3787 8222
rect 2758 8165 2816 8208
rect 2524 8093 2570 8131
rect 2524 8059 2530 8093
rect 2564 8059 2570 8093
rect 2524 8052 2570 8059
rect 2613 8113 2715 8141
rect 2613 8079 2647 8113
rect 2681 8079 2715 8113
rect 2524 8012 2574 8052
rect 2613 8051 2715 8079
rect 2758 8131 2776 8165
rect 2810 8131 2816 8165
rect 2758 8093 2816 8131
rect 2758 8059 2776 8093
rect 2810 8059 2816 8093
rect 1008 7952 1052 8006
rect 1245 7971 1328 7990
rect 852 7908 1052 7952
rect 1148 7969 1328 7971
rect 1148 7917 1155 7969
rect 1207 7959 1328 7969
rect 1207 7925 1269 7959
rect 1303 7925 1328 7959
rect 1207 7917 1328 7925
rect 1148 7916 1328 7917
rect 852 7786 896 7908
rect 1245 7895 1328 7916
rect 1568 7978 1602 8012
rect 1568 7968 1820 7978
rect 1568 7916 1758 7968
rect 1810 7916 1820 7968
rect 1568 7906 1820 7916
rect 1568 7874 1608 7906
rect 1853 7874 1892 8012
rect 2185 7874 2224 8012
rect 2255 7975 2325 7981
rect 2255 7966 2331 7975
rect 2255 7914 2270 7966
rect 2322 7914 2331 7966
rect 2255 7905 2331 7914
rect 2255 7899 2325 7905
rect 2368 7874 2407 8012
rect 2530 7978 2574 8012
rect 2758 8012 2816 8059
rect 2928 8165 2974 8212
rect 2928 8131 2934 8165
rect 2968 8152 2974 8165
rect 3114 8165 3160 8212
rect 3114 8152 3120 8165
rect 2968 8131 3120 8152
rect 3154 8131 3160 8165
rect 3272 8165 3318 8212
rect 3272 8155 3278 8165
rect 3312 8155 3318 8165
rect 3736 8175 3782 8221
rect 2928 8093 3160 8131
rect 3262 8103 3268 8155
rect 3320 8103 3326 8155
rect 3736 8141 3742 8175
rect 3776 8141 3782 8175
rect 3736 8103 3782 8141
rect 2928 8059 2934 8093
rect 2968 8059 3120 8093
rect 3154 8059 3160 8093
rect 2928 8042 3160 8059
rect 2928 8012 2974 8042
rect 3114 8012 3160 8042
rect 3272 8093 3318 8103
rect 3272 8059 3278 8093
rect 3312 8059 3318 8093
rect 3272 8012 3318 8059
rect 3736 8069 3742 8103
rect 3776 8069 3782 8103
rect 3736 8022 3782 8069
rect 3894 8175 3940 8222
rect 3894 8141 3900 8175
rect 3934 8141 3940 8175
rect 3894 8103 3940 8141
rect 3894 8069 3900 8103
rect 3934 8069 3940 8103
rect 3894 8022 3940 8069
rect 4044 8175 4090 8278
rect 4558 8222 4597 8428
rect 4738 8422 4744 8428
rect 4796 8422 4802 8474
rect 4868 8222 4907 8509
rect 6837 8467 6843 8474
rect 6516 8428 6843 8467
rect 5682 8374 6222 8418
rect 5682 8322 5734 8374
rect 5786 8364 5798 8374
rect 5850 8364 5862 8374
rect 5914 8364 5926 8374
rect 5978 8364 5990 8374
rect 6042 8364 6054 8374
rect 6106 8364 6118 8374
rect 5790 8330 5798 8364
rect 6042 8330 6044 8364
rect 6106 8330 6116 8364
rect 5786 8322 5798 8330
rect 5850 8322 5862 8330
rect 5914 8322 5926 8330
rect 5978 8322 5990 8330
rect 6042 8322 6054 8330
rect 6106 8322 6118 8330
rect 6170 8322 6222 8374
rect 5682 8278 6222 8322
rect 5700 8222 5746 8278
rect 4044 8141 4050 8175
rect 4084 8141 4090 8175
rect 4044 8103 4090 8141
rect 4044 8069 4050 8103
rect 4084 8069 4090 8103
rect 4044 8022 4090 8069
rect 4202 8175 4248 8222
rect 4202 8141 4208 8175
rect 4242 8141 4248 8175
rect 4396 8175 4442 8222
rect 4396 8149 4402 8175
rect 4202 8103 4248 8141
rect 4202 8069 4208 8103
rect 4242 8069 4248 8103
rect 4285 8147 4402 8149
rect 4285 8095 4292 8147
rect 4344 8141 4402 8147
rect 4436 8141 4442 8175
rect 4344 8103 4442 8141
rect 4344 8095 4402 8103
rect 4285 8094 4402 8095
rect 4202 8022 4248 8069
rect 4396 8069 4402 8094
rect 4436 8069 4442 8103
rect 4396 8022 4442 8069
rect 4554 8175 4600 8222
rect 4554 8141 4560 8175
rect 4594 8142 4600 8175
rect 4704 8175 4750 8222
rect 4704 8142 4710 8175
rect 4594 8141 4710 8142
rect 4744 8141 4750 8175
rect 4554 8103 4750 8141
rect 4554 8069 4560 8103
rect 4594 8076 4710 8103
rect 4594 8069 4600 8076
rect 4554 8022 4600 8069
rect 4704 8069 4710 8076
rect 4744 8069 4750 8103
rect 4704 8022 4750 8069
rect 4862 8175 4908 8222
rect 4862 8141 4868 8175
rect 4902 8141 4908 8175
rect 5694 8176 5740 8222
rect 5027 8146 5057 8155
rect 4862 8103 4908 8141
rect 4862 8069 4868 8103
rect 4902 8069 4908 8103
rect 5010 8094 5016 8146
rect 5068 8094 5074 8146
rect 5694 8142 5700 8176
rect 5734 8142 5740 8176
rect 5694 8104 5740 8142
rect 4862 8022 4908 8069
rect 5026 8053 5057 8094
rect 5694 8070 5700 8104
rect 5734 8070 5740 8104
rect 2758 7978 2802 8012
rect 2530 7934 2656 7978
rect 1242 7854 1248 7858
rect 1138 7810 1248 7854
rect 1138 7786 1182 7810
rect 1242 7806 1248 7810
rect 1300 7806 1306 7858
rect 1404 7841 1450 7874
rect 1404 7807 1410 7841
rect 1444 7807 1450 7841
rect 1404 7803 1450 7807
rect 378 7758 434 7764
rect 550 7758 622 7780
rect 434 7752 622 7758
rect 434 7712 565 7752
rect 606 7712 622 7752
rect 434 7702 622 7712
rect 378 7696 434 7702
rect 550 7682 622 7702
rect 696 7752 768 7780
rect 696 7712 712 7752
rect 753 7712 768 7752
rect 696 7682 768 7712
rect 840 7757 912 7786
rect 840 7717 856 7757
rect 897 7717 912 7757
rect 840 7688 912 7717
rect 994 7758 1182 7786
rect 994 7718 1010 7758
rect 1051 7742 1182 7758
rect 1399 7774 1450 7803
rect 1562 7841 1608 7874
rect 1562 7807 1568 7841
rect 1602 7807 1608 7841
rect 1692 7841 1738 7874
rect 1692 7812 1698 7841
rect 1562 7774 1608 7807
rect 1690 7807 1698 7812
rect 1732 7812 1738 7841
rect 1850 7841 1896 7874
rect 2024 7858 2070 7874
rect 1732 7807 1740 7812
rect 1051 7718 1066 7742
rect 1399 7728 1449 7774
rect 1690 7728 1740 7807
rect 1850 7807 1856 7841
rect 1890 7807 1896 7841
rect 1850 7774 1896 7807
rect 2014 7806 2020 7858
rect 2072 7806 2078 7858
rect 2182 7841 2228 7874
rect 2182 7807 2188 7841
rect 2222 7807 2228 7841
rect 2024 7774 2070 7806
rect 2182 7774 2228 7807
rect 2366 7841 2412 7874
rect 2524 7856 2570 7874
rect 2366 7807 2372 7841
rect 2406 7807 2412 7841
rect 2366 7774 2412 7807
rect 2516 7804 2522 7856
rect 2574 7804 2580 7856
rect 2524 7774 2570 7804
rect 2024 7742 2068 7774
rect 2612 7742 2656 7934
rect 994 7688 1066 7718
rect 1324 7673 1960 7728
rect 2024 7698 2656 7742
rect 2694 7934 2802 7978
rect 2832 7964 2904 7974
rect 2694 7736 2738 7934
rect 2832 7912 2842 7964
rect 2894 7912 2904 7964
rect 2832 7902 2904 7912
rect 2933 7874 2972 8012
rect 3118 7874 3157 8012
rect 3272 7968 3316 8012
rect 3268 7962 3320 7968
rect 3555 7937 3561 7989
rect 3613 7982 3619 7989
rect 3662 7982 3713 7994
rect 3613 7979 3713 7982
rect 3613 7945 3670 7979
rect 3704 7945 3713 7979
rect 3613 7943 3713 7945
rect 3613 7937 3619 7943
rect 3662 7931 3713 7943
rect 3897 7973 3936 8022
rect 3976 7980 4027 7985
rect 3970 7973 3976 7980
rect 3897 7934 3976 7973
rect 3268 7904 3320 7910
rect 3897 7884 3936 7934
rect 3970 7928 3976 7934
rect 4028 7928 4034 7980
rect 4206 7966 4245 8022
rect 4300 7966 4347 7977
rect 4206 7964 4347 7966
rect 4206 7931 4306 7964
rect 3976 7922 4027 7928
rect 4206 7884 4245 7931
rect 4300 7930 4306 7931
rect 4340 7930 4347 7964
rect 4300 7918 4347 7930
rect 2766 7868 2818 7874
rect 2766 7810 2776 7816
rect 2770 7807 2776 7810
rect 2810 7810 2818 7816
rect 2928 7841 2974 7874
rect 2810 7807 2816 7810
rect 2770 7774 2816 7807
rect 2928 7807 2934 7841
rect 2968 7807 2974 7841
rect 2928 7774 2974 7807
rect 3114 7841 3160 7874
rect 3114 7807 3120 7841
rect 3154 7807 3160 7841
rect 3114 7774 3160 7807
rect 3272 7841 3318 7874
rect 3272 7807 3278 7841
rect 3312 7807 3318 7841
rect 3272 7774 3318 7807
rect 3274 7736 3318 7774
rect 2694 7692 3318 7736
rect 3736 7851 3782 7884
rect 3736 7817 3742 7851
rect 3776 7817 3782 7851
rect 3736 7784 3782 7817
rect 3894 7851 3940 7884
rect 3894 7817 3900 7851
rect 3934 7817 3940 7851
rect 4044 7851 4090 7884
rect 4044 7822 4050 7851
rect 3894 7784 3940 7817
rect 4042 7817 4050 7822
rect 4084 7817 4090 7851
rect 4042 7784 4090 7817
rect 4202 7851 4248 7884
rect 4202 7817 4208 7851
rect 4242 7817 4248 7851
rect 4202 7784 4248 7817
rect 3736 7728 3780 7784
rect 4042 7728 4089 7784
rect 1324 7621 1360 7673
rect 1412 7621 1424 7673
rect 1476 7664 1488 7673
rect 1540 7664 1552 7673
rect 1604 7664 1616 7673
rect 1668 7664 1680 7673
rect 1732 7664 1744 7673
rect 1796 7664 1808 7673
rect 1479 7630 1488 7664
rect 1551 7630 1552 7664
rect 1732 7630 1733 7664
rect 1796 7630 1805 7664
rect 1476 7621 1488 7630
rect 1540 7621 1552 7630
rect 1604 7621 1616 7630
rect 1668 7621 1680 7630
rect 1732 7621 1744 7630
rect 1796 7621 1808 7630
rect 1860 7621 1872 7673
rect 1924 7621 1960 7673
rect 3704 7684 4244 7728
rect 3704 7675 3756 7684
rect 3808 7675 3820 7684
rect 1324 7588 1960 7621
rect 2346 7643 2426 7668
rect 2346 7639 3517 7643
rect 2346 7605 2369 7639
rect 2403 7605 3517 7639
rect 2346 7601 3517 7605
rect 2346 7576 2426 7601
rect 2636 7543 2702 7555
rect 272 7489 278 7543
rect 332 7489 2642 7543
rect 2696 7489 2702 7543
rect 2636 7477 2702 7489
rect 3475 7448 3517 7601
rect 3704 7641 3741 7675
rect 3808 7641 3813 7675
rect 3704 7632 3756 7641
rect 3808 7632 3820 7641
rect 3872 7632 3884 7684
rect 3936 7632 3948 7684
rect 4000 7632 4012 7684
rect 4064 7632 4076 7684
rect 4128 7675 4140 7684
rect 4192 7675 4244 7684
rect 4135 7641 4140 7675
rect 4207 7641 4244 7675
rect 4128 7632 4140 7641
rect 4192 7632 4244 7641
rect 3704 7588 4244 7632
rect 3559 7483 3565 7535
rect 3617 7528 3623 7535
rect 4306 7528 4345 7918
rect 4558 7886 4597 8022
rect 4628 7991 4680 7997
rect 4625 7942 4628 7988
rect 4680 7942 4683 7988
rect 4875 7946 4904 8022
rect 4628 7933 4680 7939
rect 4875 7918 4980 7946
rect 4396 7853 4442 7886
rect 4396 7819 4402 7853
rect 4436 7819 4442 7853
rect 4396 7786 4442 7819
rect 4554 7866 4600 7886
rect 4704 7866 4750 7886
rect 4862 7866 4908 7886
rect 4554 7853 4750 7866
rect 4554 7819 4560 7853
rect 4594 7819 4710 7853
rect 4744 7819 4750 7853
rect 4554 7800 4750 7819
rect 4856 7814 4862 7866
rect 4914 7814 4920 7866
rect 4554 7786 4600 7800
rect 4704 7786 4750 7800
rect 4862 7786 4908 7814
rect 4402 7636 4430 7786
rect 4558 7741 4597 7786
rect 4552 7735 4604 7741
rect 4552 7677 4604 7683
rect 4952 7636 4980 7918
rect 5026 7868 5056 8053
rect 5694 8022 5740 8070
rect 5852 8176 5898 8222
rect 5852 8142 5858 8176
rect 5892 8142 5898 8176
rect 5852 8104 5898 8142
rect 5852 8070 5858 8104
rect 5892 8070 5898 8104
rect 5852 8022 5898 8070
rect 6002 8176 6048 8278
rect 6516 8222 6556 8428
rect 6837 8422 6843 8428
rect 6895 8422 6901 8474
rect 6985 8462 7015 8533
rect 6985 8433 7016 8462
rect 6002 8142 6008 8176
rect 6042 8142 6048 8176
rect 6002 8104 6048 8142
rect 6002 8070 6008 8104
rect 6042 8070 6048 8104
rect 6002 8022 6048 8070
rect 6160 8176 6206 8222
rect 6160 8142 6166 8176
rect 6200 8142 6206 8176
rect 6354 8176 6400 8222
rect 6354 8150 6360 8176
rect 6160 8104 6206 8142
rect 6160 8070 6166 8104
rect 6200 8070 6206 8104
rect 6244 8148 6360 8150
rect 6244 8096 6250 8148
rect 6302 8142 6360 8148
rect 6394 8142 6400 8176
rect 6302 8104 6400 8142
rect 6302 8096 6360 8104
rect 6244 8094 6360 8096
rect 6160 8022 6206 8070
rect 6354 8070 6360 8094
rect 6394 8070 6400 8104
rect 6354 8022 6400 8070
rect 6512 8176 6558 8222
rect 6512 8142 6518 8176
rect 6552 8142 6558 8176
rect 6662 8176 6708 8222
rect 6662 8142 6668 8176
rect 6702 8142 6708 8176
rect 6512 8104 6708 8142
rect 6512 8070 6518 8104
rect 6552 8076 6668 8104
rect 6552 8070 6558 8076
rect 6512 8022 6558 8070
rect 6662 8070 6668 8076
rect 6702 8070 6708 8104
rect 6662 8022 6708 8070
rect 6820 8176 6866 8222
rect 6820 8142 6826 8176
rect 6860 8142 6866 8176
rect 6986 8146 7016 8433
rect 6820 8104 6866 8142
rect 6820 8070 6826 8104
rect 6860 8070 6866 8104
rect 6968 8094 6974 8146
rect 7026 8094 7032 8146
rect 6820 8022 6866 8070
rect 6984 8054 7016 8094
rect 5191 7937 5197 7989
rect 5249 7982 5255 7989
rect 5620 7982 5672 7994
rect 5249 7980 5672 7982
rect 5249 7946 5628 7980
rect 5662 7946 5672 7980
rect 5249 7943 5672 7946
rect 5249 7937 5255 7943
rect 5620 7932 5672 7943
rect 5856 7974 5894 8022
rect 5934 7980 5986 7986
rect 5928 7974 5934 7980
rect 5856 7934 5934 7974
rect 5856 7884 5894 7934
rect 5928 7928 5934 7934
rect 5986 7928 5992 7980
rect 6164 7966 6204 8022
rect 6258 7966 6306 7978
rect 6164 7964 6306 7966
rect 6164 7932 6264 7964
rect 5934 7922 5986 7928
rect 6164 7884 6204 7932
rect 6258 7930 6264 7932
rect 6298 7930 6306 7964
rect 6258 7918 6306 7930
rect 5009 7816 5015 7868
rect 5067 7816 5073 7868
rect 5694 7852 5740 7884
rect 5694 7818 5700 7852
rect 5734 7818 5740 7852
rect 4402 7608 4980 7636
rect 3617 7489 4345 7528
rect 3617 7483 3623 7489
rect 5021 7448 5063 7816
rect 5694 7784 5740 7818
rect 5852 7852 5898 7884
rect 5852 7818 5858 7852
rect 5892 7818 5898 7852
rect 6002 7852 6048 7884
rect 6002 7822 6008 7852
rect 5852 7784 5898 7818
rect 6000 7818 6008 7822
rect 6042 7818 6048 7852
rect 5694 7728 5738 7784
rect 6000 7728 6048 7818
rect 6160 7852 6206 7884
rect 6160 7818 6166 7852
rect 6200 7818 6206 7852
rect 6160 7784 6206 7818
rect 5662 7684 6202 7728
rect 5662 7676 5714 7684
rect 5766 7676 5778 7684
rect 5662 7642 5700 7676
rect 5766 7642 5772 7676
rect 5662 7632 5714 7642
rect 5766 7632 5778 7642
rect 5830 7632 5842 7684
rect 5894 7632 5906 7684
rect 5958 7632 5970 7684
rect 6022 7632 6034 7684
rect 6086 7676 6098 7684
rect 6150 7676 6202 7684
rect 6094 7642 6098 7676
rect 6166 7642 6202 7676
rect 6086 7632 6098 7642
rect 6150 7632 6202 7642
rect 5662 7588 6202 7632
rect 5191 7483 5197 7535
rect 5249 7528 5255 7535
rect 6264 7528 6304 7918
rect 6516 7886 6556 8022
rect 6586 7992 6638 7998
rect 6584 7942 6586 7988
rect 6638 7942 6642 7988
rect 6834 7946 6862 8022
rect 6586 7934 6638 7940
rect 6834 7918 6936 7946
rect 6354 7854 6400 7886
rect 6354 7820 6360 7854
rect 6394 7820 6400 7854
rect 6354 7786 6400 7820
rect 6512 7866 6558 7886
rect 6662 7866 6708 7886
rect 6820 7866 6866 7886
rect 6512 7854 6708 7866
rect 6512 7820 6518 7854
rect 6552 7820 6668 7854
rect 6702 7820 6708 7854
rect 6512 7800 6708 7820
rect 6814 7814 6820 7866
rect 6872 7814 6878 7866
rect 6512 7786 6558 7800
rect 6662 7786 6708 7800
rect 6820 7786 6866 7814
rect 6360 7636 6388 7786
rect 6516 7742 6556 7786
rect 6510 7736 6562 7742
rect 6510 7678 6562 7684
rect 6908 7636 6936 7918
rect 6984 7868 7014 8054
rect 6968 7816 6974 7868
rect 7026 7816 7032 7868
rect 6360 7608 6936 7636
rect 5249 7490 6304 7528
rect 5249 7489 5587 7490
rect 5249 7483 5255 7489
rect 3475 7406 5063 7448
rect 6908 7436 6936 7608
rect 7107 7448 7159 7454
rect 6908 7408 7107 7436
rect 7107 7390 7159 7396
rect 5029 7328 5081 7334
rect 3472 7281 4907 7320
rect 1348 7147 1880 7190
rect 1348 7138 1398 7147
rect 1450 7138 1462 7147
rect 1348 7104 1383 7138
rect 1450 7104 1455 7138
rect 1348 7095 1398 7104
rect 1450 7095 1462 7104
rect 1514 7095 1526 7147
rect 1578 7095 1590 7147
rect 1642 7095 1654 7147
rect 1706 7095 1718 7147
rect 1770 7138 1782 7147
rect 1834 7138 1880 7147
rect 1777 7104 1782 7138
rect 1849 7104 1880 7138
rect 3472 7123 3511 7281
rect 4738 7239 4744 7246
rect 4558 7200 4744 7239
rect 1770 7095 1782 7104
rect 1834 7095 1880 7104
rect 550 7076 622 7080
rect 550 7024 560 7076
rect 612 7024 622 7076
rect 696 7074 768 7080
rect 550 7012 566 7024
rect 607 7012 622 7024
rect 682 7072 768 7074
rect 682 7020 702 7072
rect 754 7020 768 7072
rect 682 7018 710 7020
rect 550 6982 622 7012
rect 696 7012 710 7018
rect 751 7012 768 7020
rect 696 6982 768 7012
rect 840 7057 912 7086
rect 840 7017 856 7057
rect 897 7017 912 7057
rect 840 6988 912 7017
rect 994 7057 1066 7086
rect 994 7017 1009 7057
rect 1050 7017 1066 7057
rect 1348 7050 1880 7095
rect 994 6988 1066 7017
rect 564 6942 608 6982
rect 856 6922 900 6988
rect 378 6914 433 6920
rect 846 6870 852 6922
rect 904 6870 910 6922
rect 378 6629 433 6859
rect 856 6830 900 6870
rect 1008 6830 1052 6988
rect 1407 6984 1448 7050
rect 1693 6984 1735 7050
rect 1941 7047 2687 7092
rect 1404 6937 1450 6984
rect 1404 6903 1410 6937
rect 1444 6903 1450 6937
rect 1404 6865 1450 6903
rect 1404 6831 1410 6865
rect 1444 6831 1450 6865
rect 708 6786 900 6830
rect 372 6574 378 6629
rect 433 6574 439 6629
rect 708 6552 752 6786
rect 998 6778 1004 6830
rect 1056 6778 1062 6830
rect 1404 6784 1450 6831
rect 1562 6937 1608 6984
rect 1562 6903 1568 6937
rect 1602 6903 1608 6937
rect 1562 6865 1608 6903
rect 1562 6831 1568 6865
rect 1602 6831 1608 6865
rect 1562 6784 1608 6831
rect 1692 6937 1738 6984
rect 1692 6903 1698 6937
rect 1732 6903 1738 6937
rect 1692 6865 1738 6903
rect 1692 6831 1698 6865
rect 1732 6831 1738 6865
rect 1692 6784 1738 6831
rect 1850 6981 1896 6984
rect 1941 6981 1986 7047
rect 1850 6937 1986 6981
rect 1850 6903 1856 6937
rect 1890 6936 1986 6937
rect 2024 6937 2070 6984
rect 1890 6903 1896 6936
rect 1850 6865 1896 6903
rect 2024 6903 2030 6937
rect 2064 6903 2070 6937
rect 2024 6868 2070 6903
rect 1998 6866 2070 6868
rect 1850 6831 1856 6865
rect 1890 6831 1896 6865
rect 1850 6784 1896 6831
rect 1928 6865 2070 6866
rect 1928 6841 2030 6865
rect 1928 6824 1935 6841
rect 1929 6789 1935 6824
rect 1987 6831 2030 6841
rect 2064 6831 2070 6865
rect 1987 6824 2070 6831
rect 1987 6789 1993 6824
rect 2024 6784 2070 6824
rect 2182 6940 2228 6984
rect 2366 6940 2412 6984
rect 2182 6937 2412 6940
rect 2182 6903 2188 6937
rect 2222 6903 2372 6937
rect 2406 6903 2412 6937
rect 2182 6865 2412 6903
rect 2182 6831 2188 6865
rect 2222 6831 2372 6865
rect 2406 6831 2412 6865
rect 2182 6814 2412 6831
rect 2182 6784 2228 6814
rect 2366 6784 2412 6814
rect 2524 6937 2570 6984
rect 2524 6903 2530 6937
rect 2564 6903 2570 6937
rect 2642 6913 2687 7047
rect 3118 7084 3511 7123
rect 3724 7146 4264 7190
rect 3724 7094 3776 7146
rect 3828 7137 3840 7146
rect 3892 7137 3904 7146
rect 3956 7137 3968 7146
rect 4020 7137 4032 7146
rect 4084 7137 4096 7146
rect 4148 7137 4160 7146
rect 3831 7103 3840 7137
rect 3903 7103 3904 7137
rect 4084 7103 4085 7137
rect 4148 7103 4157 7137
rect 3828 7094 3840 7103
rect 3892 7094 3904 7103
rect 3956 7094 3968 7103
rect 4020 7094 4032 7103
rect 4084 7094 4096 7103
rect 4148 7094 4160 7103
rect 4212 7094 4264 7146
rect 2774 7040 2816 7041
rect 2758 7032 2816 7040
rect 2758 6980 2769 7032
rect 2821 6980 2827 7032
rect 3118 6984 3157 7084
rect 3724 7050 4264 7094
rect 3741 6994 3787 7050
rect 3736 6993 3787 6994
rect 2758 6937 2816 6980
rect 2524 6865 2570 6903
rect 2524 6831 2530 6865
rect 2564 6831 2570 6865
rect 2524 6824 2570 6831
rect 2613 6885 2715 6913
rect 2613 6851 2647 6885
rect 2681 6851 2715 6885
rect 2524 6784 2574 6824
rect 2613 6823 2715 6851
rect 2758 6903 2776 6937
rect 2810 6903 2816 6937
rect 2758 6865 2816 6903
rect 2758 6831 2776 6865
rect 2810 6831 2816 6865
rect 1008 6724 1052 6778
rect 1245 6743 1328 6762
rect 852 6680 1052 6724
rect 1148 6741 1328 6743
rect 1148 6689 1155 6741
rect 1207 6731 1328 6741
rect 1207 6697 1269 6731
rect 1303 6697 1328 6731
rect 1207 6689 1328 6697
rect 1148 6688 1328 6689
rect 852 6558 896 6680
rect 1245 6667 1328 6688
rect 1568 6750 1602 6784
rect 1568 6740 1820 6750
rect 1568 6688 1758 6740
rect 1810 6688 1820 6740
rect 1568 6678 1820 6688
rect 1568 6646 1608 6678
rect 1853 6646 1892 6784
rect 2185 6646 2224 6784
rect 2255 6747 2325 6753
rect 2255 6738 2331 6747
rect 2255 6686 2270 6738
rect 2322 6686 2331 6738
rect 2255 6677 2331 6686
rect 2255 6671 2325 6677
rect 2368 6646 2407 6784
rect 2530 6750 2574 6784
rect 2758 6784 2816 6831
rect 2928 6937 2974 6984
rect 2928 6903 2934 6937
rect 2968 6924 2974 6937
rect 3114 6937 3160 6984
rect 3114 6924 3120 6937
rect 2968 6903 3120 6924
rect 3154 6903 3160 6937
rect 3272 6937 3318 6984
rect 3272 6927 3278 6937
rect 3312 6927 3318 6937
rect 3736 6947 3782 6993
rect 2928 6865 3160 6903
rect 3262 6875 3268 6927
rect 3320 6875 3326 6927
rect 3736 6913 3742 6947
rect 3776 6913 3782 6947
rect 3736 6875 3782 6913
rect 2928 6831 2934 6865
rect 2968 6831 3120 6865
rect 3154 6831 3160 6865
rect 2928 6814 3160 6831
rect 2928 6784 2974 6814
rect 3114 6784 3160 6814
rect 3272 6865 3318 6875
rect 3272 6831 3278 6865
rect 3312 6831 3318 6865
rect 3272 6784 3318 6831
rect 3736 6841 3742 6875
rect 3776 6841 3782 6875
rect 3736 6794 3782 6841
rect 3894 6947 3940 6994
rect 3894 6913 3900 6947
rect 3934 6913 3940 6947
rect 3894 6875 3940 6913
rect 3894 6841 3900 6875
rect 3934 6841 3940 6875
rect 3894 6794 3940 6841
rect 4044 6947 4090 7050
rect 4558 6994 4597 7200
rect 4738 7194 4744 7200
rect 4796 7194 4802 7246
rect 4868 6994 4907 7281
rect 5081 7287 7015 7317
rect 5029 7270 5081 7276
rect 6862 7239 6868 7246
rect 6516 7200 6868 7239
rect 5682 7146 6222 7190
rect 5682 7094 5734 7146
rect 5786 7136 5798 7146
rect 5850 7136 5862 7146
rect 5914 7136 5926 7146
rect 5978 7136 5990 7146
rect 6042 7136 6054 7146
rect 6106 7136 6118 7146
rect 5790 7102 5798 7136
rect 6042 7102 6044 7136
rect 6106 7102 6116 7136
rect 5786 7094 5798 7102
rect 5850 7094 5862 7102
rect 5914 7094 5926 7102
rect 5978 7094 5990 7102
rect 6042 7094 6054 7102
rect 6106 7094 6118 7102
rect 6170 7094 6222 7146
rect 5682 7050 6222 7094
rect 5700 6994 5746 7050
rect 4044 6913 4050 6947
rect 4084 6913 4090 6947
rect 4044 6875 4090 6913
rect 4044 6841 4050 6875
rect 4084 6841 4090 6875
rect 4044 6794 4090 6841
rect 4202 6947 4248 6994
rect 4202 6913 4208 6947
rect 4242 6913 4248 6947
rect 4396 6947 4442 6994
rect 4396 6921 4402 6947
rect 4202 6875 4248 6913
rect 4202 6841 4208 6875
rect 4242 6841 4248 6875
rect 4285 6919 4402 6921
rect 4285 6867 4292 6919
rect 4344 6913 4402 6919
rect 4436 6913 4442 6947
rect 4344 6875 4442 6913
rect 4344 6867 4402 6875
rect 4285 6866 4402 6867
rect 4202 6794 4248 6841
rect 4396 6841 4402 6866
rect 4436 6841 4442 6875
rect 4396 6794 4442 6841
rect 4554 6947 4600 6994
rect 4554 6913 4560 6947
rect 4594 6914 4600 6947
rect 4704 6947 4750 6994
rect 4704 6914 4710 6947
rect 4594 6913 4710 6914
rect 4744 6913 4750 6947
rect 4554 6875 4750 6913
rect 4554 6841 4560 6875
rect 4594 6848 4710 6875
rect 4594 6841 4600 6848
rect 4554 6794 4600 6841
rect 4704 6841 4710 6848
rect 4744 6841 4750 6875
rect 4704 6794 4750 6841
rect 4862 6947 4908 6994
rect 4862 6913 4868 6947
rect 4902 6913 4908 6947
rect 5694 6948 5740 6994
rect 5027 6918 5057 6927
rect 4862 6875 4908 6913
rect 4862 6841 4868 6875
rect 4902 6841 4908 6875
rect 5010 6866 5016 6918
rect 5068 6866 5074 6918
rect 5694 6914 5700 6948
rect 5734 6914 5740 6948
rect 5694 6876 5740 6914
rect 4862 6794 4908 6841
rect 5026 6825 5057 6866
rect 5694 6842 5700 6876
rect 5734 6842 5740 6876
rect 2758 6750 2802 6784
rect 2530 6706 2656 6750
rect 1242 6626 1248 6630
rect 1138 6582 1248 6626
rect 1138 6558 1182 6582
rect 1242 6578 1248 6582
rect 1300 6578 1306 6630
rect 1404 6613 1450 6646
rect 1404 6579 1410 6613
rect 1444 6579 1450 6613
rect 1404 6575 1450 6579
rect 378 6530 434 6536
rect 550 6530 622 6552
rect 434 6524 622 6530
rect 434 6484 565 6524
rect 606 6484 622 6524
rect 434 6474 622 6484
rect 378 6468 434 6474
rect 550 6454 622 6474
rect 696 6524 768 6552
rect 696 6484 712 6524
rect 753 6484 768 6524
rect 696 6454 768 6484
rect 840 6529 912 6558
rect 840 6489 856 6529
rect 897 6489 912 6529
rect 840 6460 912 6489
rect 994 6530 1182 6558
rect 994 6490 1010 6530
rect 1051 6514 1182 6530
rect 1399 6546 1450 6575
rect 1562 6613 1608 6646
rect 1562 6579 1568 6613
rect 1602 6579 1608 6613
rect 1692 6613 1738 6646
rect 1692 6584 1698 6613
rect 1562 6546 1608 6579
rect 1690 6579 1698 6584
rect 1732 6584 1738 6613
rect 1850 6613 1896 6646
rect 2024 6630 2070 6646
rect 1732 6579 1740 6584
rect 1051 6490 1066 6514
rect 1399 6500 1449 6546
rect 1690 6500 1740 6579
rect 1850 6579 1856 6613
rect 1890 6579 1896 6613
rect 1850 6546 1896 6579
rect 2014 6578 2020 6630
rect 2072 6578 2078 6630
rect 2182 6613 2228 6646
rect 2182 6579 2188 6613
rect 2222 6579 2228 6613
rect 2024 6546 2070 6578
rect 2182 6546 2228 6579
rect 2366 6613 2412 6646
rect 2524 6628 2570 6646
rect 2366 6579 2372 6613
rect 2406 6579 2412 6613
rect 2366 6546 2412 6579
rect 2516 6576 2522 6628
rect 2574 6576 2580 6628
rect 2524 6546 2570 6576
rect 2024 6514 2068 6546
rect 2612 6514 2656 6706
rect 994 6460 1066 6490
rect 1324 6445 1960 6500
rect 2024 6470 2656 6514
rect 2694 6706 2802 6750
rect 2832 6736 2904 6746
rect 2694 6508 2738 6706
rect 2832 6684 2842 6736
rect 2894 6684 2904 6736
rect 2832 6674 2904 6684
rect 2933 6646 2972 6784
rect 3118 6646 3157 6784
rect 3272 6740 3316 6784
rect 3268 6734 3320 6740
rect 3555 6709 3561 6761
rect 3613 6754 3619 6761
rect 3662 6754 3713 6766
rect 3613 6751 3713 6754
rect 3613 6717 3670 6751
rect 3704 6717 3713 6751
rect 3613 6715 3713 6717
rect 3613 6709 3619 6715
rect 3662 6703 3713 6715
rect 3897 6745 3936 6794
rect 3976 6752 4027 6757
rect 3970 6745 3976 6752
rect 3897 6706 3976 6745
rect 3268 6676 3320 6682
rect 3897 6656 3936 6706
rect 3970 6700 3976 6706
rect 4028 6700 4034 6752
rect 4206 6738 4245 6794
rect 4300 6738 4347 6749
rect 4206 6736 4347 6738
rect 4206 6703 4306 6736
rect 3976 6694 4027 6700
rect 4206 6656 4245 6703
rect 4300 6702 4306 6703
rect 4340 6702 4347 6736
rect 4300 6690 4347 6702
rect 2766 6640 2818 6646
rect 2766 6582 2776 6588
rect 2770 6579 2776 6582
rect 2810 6582 2818 6588
rect 2928 6613 2974 6646
rect 2810 6579 2816 6582
rect 2770 6546 2816 6579
rect 2928 6579 2934 6613
rect 2968 6579 2974 6613
rect 2928 6546 2974 6579
rect 3114 6613 3160 6646
rect 3114 6579 3120 6613
rect 3154 6579 3160 6613
rect 3114 6546 3160 6579
rect 3272 6613 3318 6646
rect 3272 6579 3278 6613
rect 3312 6579 3318 6613
rect 3272 6546 3318 6579
rect 3274 6508 3318 6546
rect 2694 6464 3318 6508
rect 3736 6623 3782 6656
rect 3736 6589 3742 6623
rect 3776 6589 3782 6623
rect 3736 6556 3782 6589
rect 3894 6623 3940 6656
rect 3894 6589 3900 6623
rect 3934 6589 3940 6623
rect 4044 6623 4090 6656
rect 4044 6594 4050 6623
rect 3894 6556 3940 6589
rect 4042 6589 4050 6594
rect 4084 6589 4090 6623
rect 4042 6556 4090 6589
rect 4202 6623 4248 6656
rect 4202 6589 4208 6623
rect 4242 6589 4248 6623
rect 4202 6556 4248 6589
rect 3736 6500 3780 6556
rect 4042 6500 4089 6556
rect 1324 6393 1360 6445
rect 1412 6393 1424 6445
rect 1476 6436 1488 6445
rect 1540 6436 1552 6445
rect 1604 6436 1616 6445
rect 1668 6436 1680 6445
rect 1732 6436 1744 6445
rect 1796 6436 1808 6445
rect 1479 6402 1488 6436
rect 1551 6402 1552 6436
rect 1732 6402 1733 6436
rect 1796 6402 1805 6436
rect 1476 6393 1488 6402
rect 1540 6393 1552 6402
rect 1604 6393 1616 6402
rect 1668 6393 1680 6402
rect 1732 6393 1744 6402
rect 1796 6393 1808 6402
rect 1860 6393 1872 6445
rect 1924 6393 1960 6445
rect 3704 6456 4244 6500
rect 3704 6447 3756 6456
rect 3808 6447 3820 6456
rect 1324 6360 1960 6393
rect 2346 6415 2426 6440
rect 2346 6411 3517 6415
rect 2346 6377 2369 6411
rect 2403 6377 3517 6411
rect 2346 6373 3517 6377
rect 2346 6348 2426 6373
rect 2636 6315 2702 6327
rect 272 6261 278 6315
rect 332 6261 2642 6315
rect 2696 6261 2702 6315
rect 2636 6249 2702 6261
rect 3475 6220 3517 6373
rect 3704 6413 3741 6447
rect 3808 6413 3813 6447
rect 3704 6404 3756 6413
rect 3808 6404 3820 6413
rect 3872 6404 3884 6456
rect 3936 6404 3948 6456
rect 4000 6404 4012 6456
rect 4064 6404 4076 6456
rect 4128 6447 4140 6456
rect 4192 6447 4244 6456
rect 4135 6413 4140 6447
rect 4207 6413 4244 6447
rect 4128 6404 4140 6413
rect 4192 6404 4244 6413
rect 3704 6360 4244 6404
rect 3559 6255 3565 6307
rect 3617 6300 3623 6307
rect 4306 6300 4345 6690
rect 4558 6658 4597 6794
rect 4628 6763 4680 6769
rect 4625 6714 4628 6760
rect 4680 6714 4683 6760
rect 4875 6718 4904 6794
rect 4628 6705 4680 6711
rect 4875 6690 4980 6718
rect 4396 6625 4442 6658
rect 4396 6591 4402 6625
rect 4436 6591 4442 6625
rect 4396 6558 4442 6591
rect 4554 6638 4600 6658
rect 4704 6638 4750 6658
rect 4862 6638 4908 6658
rect 4554 6625 4750 6638
rect 4554 6591 4560 6625
rect 4594 6591 4710 6625
rect 4744 6591 4750 6625
rect 4554 6572 4750 6591
rect 4856 6586 4862 6638
rect 4914 6586 4920 6638
rect 4554 6558 4600 6572
rect 4704 6558 4750 6572
rect 4862 6558 4908 6586
rect 4402 6408 4430 6558
rect 4558 6513 4597 6558
rect 4552 6507 4604 6513
rect 4552 6449 4604 6455
rect 4952 6408 4980 6690
rect 5026 6640 5056 6825
rect 5694 6794 5740 6842
rect 5852 6948 5898 6994
rect 5852 6914 5858 6948
rect 5892 6914 5898 6948
rect 5852 6876 5898 6914
rect 5852 6842 5858 6876
rect 5892 6842 5898 6876
rect 5852 6794 5898 6842
rect 6002 6948 6048 7050
rect 6516 6994 6556 7200
rect 6862 7194 6868 7200
rect 6920 7194 6926 7246
rect 6985 7234 7015 7287
rect 6985 7205 7016 7234
rect 6002 6914 6008 6948
rect 6042 6914 6048 6948
rect 6002 6876 6048 6914
rect 6002 6842 6008 6876
rect 6042 6842 6048 6876
rect 6002 6794 6048 6842
rect 6160 6948 6206 6994
rect 6160 6914 6166 6948
rect 6200 6914 6206 6948
rect 6354 6948 6400 6994
rect 6354 6922 6360 6948
rect 6160 6876 6206 6914
rect 6160 6842 6166 6876
rect 6200 6842 6206 6876
rect 6244 6920 6360 6922
rect 6244 6868 6250 6920
rect 6302 6914 6360 6920
rect 6394 6914 6400 6948
rect 6302 6876 6400 6914
rect 6302 6868 6360 6876
rect 6244 6866 6360 6868
rect 6160 6794 6206 6842
rect 6354 6842 6360 6866
rect 6394 6842 6400 6876
rect 6354 6794 6400 6842
rect 6512 6948 6558 6994
rect 6512 6914 6518 6948
rect 6552 6914 6558 6948
rect 6662 6948 6708 6994
rect 6662 6914 6668 6948
rect 6702 6914 6708 6948
rect 6512 6876 6708 6914
rect 6512 6842 6518 6876
rect 6552 6848 6668 6876
rect 6552 6842 6558 6848
rect 6512 6794 6558 6842
rect 6662 6842 6668 6848
rect 6702 6842 6708 6876
rect 6662 6794 6708 6842
rect 6820 6948 6866 6994
rect 6820 6914 6826 6948
rect 6860 6914 6866 6948
rect 6986 6918 7016 7205
rect 6820 6876 6866 6914
rect 6820 6842 6826 6876
rect 6860 6842 6866 6876
rect 6968 6866 6974 6918
rect 7026 6866 7032 6918
rect 6820 6794 6866 6842
rect 6984 6826 7016 6866
rect 5111 6709 5117 6761
rect 5169 6754 5175 6761
rect 5620 6754 5672 6766
rect 5169 6752 5672 6754
rect 5169 6718 5628 6752
rect 5662 6718 5672 6752
rect 5169 6715 5672 6718
rect 5169 6709 5175 6715
rect 5620 6704 5672 6715
rect 5856 6746 5894 6794
rect 5934 6752 5986 6758
rect 5928 6746 5934 6752
rect 5856 6706 5934 6746
rect 5856 6656 5894 6706
rect 5928 6700 5934 6706
rect 5986 6700 5992 6752
rect 6164 6738 6204 6794
rect 6258 6738 6306 6750
rect 6164 6736 6306 6738
rect 6164 6704 6264 6736
rect 5934 6694 5986 6700
rect 6164 6656 6204 6704
rect 6258 6702 6264 6704
rect 6298 6702 6306 6736
rect 6258 6690 6306 6702
rect 5009 6588 5015 6640
rect 5067 6588 5073 6640
rect 5694 6624 5740 6656
rect 5694 6590 5700 6624
rect 5734 6590 5740 6624
rect 4402 6380 4980 6408
rect 3617 6261 4345 6300
rect 3617 6255 3623 6261
rect 5021 6220 5063 6588
rect 5694 6556 5740 6590
rect 5852 6624 5898 6656
rect 5852 6590 5858 6624
rect 5892 6590 5898 6624
rect 6002 6624 6048 6656
rect 6002 6594 6008 6624
rect 5852 6556 5898 6590
rect 6000 6590 6008 6594
rect 6042 6590 6048 6624
rect 5694 6500 5738 6556
rect 6000 6500 6048 6590
rect 6160 6624 6206 6656
rect 6160 6590 6166 6624
rect 6200 6590 6206 6624
rect 6160 6556 6206 6590
rect 5662 6456 6202 6500
rect 5662 6448 5714 6456
rect 5766 6448 5778 6456
rect 5662 6414 5700 6448
rect 5766 6414 5772 6448
rect 5662 6404 5714 6414
rect 5766 6404 5778 6414
rect 5830 6404 5842 6456
rect 5894 6404 5906 6456
rect 5958 6404 5970 6456
rect 6022 6404 6034 6456
rect 6086 6448 6098 6456
rect 6150 6448 6202 6456
rect 6094 6414 6098 6448
rect 6166 6414 6202 6448
rect 6086 6404 6098 6414
rect 6150 6404 6202 6414
rect 5662 6360 6202 6404
rect 5111 6255 5117 6307
rect 5169 6300 5175 6307
rect 6264 6300 6304 6690
rect 6516 6658 6556 6794
rect 6586 6764 6638 6770
rect 6584 6714 6586 6760
rect 6638 6714 6642 6760
rect 6834 6718 6862 6794
rect 6586 6706 6638 6712
rect 6834 6690 6936 6718
rect 6354 6626 6400 6658
rect 6354 6592 6360 6626
rect 6394 6592 6400 6626
rect 6354 6558 6400 6592
rect 6512 6638 6558 6658
rect 6662 6638 6708 6658
rect 6820 6638 6866 6658
rect 6512 6626 6708 6638
rect 6512 6592 6518 6626
rect 6552 6592 6668 6626
rect 6702 6592 6708 6626
rect 6512 6572 6708 6592
rect 6814 6586 6820 6638
rect 6872 6586 6878 6638
rect 6512 6558 6558 6572
rect 6662 6558 6708 6572
rect 6820 6558 6866 6586
rect 6360 6408 6388 6558
rect 6516 6514 6556 6558
rect 6510 6508 6562 6514
rect 6510 6450 6562 6456
rect 6908 6408 6936 6690
rect 6984 6640 7014 6826
rect 6968 6588 6974 6640
rect 7026 6588 7032 6640
rect 6360 6380 6936 6408
rect 6908 6316 6936 6380
rect 5169 6262 6304 6300
rect 6346 6288 6936 6316
rect 5169 6261 5572 6262
rect 5169 6255 5175 6261
rect 3475 6178 5063 6220
rect 5035 6137 5087 6143
rect 3472 6053 4907 6092
rect 6346 6125 6374 6288
rect 6908 6286 6936 6288
rect 5087 6097 6374 6125
rect 6968 6086 6974 6138
rect 7026 6086 7032 6138
rect 5035 6079 5087 6085
rect 1348 5919 1880 5962
rect 1348 5910 1398 5919
rect 1450 5910 1462 5919
rect 1348 5876 1383 5910
rect 1450 5876 1455 5910
rect 1348 5867 1398 5876
rect 1450 5867 1462 5876
rect 1514 5867 1526 5919
rect 1578 5867 1590 5919
rect 1642 5867 1654 5919
rect 1706 5867 1718 5919
rect 1770 5910 1782 5919
rect 1834 5910 1880 5919
rect 1777 5876 1782 5910
rect 1849 5876 1880 5910
rect 3472 5895 3511 6053
rect 4738 6011 4744 6018
rect 4558 5972 4744 6011
rect 1770 5867 1782 5876
rect 1834 5867 1880 5876
rect 550 5848 622 5852
rect 550 5796 560 5848
rect 612 5796 622 5848
rect 696 5846 768 5852
rect 550 5784 566 5796
rect 607 5784 622 5796
rect 682 5844 768 5846
rect 682 5792 702 5844
rect 754 5792 768 5844
rect 682 5790 710 5792
rect 550 5754 622 5784
rect 696 5784 710 5790
rect 751 5784 768 5792
rect 696 5754 768 5784
rect 840 5829 912 5858
rect 840 5789 856 5829
rect 897 5789 912 5829
rect 840 5760 912 5789
rect 994 5829 1066 5858
rect 994 5789 1009 5829
rect 1050 5789 1066 5829
rect 1348 5822 1880 5867
rect 994 5760 1066 5789
rect 564 5714 608 5754
rect 856 5694 900 5760
rect 378 5686 433 5692
rect 846 5642 852 5694
rect 904 5642 910 5694
rect 378 5401 433 5631
rect 856 5602 900 5642
rect 1008 5602 1052 5760
rect 1407 5756 1448 5822
rect 1693 5756 1735 5822
rect 1941 5819 2687 5864
rect 1404 5709 1450 5756
rect 1404 5675 1410 5709
rect 1444 5675 1450 5709
rect 1404 5637 1450 5675
rect 1404 5603 1410 5637
rect 1444 5603 1450 5637
rect 708 5558 900 5602
rect 372 5346 378 5401
rect 433 5346 439 5401
rect 708 5324 752 5558
rect 998 5550 1004 5602
rect 1056 5550 1062 5602
rect 1404 5556 1450 5603
rect 1562 5709 1608 5756
rect 1562 5675 1568 5709
rect 1602 5675 1608 5709
rect 1562 5637 1608 5675
rect 1562 5603 1568 5637
rect 1602 5603 1608 5637
rect 1562 5556 1608 5603
rect 1692 5709 1738 5756
rect 1692 5675 1698 5709
rect 1732 5675 1738 5709
rect 1692 5637 1738 5675
rect 1692 5603 1698 5637
rect 1732 5603 1738 5637
rect 1692 5556 1738 5603
rect 1850 5753 1896 5756
rect 1941 5753 1986 5819
rect 1850 5709 1986 5753
rect 1850 5675 1856 5709
rect 1890 5708 1986 5709
rect 2024 5709 2070 5756
rect 1890 5675 1896 5708
rect 1850 5637 1896 5675
rect 2024 5675 2030 5709
rect 2064 5675 2070 5709
rect 2024 5640 2070 5675
rect 1998 5638 2070 5640
rect 1850 5603 1856 5637
rect 1890 5603 1896 5637
rect 1850 5556 1896 5603
rect 1928 5637 2070 5638
rect 1928 5613 2030 5637
rect 1928 5596 1935 5613
rect 1929 5561 1935 5596
rect 1987 5603 2030 5613
rect 2064 5603 2070 5637
rect 1987 5596 2070 5603
rect 1987 5561 1993 5596
rect 2024 5556 2070 5596
rect 2182 5712 2228 5756
rect 2366 5712 2412 5756
rect 2182 5709 2412 5712
rect 2182 5675 2188 5709
rect 2222 5675 2372 5709
rect 2406 5675 2412 5709
rect 2182 5637 2412 5675
rect 2182 5603 2188 5637
rect 2222 5603 2372 5637
rect 2406 5603 2412 5637
rect 2182 5586 2412 5603
rect 2182 5556 2228 5586
rect 2366 5556 2412 5586
rect 2524 5709 2570 5756
rect 2524 5675 2530 5709
rect 2564 5675 2570 5709
rect 2642 5685 2687 5819
rect 3118 5856 3511 5895
rect 3724 5918 4264 5962
rect 3724 5866 3776 5918
rect 3828 5909 3840 5918
rect 3892 5909 3904 5918
rect 3956 5909 3968 5918
rect 4020 5909 4032 5918
rect 4084 5909 4096 5918
rect 4148 5909 4160 5918
rect 3831 5875 3840 5909
rect 3903 5875 3904 5909
rect 4084 5875 4085 5909
rect 4148 5875 4157 5909
rect 3828 5866 3840 5875
rect 3892 5866 3904 5875
rect 3956 5866 3968 5875
rect 4020 5866 4032 5875
rect 4084 5866 4096 5875
rect 4148 5866 4160 5875
rect 4212 5866 4264 5918
rect 2774 5812 2816 5813
rect 2758 5804 2816 5812
rect 2758 5752 2769 5804
rect 2821 5752 2827 5804
rect 3118 5756 3157 5856
rect 3724 5822 4264 5866
rect 3741 5766 3787 5822
rect 3736 5765 3787 5766
rect 2758 5709 2816 5752
rect 2524 5637 2570 5675
rect 2524 5603 2530 5637
rect 2564 5603 2570 5637
rect 2524 5596 2570 5603
rect 2613 5657 2715 5685
rect 2613 5623 2647 5657
rect 2681 5623 2715 5657
rect 2524 5556 2574 5596
rect 2613 5595 2715 5623
rect 2758 5675 2776 5709
rect 2810 5675 2816 5709
rect 2758 5637 2816 5675
rect 2758 5603 2776 5637
rect 2810 5603 2816 5637
rect 1008 5496 1052 5550
rect 1245 5515 1328 5534
rect 852 5452 1052 5496
rect 1148 5513 1328 5515
rect 1148 5461 1155 5513
rect 1207 5503 1328 5513
rect 1207 5469 1269 5503
rect 1303 5469 1328 5503
rect 1207 5461 1328 5469
rect 1148 5460 1328 5461
rect 852 5330 896 5452
rect 1245 5439 1328 5460
rect 1568 5522 1602 5556
rect 1568 5512 1820 5522
rect 1568 5460 1758 5512
rect 1810 5460 1820 5512
rect 1568 5450 1820 5460
rect 1568 5418 1608 5450
rect 1853 5418 1892 5556
rect 2185 5418 2224 5556
rect 2255 5519 2325 5525
rect 2255 5510 2331 5519
rect 2255 5458 2270 5510
rect 2322 5458 2331 5510
rect 2255 5449 2331 5458
rect 2255 5443 2325 5449
rect 2368 5418 2407 5556
rect 2530 5522 2574 5556
rect 2758 5556 2816 5603
rect 2928 5709 2974 5756
rect 2928 5675 2934 5709
rect 2968 5696 2974 5709
rect 3114 5709 3160 5756
rect 3114 5696 3120 5709
rect 2968 5675 3120 5696
rect 3154 5675 3160 5709
rect 3272 5709 3318 5756
rect 3272 5699 3278 5709
rect 3312 5699 3318 5709
rect 3736 5719 3782 5765
rect 2928 5637 3160 5675
rect 3262 5647 3268 5699
rect 3320 5647 3326 5699
rect 3736 5685 3742 5719
rect 3776 5685 3782 5719
rect 3736 5647 3782 5685
rect 2928 5603 2934 5637
rect 2968 5603 3120 5637
rect 3154 5603 3160 5637
rect 2928 5586 3160 5603
rect 2928 5556 2974 5586
rect 3114 5556 3160 5586
rect 3272 5637 3318 5647
rect 3272 5603 3278 5637
rect 3312 5603 3318 5637
rect 3272 5556 3318 5603
rect 3736 5613 3742 5647
rect 3776 5613 3782 5647
rect 3736 5566 3782 5613
rect 3894 5719 3940 5766
rect 3894 5685 3900 5719
rect 3934 5685 3940 5719
rect 3894 5647 3940 5685
rect 3894 5613 3900 5647
rect 3934 5613 3940 5647
rect 3894 5566 3940 5613
rect 4044 5719 4090 5822
rect 4558 5766 4597 5972
rect 4738 5966 4744 5972
rect 4796 5966 4802 6018
rect 4868 5766 4907 6053
rect 5682 5918 6222 5962
rect 5682 5866 5734 5918
rect 5786 5908 5798 5918
rect 5850 5908 5862 5918
rect 5914 5908 5926 5918
rect 5978 5908 5990 5918
rect 6042 5908 6054 5918
rect 6106 5908 6118 5918
rect 5790 5874 5798 5908
rect 6042 5874 6044 5908
rect 6106 5874 6116 5908
rect 5786 5866 5798 5874
rect 5850 5866 5862 5874
rect 5914 5866 5926 5874
rect 5978 5866 5990 5874
rect 6042 5866 6054 5874
rect 6106 5866 6118 5874
rect 6170 5866 6222 5918
rect 5682 5822 6222 5866
rect 5700 5766 5746 5822
rect 4044 5685 4050 5719
rect 4084 5685 4090 5719
rect 4044 5647 4090 5685
rect 4044 5613 4050 5647
rect 4084 5613 4090 5647
rect 4044 5566 4090 5613
rect 4202 5719 4248 5766
rect 4202 5685 4208 5719
rect 4242 5685 4248 5719
rect 4396 5719 4442 5766
rect 4396 5693 4402 5719
rect 4202 5647 4248 5685
rect 4202 5613 4208 5647
rect 4242 5613 4248 5647
rect 4285 5691 4402 5693
rect 4285 5639 4292 5691
rect 4344 5685 4402 5691
rect 4436 5685 4442 5719
rect 4344 5647 4442 5685
rect 4344 5639 4402 5647
rect 4285 5638 4402 5639
rect 4202 5566 4248 5613
rect 4396 5613 4402 5638
rect 4436 5613 4442 5647
rect 4396 5566 4442 5613
rect 4554 5719 4600 5766
rect 4554 5685 4560 5719
rect 4594 5686 4600 5719
rect 4704 5719 4750 5766
rect 4704 5686 4710 5719
rect 4594 5685 4710 5686
rect 4744 5685 4750 5719
rect 4554 5647 4750 5685
rect 4554 5613 4560 5647
rect 4594 5620 4710 5647
rect 4594 5613 4600 5620
rect 4554 5566 4600 5613
rect 4704 5613 4710 5620
rect 4744 5613 4750 5647
rect 4704 5566 4750 5613
rect 4862 5719 4908 5766
rect 4862 5685 4868 5719
rect 4902 5685 4908 5719
rect 5694 5720 5740 5766
rect 5027 5690 5057 5699
rect 4862 5647 4908 5685
rect 4862 5613 4868 5647
rect 4902 5613 4908 5647
rect 5010 5638 5016 5690
rect 5068 5638 5074 5690
rect 5694 5686 5700 5720
rect 5734 5686 5740 5720
rect 5694 5648 5740 5686
rect 4862 5566 4908 5613
rect 5026 5597 5057 5638
rect 5694 5614 5700 5648
rect 5734 5614 5740 5648
rect 2758 5522 2802 5556
rect 2530 5478 2656 5522
rect 1242 5398 1248 5402
rect 1138 5354 1248 5398
rect 1138 5330 1182 5354
rect 1242 5350 1248 5354
rect 1300 5350 1306 5402
rect 1404 5385 1450 5418
rect 1404 5351 1410 5385
rect 1444 5351 1450 5385
rect 1404 5347 1450 5351
rect 378 5302 434 5308
rect 550 5302 622 5324
rect 434 5296 622 5302
rect 434 5256 565 5296
rect 606 5256 622 5296
rect 434 5246 622 5256
rect 378 5240 434 5246
rect 550 5226 622 5246
rect 696 5296 768 5324
rect 696 5256 712 5296
rect 753 5256 768 5296
rect 696 5226 768 5256
rect 840 5301 912 5330
rect 840 5261 856 5301
rect 897 5261 912 5301
rect 840 5232 912 5261
rect 994 5302 1182 5330
rect 994 5262 1010 5302
rect 1051 5286 1182 5302
rect 1399 5318 1450 5347
rect 1562 5385 1608 5418
rect 1562 5351 1568 5385
rect 1602 5351 1608 5385
rect 1692 5385 1738 5418
rect 1692 5356 1698 5385
rect 1562 5318 1608 5351
rect 1690 5351 1698 5356
rect 1732 5356 1738 5385
rect 1850 5385 1896 5418
rect 2024 5402 2070 5418
rect 1732 5351 1740 5356
rect 1051 5262 1066 5286
rect 1399 5272 1449 5318
rect 1690 5272 1740 5351
rect 1850 5351 1856 5385
rect 1890 5351 1896 5385
rect 1850 5318 1896 5351
rect 2014 5350 2020 5402
rect 2072 5350 2078 5402
rect 2182 5385 2228 5418
rect 2182 5351 2188 5385
rect 2222 5351 2228 5385
rect 2024 5318 2070 5350
rect 2182 5318 2228 5351
rect 2366 5385 2412 5418
rect 2524 5400 2570 5418
rect 2366 5351 2372 5385
rect 2406 5351 2412 5385
rect 2366 5318 2412 5351
rect 2516 5348 2522 5400
rect 2574 5348 2580 5400
rect 2524 5318 2570 5348
rect 2024 5286 2068 5318
rect 2612 5286 2656 5478
rect 994 5232 1066 5262
rect 1324 5217 1960 5272
rect 2024 5242 2656 5286
rect 2694 5478 2802 5522
rect 2832 5508 2904 5518
rect 2694 5280 2738 5478
rect 2832 5456 2842 5508
rect 2894 5456 2904 5508
rect 2832 5446 2904 5456
rect 2933 5418 2972 5556
rect 3118 5418 3157 5556
rect 3272 5512 3316 5556
rect 3268 5506 3320 5512
rect 3555 5481 3561 5533
rect 3613 5526 3619 5533
rect 3662 5526 3713 5538
rect 3613 5523 3713 5526
rect 3613 5489 3670 5523
rect 3704 5489 3713 5523
rect 3613 5487 3713 5489
rect 3613 5481 3619 5487
rect 3662 5475 3713 5487
rect 3897 5517 3936 5566
rect 3976 5524 4027 5529
rect 3970 5517 3976 5524
rect 3897 5478 3976 5517
rect 3268 5448 3320 5454
rect 3897 5428 3936 5478
rect 3970 5472 3976 5478
rect 4028 5472 4034 5524
rect 4206 5510 4245 5566
rect 4300 5510 4347 5521
rect 4206 5508 4347 5510
rect 4206 5475 4306 5508
rect 3976 5466 4027 5472
rect 4206 5428 4245 5475
rect 4300 5474 4306 5475
rect 4340 5474 4347 5508
rect 4300 5462 4347 5474
rect 2766 5412 2818 5418
rect 2766 5354 2776 5360
rect 2770 5351 2776 5354
rect 2810 5354 2818 5360
rect 2928 5385 2974 5418
rect 2810 5351 2816 5354
rect 2770 5318 2816 5351
rect 2928 5351 2934 5385
rect 2968 5351 2974 5385
rect 2928 5318 2974 5351
rect 3114 5385 3160 5418
rect 3114 5351 3120 5385
rect 3154 5351 3160 5385
rect 3114 5318 3160 5351
rect 3272 5385 3318 5418
rect 3272 5351 3278 5385
rect 3312 5351 3318 5385
rect 3272 5318 3318 5351
rect 3274 5280 3318 5318
rect 2694 5236 3318 5280
rect 3736 5395 3782 5428
rect 3736 5361 3742 5395
rect 3776 5361 3782 5395
rect 3736 5328 3782 5361
rect 3894 5395 3940 5428
rect 3894 5361 3900 5395
rect 3934 5361 3940 5395
rect 4044 5395 4090 5428
rect 4044 5366 4050 5395
rect 3894 5328 3940 5361
rect 4042 5361 4050 5366
rect 4084 5361 4090 5395
rect 4042 5328 4090 5361
rect 4202 5395 4248 5428
rect 4202 5361 4208 5395
rect 4242 5361 4248 5395
rect 4202 5328 4248 5361
rect 3736 5272 3780 5328
rect 4042 5272 4089 5328
rect 1324 5165 1360 5217
rect 1412 5165 1424 5217
rect 1476 5208 1488 5217
rect 1540 5208 1552 5217
rect 1604 5208 1616 5217
rect 1668 5208 1680 5217
rect 1732 5208 1744 5217
rect 1796 5208 1808 5217
rect 1479 5174 1488 5208
rect 1551 5174 1552 5208
rect 1732 5174 1733 5208
rect 1796 5174 1805 5208
rect 1476 5165 1488 5174
rect 1540 5165 1552 5174
rect 1604 5165 1616 5174
rect 1668 5165 1680 5174
rect 1732 5165 1744 5174
rect 1796 5165 1808 5174
rect 1860 5165 1872 5217
rect 1924 5165 1960 5217
rect 3704 5228 4244 5272
rect 3704 5219 3756 5228
rect 3808 5219 3820 5228
rect 1324 5132 1960 5165
rect 2346 5187 2426 5212
rect 2346 5183 3517 5187
rect 2346 5149 2369 5183
rect 2403 5149 3517 5183
rect 2346 5145 3517 5149
rect 2346 5120 2426 5145
rect 2636 5087 2702 5099
rect 272 5033 278 5087
rect 332 5033 2642 5087
rect 2696 5033 2702 5087
rect 2636 5021 2702 5033
rect 3475 4992 3517 5145
rect 3704 5185 3741 5219
rect 3808 5185 3813 5219
rect 3704 5176 3756 5185
rect 3808 5176 3820 5185
rect 3872 5176 3884 5228
rect 3936 5176 3948 5228
rect 4000 5176 4012 5228
rect 4064 5176 4076 5228
rect 4128 5219 4140 5228
rect 4192 5219 4244 5228
rect 4135 5185 4140 5219
rect 4207 5185 4244 5219
rect 4128 5176 4140 5185
rect 4192 5176 4244 5185
rect 3704 5132 4244 5176
rect 3559 5027 3565 5079
rect 3617 5072 3623 5079
rect 4306 5072 4345 5462
rect 4558 5430 4597 5566
rect 4628 5535 4680 5541
rect 4625 5486 4628 5532
rect 4680 5486 4683 5532
rect 4875 5490 4904 5566
rect 4628 5477 4680 5483
rect 4875 5462 4980 5490
rect 4396 5397 4442 5430
rect 4396 5363 4402 5397
rect 4436 5363 4442 5397
rect 4396 5330 4442 5363
rect 4554 5410 4600 5430
rect 4704 5410 4750 5430
rect 4862 5410 4908 5430
rect 4554 5397 4750 5410
rect 4554 5363 4560 5397
rect 4594 5363 4710 5397
rect 4744 5363 4750 5397
rect 4554 5344 4750 5363
rect 4856 5358 4862 5410
rect 4914 5358 4920 5410
rect 4554 5330 4600 5344
rect 4704 5330 4750 5344
rect 4862 5330 4908 5358
rect 4402 5180 4430 5330
rect 4558 5285 4597 5330
rect 4552 5279 4604 5285
rect 4552 5221 4604 5227
rect 4952 5180 4980 5462
rect 5026 5412 5056 5597
rect 5694 5566 5740 5614
rect 5852 5720 5898 5766
rect 5852 5686 5858 5720
rect 5892 5686 5898 5720
rect 5852 5648 5898 5686
rect 5852 5614 5858 5648
rect 5892 5614 5898 5648
rect 5852 5566 5898 5614
rect 6002 5720 6048 5822
rect 6516 5766 6556 6010
rect 6985 6006 7015 6086
rect 6985 5977 7016 6006
rect 6002 5686 6008 5720
rect 6042 5686 6048 5720
rect 6002 5648 6048 5686
rect 6002 5614 6008 5648
rect 6042 5614 6048 5648
rect 6002 5566 6048 5614
rect 6160 5720 6206 5766
rect 6160 5686 6166 5720
rect 6200 5686 6206 5720
rect 6354 5720 6400 5766
rect 6354 5694 6360 5720
rect 6160 5648 6206 5686
rect 6160 5614 6166 5648
rect 6200 5614 6206 5648
rect 6244 5692 6360 5694
rect 6244 5640 6250 5692
rect 6302 5686 6360 5692
rect 6394 5686 6400 5720
rect 6302 5648 6400 5686
rect 6302 5640 6360 5648
rect 6244 5638 6360 5640
rect 6160 5566 6206 5614
rect 6354 5614 6360 5638
rect 6394 5614 6400 5648
rect 6354 5566 6400 5614
rect 6512 5720 6558 5766
rect 6512 5686 6518 5720
rect 6552 5686 6558 5720
rect 6662 5720 6708 5766
rect 6662 5686 6668 5720
rect 6702 5686 6708 5720
rect 6512 5648 6708 5686
rect 6512 5614 6518 5648
rect 6552 5620 6668 5648
rect 6552 5614 6558 5620
rect 6512 5566 6558 5614
rect 6662 5614 6668 5620
rect 6702 5614 6708 5648
rect 6662 5566 6708 5614
rect 6820 5720 6866 5766
rect 6820 5686 6826 5720
rect 6860 5686 6866 5720
rect 6986 5690 7016 5977
rect 6820 5648 6866 5686
rect 6820 5614 6826 5648
rect 6860 5614 6866 5648
rect 6968 5638 6974 5690
rect 7026 5638 7032 5690
rect 6820 5566 6866 5614
rect 6984 5598 7016 5638
rect 5273 5481 5279 5533
rect 5331 5526 5337 5533
rect 5620 5526 5672 5538
rect 5331 5524 5672 5526
rect 5331 5490 5628 5524
rect 5662 5490 5672 5524
rect 5331 5487 5672 5490
rect 5331 5481 5337 5487
rect 5620 5476 5672 5487
rect 5856 5518 5894 5566
rect 5934 5524 5986 5530
rect 5928 5518 5934 5524
rect 5856 5478 5934 5518
rect 5856 5428 5894 5478
rect 5928 5472 5934 5478
rect 5986 5472 5992 5524
rect 6164 5510 6204 5566
rect 6258 5510 6306 5522
rect 6164 5508 6306 5510
rect 6164 5476 6264 5508
rect 5934 5466 5986 5472
rect 6164 5428 6204 5476
rect 6258 5474 6264 5476
rect 6298 5474 6306 5508
rect 6258 5462 6306 5474
rect 5009 5360 5015 5412
rect 5067 5360 5073 5412
rect 5694 5396 5740 5428
rect 5694 5362 5700 5396
rect 5734 5362 5740 5396
rect 4402 5152 4980 5180
rect 3617 5033 4345 5072
rect 3617 5027 3623 5033
rect 5021 4992 5063 5360
rect 5694 5328 5740 5362
rect 5852 5396 5898 5428
rect 5852 5362 5858 5396
rect 5892 5362 5898 5396
rect 6002 5396 6048 5428
rect 6002 5366 6008 5396
rect 5852 5328 5898 5362
rect 6000 5362 6008 5366
rect 6042 5362 6048 5396
rect 5694 5272 5738 5328
rect 6000 5272 6048 5362
rect 6160 5396 6206 5428
rect 6160 5362 6166 5396
rect 6200 5362 6206 5396
rect 6160 5328 6206 5362
rect 5662 5228 6202 5272
rect 5662 5220 5714 5228
rect 5766 5220 5778 5228
rect 5662 5186 5700 5220
rect 5766 5186 5772 5220
rect 5662 5176 5714 5186
rect 5766 5176 5778 5186
rect 5830 5176 5842 5228
rect 5894 5176 5906 5228
rect 5958 5176 5970 5228
rect 6022 5176 6034 5228
rect 6086 5220 6098 5228
rect 6150 5220 6202 5228
rect 6094 5186 6098 5220
rect 6166 5186 6202 5220
rect 6086 5176 6098 5186
rect 6150 5176 6202 5186
rect 5662 5132 6202 5176
rect 5273 5027 5279 5079
rect 5331 5072 5337 5079
rect 6264 5072 6304 5462
rect 6516 5430 6556 5566
rect 6586 5536 6638 5542
rect 6584 5486 6586 5532
rect 6638 5486 6642 5532
rect 6834 5490 6862 5566
rect 6586 5478 6638 5484
rect 6834 5462 6936 5490
rect 6354 5398 6400 5430
rect 6354 5364 6360 5398
rect 6394 5364 6400 5398
rect 6354 5330 6400 5364
rect 6512 5410 6558 5430
rect 6662 5410 6708 5430
rect 6820 5410 6866 5430
rect 6512 5398 6708 5410
rect 6512 5364 6518 5398
rect 6552 5364 6668 5398
rect 6702 5364 6708 5398
rect 6512 5344 6708 5364
rect 6814 5358 6820 5410
rect 6872 5358 6878 5410
rect 6512 5330 6558 5344
rect 6662 5330 6708 5344
rect 6820 5330 6866 5358
rect 6360 5180 6388 5330
rect 6516 5286 6556 5330
rect 6510 5280 6562 5286
rect 6510 5222 6562 5228
rect 6908 5180 6936 5462
rect 6984 5412 7014 5598
rect 6968 5360 6974 5412
rect 7026 5360 7032 5412
rect 6360 5152 6936 5180
rect 5331 5034 6304 5072
rect 5331 5033 5584 5034
rect 5331 5027 5337 5033
rect 3475 4950 5063 4992
rect 6908 4964 6936 5152
rect 6908 4936 7234 4964
rect 5029 4872 5081 4878
rect 3472 4825 4907 4864
rect 1348 4691 1880 4734
rect 1348 4682 1398 4691
rect 1450 4682 1462 4691
rect 1348 4648 1383 4682
rect 1450 4648 1455 4682
rect 1348 4639 1398 4648
rect 1450 4639 1462 4648
rect 1514 4639 1526 4691
rect 1578 4639 1590 4691
rect 1642 4639 1654 4691
rect 1706 4639 1718 4691
rect 1770 4682 1782 4691
rect 1834 4682 1880 4691
rect 1777 4648 1782 4682
rect 1849 4648 1880 4682
rect 3472 4667 3511 4825
rect 4738 4783 4744 4790
rect 4558 4744 4744 4783
rect 1770 4639 1782 4648
rect 1834 4639 1880 4648
rect 550 4620 622 4624
rect 550 4568 560 4620
rect 612 4568 622 4620
rect 696 4618 768 4624
rect 550 4556 566 4568
rect 607 4556 622 4568
rect 682 4616 768 4618
rect 682 4564 702 4616
rect 754 4564 768 4616
rect 682 4562 710 4564
rect 550 4526 622 4556
rect 696 4556 710 4562
rect 751 4556 768 4564
rect 696 4526 768 4556
rect 840 4601 912 4630
rect 840 4561 856 4601
rect 897 4561 912 4601
rect 840 4532 912 4561
rect 994 4601 1066 4630
rect 994 4561 1009 4601
rect 1050 4561 1066 4601
rect 1348 4594 1880 4639
rect 994 4532 1066 4561
rect 564 4486 608 4526
rect 856 4466 900 4532
rect 378 4458 433 4464
rect 846 4414 852 4466
rect 904 4414 910 4466
rect 378 4173 433 4403
rect 856 4374 900 4414
rect 1008 4374 1052 4532
rect 1407 4528 1448 4594
rect 1693 4528 1735 4594
rect 1941 4591 2687 4636
rect 1404 4481 1450 4528
rect 1404 4447 1410 4481
rect 1444 4447 1450 4481
rect 1404 4409 1450 4447
rect 1404 4375 1410 4409
rect 1444 4375 1450 4409
rect 708 4330 900 4374
rect 372 4118 378 4173
rect 433 4118 439 4173
rect 708 4096 752 4330
rect 998 4322 1004 4374
rect 1056 4322 1062 4374
rect 1404 4328 1450 4375
rect 1562 4481 1608 4528
rect 1562 4447 1568 4481
rect 1602 4447 1608 4481
rect 1562 4409 1608 4447
rect 1562 4375 1568 4409
rect 1602 4375 1608 4409
rect 1562 4328 1608 4375
rect 1692 4481 1738 4528
rect 1692 4447 1698 4481
rect 1732 4447 1738 4481
rect 1692 4409 1738 4447
rect 1692 4375 1698 4409
rect 1732 4375 1738 4409
rect 1692 4328 1738 4375
rect 1850 4525 1896 4528
rect 1941 4525 1986 4591
rect 1850 4481 1986 4525
rect 1850 4447 1856 4481
rect 1890 4480 1986 4481
rect 2024 4481 2070 4528
rect 1890 4447 1896 4480
rect 1850 4409 1896 4447
rect 2024 4447 2030 4481
rect 2064 4447 2070 4481
rect 2024 4412 2070 4447
rect 1998 4410 2070 4412
rect 1850 4375 1856 4409
rect 1890 4375 1896 4409
rect 1850 4328 1896 4375
rect 1928 4409 2070 4410
rect 1928 4385 2030 4409
rect 1928 4368 1935 4385
rect 1929 4333 1935 4368
rect 1987 4375 2030 4385
rect 2064 4375 2070 4409
rect 1987 4368 2070 4375
rect 1987 4333 1993 4368
rect 2024 4328 2070 4368
rect 2182 4484 2228 4528
rect 2366 4484 2412 4528
rect 2182 4481 2412 4484
rect 2182 4447 2188 4481
rect 2222 4447 2372 4481
rect 2406 4447 2412 4481
rect 2182 4409 2412 4447
rect 2182 4375 2188 4409
rect 2222 4375 2372 4409
rect 2406 4375 2412 4409
rect 2182 4358 2412 4375
rect 2182 4328 2228 4358
rect 2366 4328 2412 4358
rect 2524 4481 2570 4528
rect 2524 4447 2530 4481
rect 2564 4447 2570 4481
rect 2642 4457 2687 4591
rect 3118 4628 3511 4667
rect 3724 4690 4264 4734
rect 3724 4638 3776 4690
rect 3828 4681 3840 4690
rect 3892 4681 3904 4690
rect 3956 4681 3968 4690
rect 4020 4681 4032 4690
rect 4084 4681 4096 4690
rect 4148 4681 4160 4690
rect 3831 4647 3840 4681
rect 3903 4647 3904 4681
rect 4084 4647 4085 4681
rect 4148 4647 4157 4681
rect 3828 4638 3840 4647
rect 3892 4638 3904 4647
rect 3956 4638 3968 4647
rect 4020 4638 4032 4647
rect 4084 4638 4096 4647
rect 4148 4638 4160 4647
rect 4212 4638 4264 4690
rect 2774 4584 2816 4585
rect 2758 4576 2816 4584
rect 2758 4524 2769 4576
rect 2821 4524 2827 4576
rect 3118 4528 3157 4628
rect 3724 4594 4264 4638
rect 3741 4538 3787 4594
rect 3736 4537 3787 4538
rect 2758 4481 2816 4524
rect 2524 4409 2570 4447
rect 2524 4375 2530 4409
rect 2564 4375 2570 4409
rect 2524 4368 2570 4375
rect 2613 4429 2715 4457
rect 2613 4395 2647 4429
rect 2681 4395 2715 4429
rect 2524 4328 2574 4368
rect 2613 4367 2715 4395
rect 2758 4447 2776 4481
rect 2810 4447 2816 4481
rect 2758 4409 2816 4447
rect 2758 4375 2776 4409
rect 2810 4375 2816 4409
rect 1008 4268 1052 4322
rect 1245 4287 1328 4306
rect 852 4224 1052 4268
rect 1148 4285 1328 4287
rect 1148 4233 1155 4285
rect 1207 4275 1328 4285
rect 1207 4241 1269 4275
rect 1303 4241 1328 4275
rect 1207 4233 1328 4241
rect 1148 4232 1328 4233
rect 852 4102 896 4224
rect 1245 4211 1328 4232
rect 1568 4294 1602 4328
rect 1568 4284 1820 4294
rect 1568 4232 1758 4284
rect 1810 4232 1820 4284
rect 1568 4222 1820 4232
rect 1568 4190 1608 4222
rect 1853 4190 1892 4328
rect 2185 4190 2224 4328
rect 2255 4291 2325 4297
rect 2255 4282 2331 4291
rect 2255 4230 2270 4282
rect 2322 4230 2331 4282
rect 2255 4221 2331 4230
rect 2255 4215 2325 4221
rect 2368 4190 2407 4328
rect 2530 4294 2574 4328
rect 2758 4328 2816 4375
rect 2928 4481 2974 4528
rect 2928 4447 2934 4481
rect 2968 4468 2974 4481
rect 3114 4481 3160 4528
rect 3114 4468 3120 4481
rect 2968 4447 3120 4468
rect 3154 4447 3160 4481
rect 3272 4481 3318 4528
rect 3272 4471 3278 4481
rect 3312 4471 3318 4481
rect 3736 4491 3782 4537
rect 2928 4409 3160 4447
rect 3262 4419 3268 4471
rect 3320 4419 3326 4471
rect 3736 4457 3742 4491
rect 3776 4457 3782 4491
rect 3736 4419 3782 4457
rect 2928 4375 2934 4409
rect 2968 4375 3120 4409
rect 3154 4375 3160 4409
rect 2928 4358 3160 4375
rect 2928 4328 2974 4358
rect 3114 4328 3160 4358
rect 3272 4409 3318 4419
rect 3272 4375 3278 4409
rect 3312 4375 3318 4409
rect 3272 4328 3318 4375
rect 3736 4385 3742 4419
rect 3776 4385 3782 4419
rect 3736 4338 3782 4385
rect 3894 4491 3940 4538
rect 3894 4457 3900 4491
rect 3934 4457 3940 4491
rect 3894 4419 3940 4457
rect 3894 4385 3900 4419
rect 3934 4385 3940 4419
rect 3894 4338 3940 4385
rect 4044 4491 4090 4594
rect 4558 4538 4597 4744
rect 4738 4738 4744 4744
rect 4796 4738 4802 4790
rect 4868 4538 4907 4825
rect 5081 4831 7015 4861
rect 5029 4814 5081 4820
rect 6862 4783 6868 4790
rect 6516 4744 6868 4783
rect 5682 4690 6222 4734
rect 5682 4638 5734 4690
rect 5786 4680 5798 4690
rect 5850 4680 5862 4690
rect 5914 4680 5926 4690
rect 5978 4680 5990 4690
rect 6042 4680 6054 4690
rect 6106 4680 6118 4690
rect 5790 4646 5798 4680
rect 6042 4646 6044 4680
rect 6106 4646 6116 4680
rect 5786 4638 5798 4646
rect 5850 4638 5862 4646
rect 5914 4638 5926 4646
rect 5978 4638 5990 4646
rect 6042 4638 6054 4646
rect 6106 4638 6118 4646
rect 6170 4638 6222 4690
rect 5682 4594 6222 4638
rect 5700 4538 5746 4594
rect 4044 4457 4050 4491
rect 4084 4457 4090 4491
rect 4044 4419 4090 4457
rect 4044 4385 4050 4419
rect 4084 4385 4090 4419
rect 4044 4338 4090 4385
rect 4202 4491 4248 4538
rect 4202 4457 4208 4491
rect 4242 4457 4248 4491
rect 4396 4491 4442 4538
rect 4396 4465 4402 4491
rect 4202 4419 4248 4457
rect 4202 4385 4208 4419
rect 4242 4385 4248 4419
rect 4285 4463 4402 4465
rect 4285 4411 4292 4463
rect 4344 4457 4402 4463
rect 4436 4457 4442 4491
rect 4344 4419 4442 4457
rect 4344 4411 4402 4419
rect 4285 4410 4402 4411
rect 4202 4338 4248 4385
rect 4396 4385 4402 4410
rect 4436 4385 4442 4419
rect 4396 4338 4442 4385
rect 4554 4491 4600 4538
rect 4554 4457 4560 4491
rect 4594 4458 4600 4491
rect 4704 4491 4750 4538
rect 4704 4458 4710 4491
rect 4594 4457 4710 4458
rect 4744 4457 4750 4491
rect 4554 4419 4750 4457
rect 4554 4385 4560 4419
rect 4594 4392 4710 4419
rect 4594 4385 4600 4392
rect 4554 4338 4600 4385
rect 4704 4385 4710 4392
rect 4744 4385 4750 4419
rect 4704 4338 4750 4385
rect 4862 4491 4908 4538
rect 4862 4457 4868 4491
rect 4902 4457 4908 4491
rect 5694 4492 5740 4538
rect 5027 4462 5057 4471
rect 4862 4419 4908 4457
rect 4862 4385 4868 4419
rect 4902 4385 4908 4419
rect 5010 4410 5016 4462
rect 5068 4410 5074 4462
rect 5694 4458 5700 4492
rect 5734 4458 5740 4492
rect 5694 4420 5740 4458
rect 4862 4338 4908 4385
rect 5026 4369 5057 4410
rect 5694 4386 5700 4420
rect 5734 4386 5740 4420
rect 2758 4294 2802 4328
rect 2530 4250 2656 4294
rect 1242 4170 1248 4174
rect 1138 4126 1248 4170
rect 1138 4102 1182 4126
rect 1242 4122 1248 4126
rect 1300 4122 1306 4174
rect 1404 4157 1450 4190
rect 1404 4123 1410 4157
rect 1444 4123 1450 4157
rect 1404 4119 1450 4123
rect 378 4074 434 4080
rect 550 4074 622 4096
rect 434 4068 622 4074
rect 434 4028 565 4068
rect 606 4028 622 4068
rect 434 4018 622 4028
rect 378 4012 434 4018
rect 550 3998 622 4018
rect 696 4068 768 4096
rect 696 4028 712 4068
rect 753 4028 768 4068
rect 696 3998 768 4028
rect 840 4073 912 4102
rect 840 4033 856 4073
rect 897 4033 912 4073
rect 840 4004 912 4033
rect 994 4074 1182 4102
rect 994 4034 1010 4074
rect 1051 4058 1182 4074
rect 1399 4090 1450 4119
rect 1562 4157 1608 4190
rect 1562 4123 1568 4157
rect 1602 4123 1608 4157
rect 1692 4157 1738 4190
rect 1692 4128 1698 4157
rect 1562 4090 1608 4123
rect 1690 4123 1698 4128
rect 1732 4128 1738 4157
rect 1850 4157 1896 4190
rect 2024 4174 2070 4190
rect 1732 4123 1740 4128
rect 1051 4034 1066 4058
rect 1399 4044 1449 4090
rect 1690 4044 1740 4123
rect 1850 4123 1856 4157
rect 1890 4123 1896 4157
rect 1850 4090 1896 4123
rect 2014 4122 2020 4174
rect 2072 4122 2078 4174
rect 2182 4157 2228 4190
rect 2182 4123 2188 4157
rect 2222 4123 2228 4157
rect 2024 4090 2070 4122
rect 2182 4090 2228 4123
rect 2366 4157 2412 4190
rect 2524 4172 2570 4190
rect 2366 4123 2372 4157
rect 2406 4123 2412 4157
rect 2366 4090 2412 4123
rect 2516 4120 2522 4172
rect 2574 4120 2580 4172
rect 2524 4090 2570 4120
rect 2024 4058 2068 4090
rect 2612 4058 2656 4250
rect 994 4004 1066 4034
rect 1324 3989 1960 4044
rect 2024 4014 2656 4058
rect 2694 4250 2802 4294
rect 2832 4280 2904 4290
rect 2694 4052 2738 4250
rect 2832 4228 2842 4280
rect 2894 4228 2904 4280
rect 2832 4218 2904 4228
rect 2933 4190 2972 4328
rect 3118 4190 3157 4328
rect 3272 4284 3316 4328
rect 3268 4278 3320 4284
rect 3555 4253 3561 4305
rect 3613 4298 3619 4305
rect 3662 4298 3713 4310
rect 3613 4295 3713 4298
rect 3613 4261 3670 4295
rect 3704 4261 3713 4295
rect 3613 4259 3713 4261
rect 3613 4253 3619 4259
rect 3662 4247 3713 4259
rect 3897 4289 3936 4338
rect 3976 4296 4027 4301
rect 3970 4289 3976 4296
rect 3897 4250 3976 4289
rect 3268 4220 3320 4226
rect 3897 4200 3936 4250
rect 3970 4244 3976 4250
rect 4028 4244 4034 4296
rect 4206 4282 4245 4338
rect 4300 4282 4347 4293
rect 4206 4280 4347 4282
rect 4206 4247 4306 4280
rect 3976 4238 4027 4244
rect 4206 4200 4245 4247
rect 4300 4246 4306 4247
rect 4340 4246 4347 4280
rect 4300 4234 4347 4246
rect 2766 4184 2818 4190
rect 2766 4126 2776 4132
rect 2770 4123 2776 4126
rect 2810 4126 2818 4132
rect 2928 4157 2974 4190
rect 2810 4123 2816 4126
rect 2770 4090 2816 4123
rect 2928 4123 2934 4157
rect 2968 4123 2974 4157
rect 2928 4090 2974 4123
rect 3114 4157 3160 4190
rect 3114 4123 3120 4157
rect 3154 4123 3160 4157
rect 3114 4090 3160 4123
rect 3272 4157 3318 4190
rect 3272 4123 3278 4157
rect 3312 4123 3318 4157
rect 3272 4090 3318 4123
rect 3274 4052 3318 4090
rect 2694 4008 3318 4052
rect 3736 4167 3782 4200
rect 3736 4133 3742 4167
rect 3776 4133 3782 4167
rect 3736 4100 3782 4133
rect 3894 4167 3940 4200
rect 3894 4133 3900 4167
rect 3934 4133 3940 4167
rect 4044 4167 4090 4200
rect 4044 4138 4050 4167
rect 3894 4100 3940 4133
rect 4042 4133 4050 4138
rect 4084 4133 4090 4167
rect 4042 4100 4090 4133
rect 4202 4167 4248 4200
rect 4202 4133 4208 4167
rect 4242 4133 4248 4167
rect 4202 4100 4248 4133
rect 3736 4044 3780 4100
rect 4042 4044 4089 4100
rect 1324 3937 1360 3989
rect 1412 3937 1424 3989
rect 1476 3980 1488 3989
rect 1540 3980 1552 3989
rect 1604 3980 1616 3989
rect 1668 3980 1680 3989
rect 1732 3980 1744 3989
rect 1796 3980 1808 3989
rect 1479 3946 1488 3980
rect 1551 3946 1552 3980
rect 1732 3946 1733 3980
rect 1796 3946 1805 3980
rect 1476 3937 1488 3946
rect 1540 3937 1552 3946
rect 1604 3937 1616 3946
rect 1668 3937 1680 3946
rect 1732 3937 1744 3946
rect 1796 3937 1808 3946
rect 1860 3937 1872 3989
rect 1924 3937 1960 3989
rect 3704 4000 4244 4044
rect 3704 3991 3756 4000
rect 3808 3991 3820 4000
rect 1324 3904 1960 3937
rect 2346 3959 2426 3984
rect 2346 3955 3517 3959
rect 2346 3921 2369 3955
rect 2403 3921 3517 3955
rect 2346 3917 3517 3921
rect 2346 3892 2426 3917
rect 2636 3859 2702 3871
rect 272 3805 278 3859
rect 332 3805 2642 3859
rect 2696 3805 2702 3859
rect 2636 3793 2702 3805
rect 3475 3764 3517 3917
rect 3704 3957 3741 3991
rect 3808 3957 3813 3991
rect 3704 3948 3756 3957
rect 3808 3948 3820 3957
rect 3872 3948 3884 4000
rect 3936 3948 3948 4000
rect 4000 3948 4012 4000
rect 4064 3948 4076 4000
rect 4128 3991 4140 4000
rect 4192 3991 4244 4000
rect 4135 3957 4140 3991
rect 4207 3957 4244 3991
rect 4128 3948 4140 3957
rect 4192 3948 4244 3957
rect 3704 3904 4244 3948
rect 3559 3799 3565 3851
rect 3617 3844 3623 3851
rect 4306 3844 4345 4234
rect 4558 4202 4597 4338
rect 4628 4307 4680 4313
rect 4625 4258 4628 4304
rect 4680 4258 4683 4304
rect 4875 4262 4904 4338
rect 4628 4249 4680 4255
rect 4875 4234 4980 4262
rect 4396 4169 4442 4202
rect 4396 4135 4402 4169
rect 4436 4135 4442 4169
rect 4396 4102 4442 4135
rect 4554 4182 4600 4202
rect 4704 4182 4750 4202
rect 4862 4182 4908 4202
rect 4554 4169 4750 4182
rect 4554 4135 4560 4169
rect 4594 4135 4710 4169
rect 4744 4135 4750 4169
rect 4554 4116 4750 4135
rect 4856 4130 4862 4182
rect 4914 4130 4920 4182
rect 4554 4102 4600 4116
rect 4704 4102 4750 4116
rect 4862 4102 4908 4130
rect 4402 3952 4430 4102
rect 4558 4057 4597 4102
rect 4552 4051 4604 4057
rect 4552 3993 4604 3999
rect 4952 3952 4980 4234
rect 5026 4184 5056 4369
rect 5694 4338 5740 4386
rect 5852 4492 5898 4538
rect 5852 4458 5858 4492
rect 5892 4458 5898 4492
rect 5852 4420 5898 4458
rect 5852 4386 5858 4420
rect 5892 4386 5898 4420
rect 5852 4338 5898 4386
rect 6002 4492 6048 4594
rect 6516 4538 6556 4744
rect 6862 4738 6868 4744
rect 6920 4738 6926 4790
rect 6985 4778 7015 4831
rect 6985 4749 7016 4778
rect 6002 4458 6008 4492
rect 6042 4458 6048 4492
rect 6002 4420 6048 4458
rect 6002 4386 6008 4420
rect 6042 4386 6048 4420
rect 6002 4338 6048 4386
rect 6160 4492 6206 4538
rect 6160 4458 6166 4492
rect 6200 4458 6206 4492
rect 6354 4492 6400 4538
rect 6354 4466 6360 4492
rect 6160 4420 6206 4458
rect 6160 4386 6166 4420
rect 6200 4386 6206 4420
rect 6244 4464 6360 4466
rect 6244 4412 6250 4464
rect 6302 4458 6360 4464
rect 6394 4458 6400 4492
rect 6302 4420 6400 4458
rect 6302 4412 6360 4420
rect 6244 4410 6360 4412
rect 6160 4338 6206 4386
rect 6354 4386 6360 4410
rect 6394 4386 6400 4420
rect 6354 4338 6400 4386
rect 6512 4492 6558 4538
rect 6512 4458 6518 4492
rect 6552 4458 6558 4492
rect 6662 4492 6708 4538
rect 6662 4458 6668 4492
rect 6702 4458 6708 4492
rect 6512 4420 6708 4458
rect 6512 4386 6518 4420
rect 6552 4392 6668 4420
rect 6552 4386 6558 4392
rect 6512 4338 6558 4386
rect 6662 4386 6668 4392
rect 6702 4386 6708 4420
rect 6662 4338 6708 4386
rect 6820 4492 6866 4538
rect 6820 4458 6826 4492
rect 6860 4458 6866 4492
rect 6986 4462 7016 4749
rect 7206 4678 7234 4936
rect 7194 4672 7246 4678
rect 7194 4614 7246 4620
rect 6820 4420 6866 4458
rect 6820 4386 6826 4420
rect 6860 4386 6866 4420
rect 6968 4410 6974 4462
rect 7026 4410 7032 4462
rect 6820 4338 6866 4386
rect 6984 4370 7016 4410
rect 5111 4253 5117 4305
rect 5169 4298 5175 4305
rect 5620 4298 5672 4310
rect 5169 4296 5672 4298
rect 5169 4262 5628 4296
rect 5662 4262 5672 4296
rect 5169 4259 5672 4262
rect 5169 4253 5175 4259
rect 5620 4248 5672 4259
rect 5856 4290 5894 4338
rect 5934 4296 5986 4302
rect 5928 4290 5934 4296
rect 5856 4250 5934 4290
rect 5856 4200 5894 4250
rect 5928 4244 5934 4250
rect 5986 4244 5992 4296
rect 6164 4282 6204 4338
rect 6258 4282 6306 4294
rect 6164 4280 6306 4282
rect 6164 4248 6264 4280
rect 5934 4238 5986 4244
rect 6164 4200 6204 4248
rect 6258 4246 6264 4248
rect 6298 4246 6306 4280
rect 6258 4234 6306 4246
rect 5009 4132 5015 4184
rect 5067 4132 5073 4184
rect 5694 4168 5740 4200
rect 5694 4134 5700 4168
rect 5734 4134 5740 4168
rect 4402 3924 4980 3952
rect 3617 3805 4345 3844
rect 3617 3799 3623 3805
rect 5021 3764 5063 4132
rect 5694 4100 5740 4134
rect 5852 4168 5898 4200
rect 5852 4134 5858 4168
rect 5892 4134 5898 4168
rect 6002 4168 6048 4200
rect 6002 4138 6008 4168
rect 5852 4100 5898 4134
rect 6000 4134 6008 4138
rect 6042 4134 6048 4168
rect 5694 4044 5738 4100
rect 6000 4044 6048 4134
rect 6160 4168 6206 4200
rect 6160 4134 6166 4168
rect 6200 4134 6206 4168
rect 6160 4100 6206 4134
rect 5662 4000 6202 4044
rect 5662 3992 5714 4000
rect 5766 3992 5778 4000
rect 5662 3958 5700 3992
rect 5766 3958 5772 3992
rect 5662 3948 5714 3958
rect 5766 3948 5778 3958
rect 5830 3948 5842 4000
rect 5894 3948 5906 4000
rect 5958 3948 5970 4000
rect 6022 3948 6034 4000
rect 6086 3992 6098 4000
rect 6150 3992 6202 4000
rect 6094 3958 6098 3992
rect 6166 3958 6202 3992
rect 6086 3948 6098 3958
rect 6150 3948 6202 3958
rect 5662 3904 6202 3948
rect 5111 3799 5117 3851
rect 5169 3844 5175 3851
rect 6264 3844 6304 4234
rect 6516 4202 6556 4338
rect 6586 4308 6638 4314
rect 6584 4258 6586 4304
rect 6638 4258 6642 4304
rect 6834 4262 6862 4338
rect 6586 4250 6638 4256
rect 6834 4234 6936 4262
rect 6354 4170 6400 4202
rect 6354 4136 6360 4170
rect 6394 4136 6400 4170
rect 6354 4102 6400 4136
rect 6512 4182 6558 4202
rect 6662 4182 6708 4202
rect 6820 4182 6866 4202
rect 6512 4170 6708 4182
rect 6512 4136 6518 4170
rect 6552 4136 6668 4170
rect 6702 4136 6708 4170
rect 6512 4116 6708 4136
rect 6814 4130 6820 4182
rect 6872 4130 6878 4182
rect 6512 4102 6558 4116
rect 6662 4102 6708 4116
rect 6820 4102 6866 4130
rect 6360 3952 6388 4102
rect 6516 4058 6556 4102
rect 6510 4052 6562 4058
rect 6510 3994 6562 4000
rect 6908 3952 6936 4234
rect 6984 4184 7014 4370
rect 6968 4132 6974 4184
rect 7026 4132 7032 4184
rect 6360 3924 6936 3952
rect 6908 3860 6936 3924
rect 5169 3806 6304 3844
rect 6346 3832 6936 3860
rect 5169 3805 5572 3806
rect 5169 3799 5175 3805
rect 3475 3722 5063 3764
rect 5035 3681 5087 3687
rect 3472 3597 4907 3636
rect 6346 3669 6374 3832
rect 6908 3830 6936 3832
rect 6512 3766 6564 3772
rect 6512 3708 6564 3714
rect 5087 3641 6374 3669
rect 6523 3651 6553 3708
rect 5035 3623 5087 3629
rect 6523 3621 7015 3651
rect 1348 3463 1880 3506
rect 1348 3454 1398 3463
rect 1450 3454 1462 3463
rect 1348 3420 1383 3454
rect 1450 3420 1455 3454
rect 1348 3411 1398 3420
rect 1450 3411 1462 3420
rect 1514 3411 1526 3463
rect 1578 3411 1590 3463
rect 1642 3411 1654 3463
rect 1706 3411 1718 3463
rect 1770 3454 1782 3463
rect 1834 3454 1880 3463
rect 1777 3420 1782 3454
rect 1849 3420 1880 3454
rect 3472 3439 3511 3597
rect 4738 3555 4744 3562
rect 4558 3516 4744 3555
rect 1770 3411 1782 3420
rect 1834 3411 1880 3420
rect 550 3392 622 3396
rect 550 3340 560 3392
rect 612 3340 622 3392
rect 696 3390 768 3396
rect 550 3328 566 3340
rect 607 3328 622 3340
rect 682 3388 768 3390
rect 682 3336 702 3388
rect 754 3336 768 3388
rect 682 3334 710 3336
rect 550 3298 622 3328
rect 696 3328 710 3334
rect 751 3328 768 3336
rect 696 3298 768 3328
rect 840 3373 912 3402
rect 840 3333 856 3373
rect 897 3333 912 3373
rect 840 3304 912 3333
rect 994 3373 1066 3402
rect 994 3333 1009 3373
rect 1050 3333 1066 3373
rect 1348 3366 1880 3411
rect 994 3304 1066 3333
rect 564 3258 608 3298
rect 856 3238 900 3304
rect 378 3230 433 3236
rect 846 3186 852 3238
rect 904 3186 910 3238
rect 378 2945 433 3175
rect 856 3146 900 3186
rect 1008 3146 1052 3304
rect 1407 3300 1448 3366
rect 1693 3300 1735 3366
rect 1941 3363 2687 3408
rect 1404 3253 1450 3300
rect 1404 3219 1410 3253
rect 1444 3219 1450 3253
rect 1404 3181 1450 3219
rect 1404 3147 1410 3181
rect 1444 3147 1450 3181
rect 708 3102 900 3146
rect 372 2890 378 2945
rect 433 2890 439 2945
rect 708 2868 752 3102
rect 998 3094 1004 3146
rect 1056 3094 1062 3146
rect 1404 3100 1450 3147
rect 1562 3253 1608 3300
rect 1562 3219 1568 3253
rect 1602 3219 1608 3253
rect 1562 3181 1608 3219
rect 1562 3147 1568 3181
rect 1602 3147 1608 3181
rect 1562 3100 1608 3147
rect 1692 3253 1738 3300
rect 1692 3219 1698 3253
rect 1732 3219 1738 3253
rect 1692 3181 1738 3219
rect 1692 3147 1698 3181
rect 1732 3147 1738 3181
rect 1692 3100 1738 3147
rect 1850 3297 1896 3300
rect 1941 3297 1986 3363
rect 1850 3253 1986 3297
rect 1850 3219 1856 3253
rect 1890 3252 1986 3253
rect 2024 3253 2070 3300
rect 1890 3219 1896 3252
rect 1850 3181 1896 3219
rect 2024 3219 2030 3253
rect 2064 3219 2070 3253
rect 2024 3184 2070 3219
rect 1998 3182 2070 3184
rect 1850 3147 1856 3181
rect 1890 3147 1896 3181
rect 1850 3100 1896 3147
rect 1928 3181 2070 3182
rect 1928 3157 2030 3181
rect 1928 3140 1935 3157
rect 1929 3105 1935 3140
rect 1987 3147 2030 3157
rect 2064 3147 2070 3181
rect 1987 3140 2070 3147
rect 1987 3105 1993 3140
rect 2024 3100 2070 3140
rect 2182 3256 2228 3300
rect 2366 3256 2412 3300
rect 2182 3253 2412 3256
rect 2182 3219 2188 3253
rect 2222 3219 2372 3253
rect 2406 3219 2412 3253
rect 2182 3181 2412 3219
rect 2182 3147 2188 3181
rect 2222 3147 2372 3181
rect 2406 3147 2412 3181
rect 2182 3130 2412 3147
rect 2182 3100 2228 3130
rect 2366 3100 2412 3130
rect 2524 3253 2570 3300
rect 2524 3219 2530 3253
rect 2564 3219 2570 3253
rect 2642 3229 2687 3363
rect 3118 3400 3511 3439
rect 3724 3462 4264 3506
rect 3724 3410 3776 3462
rect 3828 3453 3840 3462
rect 3892 3453 3904 3462
rect 3956 3453 3968 3462
rect 4020 3453 4032 3462
rect 4084 3453 4096 3462
rect 4148 3453 4160 3462
rect 3831 3419 3840 3453
rect 3903 3419 3904 3453
rect 4084 3419 4085 3453
rect 4148 3419 4157 3453
rect 3828 3410 3840 3419
rect 3892 3410 3904 3419
rect 3956 3410 3968 3419
rect 4020 3410 4032 3419
rect 4084 3410 4096 3419
rect 4148 3410 4160 3419
rect 4212 3410 4264 3462
rect 2774 3356 2816 3357
rect 2758 3348 2816 3356
rect 2758 3296 2769 3348
rect 2821 3296 2827 3348
rect 3118 3300 3157 3400
rect 3724 3366 4264 3410
rect 3741 3310 3787 3366
rect 3736 3309 3787 3310
rect 2758 3253 2816 3296
rect 2524 3181 2570 3219
rect 2524 3147 2530 3181
rect 2564 3147 2570 3181
rect 2524 3140 2570 3147
rect 2613 3201 2715 3229
rect 2613 3167 2647 3201
rect 2681 3167 2715 3201
rect 2524 3100 2574 3140
rect 2613 3139 2715 3167
rect 2758 3219 2776 3253
rect 2810 3219 2816 3253
rect 2758 3181 2816 3219
rect 2758 3147 2776 3181
rect 2810 3147 2816 3181
rect 1008 3040 1052 3094
rect 1245 3059 1328 3078
rect 852 2996 1052 3040
rect 1148 3057 1328 3059
rect 1148 3005 1155 3057
rect 1207 3047 1328 3057
rect 1207 3013 1269 3047
rect 1303 3013 1328 3047
rect 1207 3005 1328 3013
rect 1148 3004 1328 3005
rect 852 2874 896 2996
rect 1245 2983 1328 3004
rect 1568 3066 1602 3100
rect 1568 3056 1820 3066
rect 1568 3004 1758 3056
rect 1810 3004 1820 3056
rect 1568 2994 1820 3004
rect 1568 2962 1608 2994
rect 1853 2962 1892 3100
rect 2185 2962 2224 3100
rect 2255 3063 2325 3069
rect 2255 3054 2331 3063
rect 2255 3002 2270 3054
rect 2322 3002 2331 3054
rect 2255 2993 2331 3002
rect 2255 2987 2325 2993
rect 2368 2962 2407 3100
rect 2530 3066 2574 3100
rect 2758 3100 2816 3147
rect 2928 3253 2974 3300
rect 2928 3219 2934 3253
rect 2968 3240 2974 3253
rect 3114 3253 3160 3300
rect 3114 3240 3120 3253
rect 2968 3219 3120 3240
rect 3154 3219 3160 3253
rect 3272 3253 3318 3300
rect 3272 3243 3278 3253
rect 3312 3243 3318 3253
rect 3736 3263 3782 3309
rect 2928 3181 3160 3219
rect 3262 3191 3268 3243
rect 3320 3191 3326 3243
rect 3736 3229 3742 3263
rect 3776 3229 3782 3263
rect 3736 3191 3782 3229
rect 2928 3147 2934 3181
rect 2968 3147 3120 3181
rect 3154 3147 3160 3181
rect 2928 3130 3160 3147
rect 2928 3100 2974 3130
rect 3114 3100 3160 3130
rect 3272 3181 3318 3191
rect 3272 3147 3278 3181
rect 3312 3147 3318 3181
rect 3272 3100 3318 3147
rect 3736 3157 3742 3191
rect 3776 3157 3782 3191
rect 3736 3110 3782 3157
rect 3894 3263 3940 3310
rect 3894 3229 3900 3263
rect 3934 3229 3940 3263
rect 3894 3191 3940 3229
rect 3894 3157 3900 3191
rect 3934 3157 3940 3191
rect 3894 3110 3940 3157
rect 4044 3263 4090 3366
rect 4558 3310 4597 3516
rect 4738 3510 4744 3516
rect 4796 3510 4802 3562
rect 4868 3310 4907 3597
rect 6837 3555 6843 3562
rect 6516 3516 6843 3555
rect 5682 3462 6222 3506
rect 5682 3410 5734 3462
rect 5786 3452 5798 3462
rect 5850 3452 5862 3462
rect 5914 3452 5926 3462
rect 5978 3452 5990 3462
rect 6042 3452 6054 3462
rect 6106 3452 6118 3462
rect 5790 3418 5798 3452
rect 6042 3418 6044 3452
rect 6106 3418 6116 3452
rect 5786 3410 5798 3418
rect 5850 3410 5862 3418
rect 5914 3410 5926 3418
rect 5978 3410 5990 3418
rect 6042 3410 6054 3418
rect 6106 3410 6118 3418
rect 6170 3410 6222 3462
rect 5682 3366 6222 3410
rect 5700 3310 5746 3366
rect 4044 3229 4050 3263
rect 4084 3229 4090 3263
rect 4044 3191 4090 3229
rect 4044 3157 4050 3191
rect 4084 3157 4090 3191
rect 4044 3110 4090 3157
rect 4202 3263 4248 3310
rect 4202 3229 4208 3263
rect 4242 3229 4248 3263
rect 4396 3263 4442 3310
rect 4396 3237 4402 3263
rect 4202 3191 4248 3229
rect 4202 3157 4208 3191
rect 4242 3157 4248 3191
rect 4285 3235 4402 3237
rect 4285 3183 4292 3235
rect 4344 3229 4402 3235
rect 4436 3229 4442 3263
rect 4344 3191 4442 3229
rect 4344 3183 4402 3191
rect 4285 3182 4402 3183
rect 4202 3110 4248 3157
rect 4396 3157 4402 3182
rect 4436 3157 4442 3191
rect 4396 3110 4442 3157
rect 4554 3263 4600 3310
rect 4554 3229 4560 3263
rect 4594 3230 4600 3263
rect 4704 3263 4750 3310
rect 4704 3230 4710 3263
rect 4594 3229 4710 3230
rect 4744 3229 4750 3263
rect 4554 3191 4750 3229
rect 4554 3157 4560 3191
rect 4594 3164 4710 3191
rect 4594 3157 4600 3164
rect 4554 3110 4600 3157
rect 4704 3157 4710 3164
rect 4744 3157 4750 3191
rect 4704 3110 4750 3157
rect 4862 3263 4908 3310
rect 4862 3229 4868 3263
rect 4902 3229 4908 3263
rect 5694 3264 5740 3310
rect 5027 3234 5057 3243
rect 4862 3191 4908 3229
rect 4862 3157 4868 3191
rect 4902 3157 4908 3191
rect 5010 3182 5016 3234
rect 5068 3182 5074 3234
rect 5694 3230 5700 3264
rect 5734 3230 5740 3264
rect 5694 3192 5740 3230
rect 4862 3110 4908 3157
rect 5026 3141 5057 3182
rect 5694 3158 5700 3192
rect 5734 3158 5740 3192
rect 2758 3066 2802 3100
rect 2530 3022 2656 3066
rect 1242 2942 1248 2946
rect 1138 2898 1248 2942
rect 1138 2874 1182 2898
rect 1242 2894 1248 2898
rect 1300 2894 1306 2946
rect 1404 2929 1450 2962
rect 1404 2895 1410 2929
rect 1444 2895 1450 2929
rect 1404 2891 1450 2895
rect 378 2846 434 2852
rect 550 2846 622 2868
rect 434 2840 622 2846
rect 434 2800 565 2840
rect 606 2800 622 2840
rect 434 2790 622 2800
rect 378 2784 434 2790
rect 550 2770 622 2790
rect 696 2840 768 2868
rect 696 2800 712 2840
rect 753 2800 768 2840
rect 696 2770 768 2800
rect 840 2845 912 2874
rect 840 2805 856 2845
rect 897 2805 912 2845
rect 840 2776 912 2805
rect 994 2846 1182 2874
rect 994 2806 1010 2846
rect 1051 2830 1182 2846
rect 1399 2862 1450 2891
rect 1562 2929 1608 2962
rect 1562 2895 1568 2929
rect 1602 2895 1608 2929
rect 1692 2929 1738 2962
rect 1692 2900 1698 2929
rect 1562 2862 1608 2895
rect 1690 2895 1698 2900
rect 1732 2900 1738 2929
rect 1850 2929 1896 2962
rect 2024 2946 2070 2962
rect 1732 2895 1740 2900
rect 1051 2806 1066 2830
rect 1399 2816 1449 2862
rect 1690 2816 1740 2895
rect 1850 2895 1856 2929
rect 1890 2895 1896 2929
rect 1850 2862 1896 2895
rect 2014 2894 2020 2946
rect 2072 2894 2078 2946
rect 2182 2929 2228 2962
rect 2182 2895 2188 2929
rect 2222 2895 2228 2929
rect 2024 2862 2070 2894
rect 2182 2862 2228 2895
rect 2366 2929 2412 2962
rect 2524 2944 2570 2962
rect 2366 2895 2372 2929
rect 2406 2895 2412 2929
rect 2366 2862 2412 2895
rect 2516 2892 2522 2944
rect 2574 2892 2580 2944
rect 2524 2862 2570 2892
rect 2024 2830 2068 2862
rect 2612 2830 2656 3022
rect 994 2776 1066 2806
rect 1324 2761 1960 2816
rect 2024 2786 2656 2830
rect 2694 3022 2802 3066
rect 2832 3052 2904 3062
rect 2694 2824 2738 3022
rect 2832 3000 2842 3052
rect 2894 3000 2904 3052
rect 2832 2990 2904 3000
rect 2933 2962 2972 3100
rect 3118 2962 3157 3100
rect 3272 3056 3316 3100
rect 3268 3050 3320 3056
rect 3555 3025 3561 3077
rect 3613 3070 3619 3077
rect 3662 3070 3713 3082
rect 3613 3067 3713 3070
rect 3613 3033 3670 3067
rect 3704 3033 3713 3067
rect 3613 3031 3713 3033
rect 3613 3025 3619 3031
rect 3662 3019 3713 3031
rect 3897 3061 3936 3110
rect 3976 3068 4027 3073
rect 3970 3061 3976 3068
rect 3897 3022 3976 3061
rect 3268 2992 3320 2998
rect 3897 2972 3936 3022
rect 3970 3016 3976 3022
rect 4028 3016 4034 3068
rect 4206 3054 4245 3110
rect 4300 3054 4347 3065
rect 4206 3052 4347 3054
rect 4206 3019 4306 3052
rect 3976 3010 4027 3016
rect 4206 2972 4245 3019
rect 4300 3018 4306 3019
rect 4340 3018 4347 3052
rect 4300 3006 4347 3018
rect 2766 2956 2818 2962
rect 2766 2898 2776 2904
rect 2770 2895 2776 2898
rect 2810 2898 2818 2904
rect 2928 2929 2974 2962
rect 2810 2895 2816 2898
rect 2770 2862 2816 2895
rect 2928 2895 2934 2929
rect 2968 2895 2974 2929
rect 2928 2862 2974 2895
rect 3114 2929 3160 2962
rect 3114 2895 3120 2929
rect 3154 2895 3160 2929
rect 3114 2862 3160 2895
rect 3272 2929 3318 2962
rect 3272 2895 3278 2929
rect 3312 2895 3318 2929
rect 3272 2862 3318 2895
rect 3274 2824 3318 2862
rect 2694 2780 3318 2824
rect 3736 2939 3782 2972
rect 3736 2905 3742 2939
rect 3776 2905 3782 2939
rect 3736 2872 3782 2905
rect 3894 2939 3940 2972
rect 3894 2905 3900 2939
rect 3934 2905 3940 2939
rect 4044 2939 4090 2972
rect 4044 2910 4050 2939
rect 3894 2872 3940 2905
rect 4042 2905 4050 2910
rect 4084 2905 4090 2939
rect 4042 2872 4090 2905
rect 4202 2939 4248 2972
rect 4202 2905 4208 2939
rect 4242 2905 4248 2939
rect 4202 2872 4248 2905
rect 3736 2816 3780 2872
rect 4042 2816 4089 2872
rect 1324 2709 1360 2761
rect 1412 2709 1424 2761
rect 1476 2752 1488 2761
rect 1540 2752 1552 2761
rect 1604 2752 1616 2761
rect 1668 2752 1680 2761
rect 1732 2752 1744 2761
rect 1796 2752 1808 2761
rect 1479 2718 1488 2752
rect 1551 2718 1552 2752
rect 1732 2718 1733 2752
rect 1796 2718 1805 2752
rect 1476 2709 1488 2718
rect 1540 2709 1552 2718
rect 1604 2709 1616 2718
rect 1668 2709 1680 2718
rect 1732 2709 1744 2718
rect 1796 2709 1808 2718
rect 1860 2709 1872 2761
rect 1924 2709 1960 2761
rect 3704 2772 4244 2816
rect 3704 2763 3756 2772
rect 3808 2763 3820 2772
rect 1324 2676 1960 2709
rect 2346 2731 2426 2756
rect 2346 2727 3517 2731
rect 2346 2693 2369 2727
rect 2403 2693 3517 2727
rect 2346 2689 3517 2693
rect 2346 2664 2426 2689
rect 2636 2631 2702 2643
rect 272 2577 278 2631
rect 332 2577 2642 2631
rect 2696 2577 2702 2631
rect 2636 2565 2702 2577
rect 3475 2536 3517 2689
rect 3704 2729 3741 2763
rect 3808 2729 3813 2763
rect 3704 2720 3756 2729
rect 3808 2720 3820 2729
rect 3872 2720 3884 2772
rect 3936 2720 3948 2772
rect 4000 2720 4012 2772
rect 4064 2720 4076 2772
rect 4128 2763 4140 2772
rect 4192 2763 4244 2772
rect 4135 2729 4140 2763
rect 4207 2729 4244 2763
rect 4128 2720 4140 2729
rect 4192 2720 4244 2729
rect 3704 2676 4244 2720
rect 3559 2571 3565 2623
rect 3617 2616 3623 2623
rect 4306 2616 4345 3006
rect 4558 2974 4597 3110
rect 4628 3079 4680 3085
rect 4625 3030 4628 3076
rect 4680 3030 4683 3076
rect 4875 3034 4904 3110
rect 4628 3021 4680 3027
rect 4875 3006 4980 3034
rect 4396 2941 4442 2974
rect 4396 2907 4402 2941
rect 4436 2907 4442 2941
rect 4396 2874 4442 2907
rect 4554 2954 4600 2974
rect 4704 2954 4750 2974
rect 4862 2954 4908 2974
rect 4554 2941 4750 2954
rect 4554 2907 4560 2941
rect 4594 2907 4710 2941
rect 4744 2907 4750 2941
rect 4554 2888 4750 2907
rect 4856 2902 4862 2954
rect 4914 2902 4920 2954
rect 4554 2874 4600 2888
rect 4704 2874 4750 2888
rect 4862 2874 4908 2902
rect 4402 2724 4430 2874
rect 4558 2829 4597 2874
rect 4552 2823 4604 2829
rect 4552 2765 4604 2771
rect 4952 2724 4980 3006
rect 5026 2956 5056 3141
rect 5694 3110 5740 3158
rect 5852 3264 5898 3310
rect 5852 3230 5858 3264
rect 5892 3230 5898 3264
rect 5852 3192 5898 3230
rect 5852 3158 5858 3192
rect 5892 3158 5898 3192
rect 5852 3110 5898 3158
rect 6002 3264 6048 3366
rect 6516 3310 6556 3516
rect 6837 3510 6843 3516
rect 6895 3510 6901 3562
rect 6985 3550 7015 3621
rect 6985 3521 7016 3550
rect 6002 3230 6008 3264
rect 6042 3230 6048 3264
rect 6002 3192 6048 3230
rect 6002 3158 6008 3192
rect 6042 3158 6048 3192
rect 6002 3110 6048 3158
rect 6160 3264 6206 3310
rect 6160 3230 6166 3264
rect 6200 3230 6206 3264
rect 6354 3264 6400 3310
rect 6354 3238 6360 3264
rect 6160 3192 6206 3230
rect 6160 3158 6166 3192
rect 6200 3158 6206 3192
rect 6244 3236 6360 3238
rect 6244 3184 6250 3236
rect 6302 3230 6360 3236
rect 6394 3230 6400 3264
rect 6302 3192 6400 3230
rect 6302 3184 6360 3192
rect 6244 3182 6360 3184
rect 6160 3110 6206 3158
rect 6354 3158 6360 3182
rect 6394 3158 6400 3192
rect 6354 3110 6400 3158
rect 6512 3264 6558 3310
rect 6512 3230 6518 3264
rect 6552 3230 6558 3264
rect 6662 3264 6708 3310
rect 6662 3230 6668 3264
rect 6702 3230 6708 3264
rect 6512 3192 6708 3230
rect 6512 3158 6518 3192
rect 6552 3164 6668 3192
rect 6552 3158 6558 3164
rect 6512 3110 6558 3158
rect 6662 3158 6668 3164
rect 6702 3158 6708 3192
rect 6662 3110 6708 3158
rect 6820 3264 6866 3310
rect 6820 3230 6826 3264
rect 6860 3230 6866 3264
rect 6986 3234 7016 3521
rect 6820 3192 6866 3230
rect 6820 3158 6826 3192
rect 6860 3158 6866 3192
rect 6968 3182 6974 3234
rect 7026 3182 7032 3234
rect 6820 3110 6866 3158
rect 6984 3142 7016 3182
rect 5191 3025 5197 3077
rect 5249 3070 5255 3077
rect 5620 3070 5672 3082
rect 5249 3068 5672 3070
rect 5249 3034 5628 3068
rect 5662 3034 5672 3068
rect 5249 3031 5672 3034
rect 5249 3025 5255 3031
rect 5620 3020 5672 3031
rect 5856 3062 5894 3110
rect 5934 3068 5986 3074
rect 5928 3062 5934 3068
rect 5856 3022 5934 3062
rect 5856 2972 5894 3022
rect 5928 3016 5934 3022
rect 5986 3016 5992 3068
rect 6164 3054 6204 3110
rect 6258 3054 6306 3066
rect 6164 3052 6306 3054
rect 6164 3020 6264 3052
rect 5934 3010 5986 3016
rect 6164 2972 6204 3020
rect 6258 3018 6264 3020
rect 6298 3018 6306 3052
rect 6258 3006 6306 3018
rect 5009 2904 5015 2956
rect 5067 2904 5073 2956
rect 5694 2940 5740 2972
rect 5694 2906 5700 2940
rect 5734 2906 5740 2940
rect 4402 2696 4980 2724
rect 3617 2577 4345 2616
rect 3617 2571 3623 2577
rect 5021 2536 5063 2904
rect 5694 2872 5740 2906
rect 5852 2940 5898 2972
rect 5852 2906 5858 2940
rect 5892 2906 5898 2940
rect 6002 2940 6048 2972
rect 6002 2910 6008 2940
rect 5852 2872 5898 2906
rect 6000 2906 6008 2910
rect 6042 2906 6048 2940
rect 5694 2816 5738 2872
rect 6000 2816 6048 2906
rect 6160 2940 6206 2972
rect 6160 2906 6166 2940
rect 6200 2906 6206 2940
rect 6160 2872 6206 2906
rect 5662 2772 6202 2816
rect 5662 2764 5714 2772
rect 5766 2764 5778 2772
rect 5662 2730 5700 2764
rect 5766 2730 5772 2764
rect 5662 2720 5714 2730
rect 5766 2720 5778 2730
rect 5830 2720 5842 2772
rect 5894 2720 5906 2772
rect 5958 2720 5970 2772
rect 6022 2720 6034 2772
rect 6086 2764 6098 2772
rect 6150 2764 6202 2772
rect 6094 2730 6098 2764
rect 6166 2730 6202 2764
rect 6086 2720 6098 2730
rect 6150 2720 6202 2730
rect 5662 2676 6202 2720
rect 5191 2571 5197 2623
rect 5249 2616 5255 2623
rect 6264 2616 6304 3006
rect 6516 2974 6556 3110
rect 6586 3080 6638 3086
rect 6584 3030 6586 3076
rect 6638 3030 6642 3076
rect 6834 3034 6862 3110
rect 6586 3022 6638 3028
rect 6834 3006 6936 3034
rect 6354 2942 6400 2974
rect 6354 2908 6360 2942
rect 6394 2908 6400 2942
rect 6354 2874 6400 2908
rect 6512 2954 6558 2974
rect 6662 2954 6708 2974
rect 6820 2954 6866 2974
rect 6512 2942 6708 2954
rect 6512 2908 6518 2942
rect 6552 2908 6668 2942
rect 6702 2908 6708 2942
rect 6512 2888 6708 2908
rect 6814 2902 6820 2954
rect 6872 2902 6878 2954
rect 6512 2874 6558 2888
rect 6662 2874 6708 2888
rect 6820 2874 6866 2902
rect 6360 2724 6388 2874
rect 6516 2830 6556 2874
rect 6510 2824 6562 2830
rect 6510 2766 6562 2772
rect 6908 2724 6936 3006
rect 6984 2956 7014 3142
rect 6968 2904 6974 2956
rect 7026 2904 7032 2956
rect 6360 2696 6936 2724
rect 5249 2578 6304 2616
rect 5249 2577 5587 2578
rect 5249 2571 5255 2577
rect 3475 2494 5063 2536
rect 6908 2524 6936 2696
rect 7107 2536 7159 2542
rect 6908 2496 7107 2524
rect 7107 2478 7159 2484
rect 5029 2416 5081 2422
rect 3472 2369 4907 2408
rect 1348 2235 1880 2278
rect 1348 2226 1398 2235
rect 1450 2226 1462 2235
rect 1348 2192 1383 2226
rect 1450 2192 1455 2226
rect 1348 2183 1398 2192
rect 1450 2183 1462 2192
rect 1514 2183 1526 2235
rect 1578 2183 1590 2235
rect 1642 2183 1654 2235
rect 1706 2183 1718 2235
rect 1770 2226 1782 2235
rect 1834 2226 1880 2235
rect 1777 2192 1782 2226
rect 1849 2192 1880 2226
rect 3472 2211 3511 2369
rect 4738 2327 4744 2334
rect 4558 2288 4744 2327
rect 1770 2183 1782 2192
rect 1834 2183 1880 2192
rect 550 2164 622 2168
rect 550 2112 560 2164
rect 612 2112 622 2164
rect 696 2162 768 2168
rect 550 2100 566 2112
rect 607 2100 622 2112
rect 682 2160 768 2162
rect 682 2108 702 2160
rect 754 2108 768 2160
rect 682 2106 710 2108
rect 550 2070 622 2100
rect 696 2100 710 2106
rect 751 2100 768 2108
rect 696 2070 768 2100
rect 840 2145 912 2174
rect 840 2105 856 2145
rect 897 2105 912 2145
rect 840 2076 912 2105
rect 994 2145 1066 2174
rect 994 2105 1009 2145
rect 1050 2105 1066 2145
rect 1348 2138 1880 2183
rect 994 2076 1066 2105
rect 564 2030 608 2070
rect 856 2010 900 2076
rect 378 2002 433 2008
rect 846 1958 852 2010
rect 904 1958 910 2010
rect 378 1717 433 1947
rect 856 1918 900 1958
rect 1008 1918 1052 2076
rect 1407 2072 1448 2138
rect 1693 2072 1735 2138
rect 1941 2135 2687 2180
rect 1404 2025 1450 2072
rect 1404 1991 1410 2025
rect 1444 1991 1450 2025
rect 1404 1953 1450 1991
rect 1404 1919 1410 1953
rect 1444 1919 1450 1953
rect 708 1874 900 1918
rect 372 1662 378 1717
rect 433 1662 439 1717
rect 708 1640 752 1874
rect 998 1866 1004 1918
rect 1056 1866 1062 1918
rect 1404 1872 1450 1919
rect 1562 2025 1608 2072
rect 1562 1991 1568 2025
rect 1602 1991 1608 2025
rect 1562 1953 1608 1991
rect 1562 1919 1568 1953
rect 1602 1919 1608 1953
rect 1562 1872 1608 1919
rect 1692 2025 1738 2072
rect 1692 1991 1698 2025
rect 1732 1991 1738 2025
rect 1692 1953 1738 1991
rect 1692 1919 1698 1953
rect 1732 1919 1738 1953
rect 1692 1872 1738 1919
rect 1850 2069 1896 2072
rect 1941 2069 1986 2135
rect 1850 2025 1986 2069
rect 1850 1991 1856 2025
rect 1890 2024 1986 2025
rect 2024 2025 2070 2072
rect 1890 1991 1896 2024
rect 1850 1953 1896 1991
rect 2024 1991 2030 2025
rect 2064 1991 2070 2025
rect 2024 1956 2070 1991
rect 1998 1954 2070 1956
rect 1850 1919 1856 1953
rect 1890 1919 1896 1953
rect 1850 1872 1896 1919
rect 1928 1953 2070 1954
rect 1928 1929 2030 1953
rect 1928 1912 1935 1929
rect 1929 1877 1935 1912
rect 1987 1919 2030 1929
rect 2064 1919 2070 1953
rect 1987 1912 2070 1919
rect 1987 1877 1993 1912
rect 2024 1872 2070 1912
rect 2182 2028 2228 2072
rect 2366 2028 2412 2072
rect 2182 2025 2412 2028
rect 2182 1991 2188 2025
rect 2222 1991 2372 2025
rect 2406 1991 2412 2025
rect 2182 1953 2412 1991
rect 2182 1919 2188 1953
rect 2222 1919 2372 1953
rect 2406 1919 2412 1953
rect 2182 1902 2412 1919
rect 2182 1872 2228 1902
rect 2366 1872 2412 1902
rect 2524 2025 2570 2072
rect 2524 1991 2530 2025
rect 2564 1991 2570 2025
rect 2642 2001 2687 2135
rect 3118 2172 3511 2211
rect 3724 2234 4264 2278
rect 3724 2182 3776 2234
rect 3828 2225 3840 2234
rect 3892 2225 3904 2234
rect 3956 2225 3968 2234
rect 4020 2225 4032 2234
rect 4084 2225 4096 2234
rect 4148 2225 4160 2234
rect 3831 2191 3840 2225
rect 3903 2191 3904 2225
rect 4084 2191 4085 2225
rect 4148 2191 4157 2225
rect 3828 2182 3840 2191
rect 3892 2182 3904 2191
rect 3956 2182 3968 2191
rect 4020 2182 4032 2191
rect 4084 2182 4096 2191
rect 4148 2182 4160 2191
rect 4212 2182 4264 2234
rect 2774 2128 2816 2129
rect 2758 2120 2816 2128
rect 2758 2068 2769 2120
rect 2821 2068 2827 2120
rect 3118 2072 3157 2172
rect 3724 2138 4264 2182
rect 3741 2082 3787 2138
rect 3736 2081 3787 2082
rect 2758 2025 2816 2068
rect 2524 1953 2570 1991
rect 2524 1919 2530 1953
rect 2564 1919 2570 1953
rect 2524 1912 2570 1919
rect 2613 1973 2715 2001
rect 2613 1939 2647 1973
rect 2681 1939 2715 1973
rect 2524 1872 2574 1912
rect 2613 1911 2715 1939
rect 2758 1991 2776 2025
rect 2810 1991 2816 2025
rect 2758 1953 2816 1991
rect 2758 1919 2776 1953
rect 2810 1919 2816 1953
rect 1008 1812 1052 1866
rect 1245 1831 1328 1850
rect 852 1768 1052 1812
rect 1148 1829 1328 1831
rect 1148 1777 1155 1829
rect 1207 1819 1328 1829
rect 1207 1785 1269 1819
rect 1303 1785 1328 1819
rect 1207 1777 1328 1785
rect 1148 1776 1328 1777
rect 852 1646 896 1768
rect 1245 1755 1328 1776
rect 1568 1838 1602 1872
rect 1568 1828 1820 1838
rect 1568 1776 1758 1828
rect 1810 1776 1820 1828
rect 1568 1766 1820 1776
rect 1568 1734 1608 1766
rect 1853 1734 1892 1872
rect 2185 1734 2224 1872
rect 2255 1835 2325 1841
rect 2255 1826 2331 1835
rect 2255 1774 2270 1826
rect 2322 1774 2331 1826
rect 2255 1765 2331 1774
rect 2255 1759 2325 1765
rect 2368 1734 2407 1872
rect 2530 1838 2574 1872
rect 2758 1872 2816 1919
rect 2928 2025 2974 2072
rect 2928 1991 2934 2025
rect 2968 2012 2974 2025
rect 3114 2025 3160 2072
rect 3114 2012 3120 2025
rect 2968 1991 3120 2012
rect 3154 1991 3160 2025
rect 3272 2025 3318 2072
rect 3272 2015 3278 2025
rect 3312 2015 3318 2025
rect 3736 2035 3782 2081
rect 2928 1953 3160 1991
rect 3262 1963 3268 2015
rect 3320 1963 3326 2015
rect 3736 2001 3742 2035
rect 3776 2001 3782 2035
rect 3736 1963 3782 2001
rect 2928 1919 2934 1953
rect 2968 1919 3120 1953
rect 3154 1919 3160 1953
rect 2928 1902 3160 1919
rect 2928 1872 2974 1902
rect 3114 1872 3160 1902
rect 3272 1953 3318 1963
rect 3272 1919 3278 1953
rect 3312 1919 3318 1953
rect 3272 1872 3318 1919
rect 3736 1929 3742 1963
rect 3776 1929 3782 1963
rect 3736 1882 3782 1929
rect 3894 2035 3940 2082
rect 3894 2001 3900 2035
rect 3934 2001 3940 2035
rect 3894 1963 3940 2001
rect 3894 1929 3900 1963
rect 3934 1929 3940 1963
rect 3894 1882 3940 1929
rect 4044 2035 4090 2138
rect 4558 2082 4597 2288
rect 4738 2282 4744 2288
rect 4796 2282 4802 2334
rect 4868 2082 4907 2369
rect 5081 2375 7015 2405
rect 5029 2358 5081 2364
rect 6862 2327 6868 2334
rect 6516 2288 6868 2327
rect 5682 2234 6222 2278
rect 5682 2182 5734 2234
rect 5786 2224 5798 2234
rect 5850 2224 5862 2234
rect 5914 2224 5926 2234
rect 5978 2224 5990 2234
rect 6042 2224 6054 2234
rect 6106 2224 6118 2234
rect 5790 2190 5798 2224
rect 6042 2190 6044 2224
rect 6106 2190 6116 2224
rect 5786 2182 5798 2190
rect 5850 2182 5862 2190
rect 5914 2182 5926 2190
rect 5978 2182 5990 2190
rect 6042 2182 6054 2190
rect 6106 2182 6118 2190
rect 6170 2182 6222 2234
rect 5682 2138 6222 2182
rect 5700 2082 5746 2138
rect 4044 2001 4050 2035
rect 4084 2001 4090 2035
rect 4044 1963 4090 2001
rect 4044 1929 4050 1963
rect 4084 1929 4090 1963
rect 4044 1882 4090 1929
rect 4202 2035 4248 2082
rect 4202 2001 4208 2035
rect 4242 2001 4248 2035
rect 4396 2035 4442 2082
rect 4396 2009 4402 2035
rect 4202 1963 4248 2001
rect 4202 1929 4208 1963
rect 4242 1929 4248 1963
rect 4285 2007 4402 2009
rect 4285 1955 4292 2007
rect 4344 2001 4402 2007
rect 4436 2001 4442 2035
rect 4344 1963 4442 2001
rect 4344 1955 4402 1963
rect 4285 1954 4402 1955
rect 4202 1882 4248 1929
rect 4396 1929 4402 1954
rect 4436 1929 4442 1963
rect 4396 1882 4442 1929
rect 4554 2035 4600 2082
rect 4554 2001 4560 2035
rect 4594 2002 4600 2035
rect 4704 2035 4750 2082
rect 4704 2002 4710 2035
rect 4594 2001 4710 2002
rect 4744 2001 4750 2035
rect 4554 1963 4750 2001
rect 4554 1929 4560 1963
rect 4594 1936 4710 1963
rect 4594 1929 4600 1936
rect 4554 1882 4600 1929
rect 4704 1929 4710 1936
rect 4744 1929 4750 1963
rect 4704 1882 4750 1929
rect 4862 2035 4908 2082
rect 4862 2001 4868 2035
rect 4902 2001 4908 2035
rect 5694 2036 5740 2082
rect 5027 2006 5057 2015
rect 4862 1963 4908 2001
rect 4862 1929 4868 1963
rect 4902 1929 4908 1963
rect 5010 1954 5016 2006
rect 5068 1954 5074 2006
rect 5694 2002 5700 2036
rect 5734 2002 5740 2036
rect 5694 1964 5740 2002
rect 4862 1882 4908 1929
rect 5026 1913 5057 1954
rect 5694 1930 5700 1964
rect 5734 1930 5740 1964
rect 2758 1838 2802 1872
rect 2530 1794 2656 1838
rect 1242 1714 1248 1718
rect 1138 1670 1248 1714
rect 1138 1646 1182 1670
rect 1242 1666 1248 1670
rect 1300 1666 1306 1718
rect 1404 1701 1450 1734
rect 1404 1667 1410 1701
rect 1444 1667 1450 1701
rect 1404 1663 1450 1667
rect 378 1618 434 1624
rect 550 1618 622 1640
rect 434 1612 622 1618
rect 434 1572 565 1612
rect 606 1572 622 1612
rect 434 1562 622 1572
rect 378 1556 434 1562
rect 550 1542 622 1562
rect 696 1612 768 1640
rect 696 1572 712 1612
rect 753 1572 768 1612
rect 696 1542 768 1572
rect 840 1617 912 1646
rect 840 1577 856 1617
rect 897 1577 912 1617
rect 840 1548 912 1577
rect 994 1618 1182 1646
rect 994 1578 1010 1618
rect 1051 1602 1182 1618
rect 1399 1634 1450 1663
rect 1562 1701 1608 1734
rect 1562 1667 1568 1701
rect 1602 1667 1608 1701
rect 1692 1701 1738 1734
rect 1692 1672 1698 1701
rect 1562 1634 1608 1667
rect 1690 1667 1698 1672
rect 1732 1672 1738 1701
rect 1850 1701 1896 1734
rect 2024 1718 2070 1734
rect 1732 1667 1740 1672
rect 1051 1578 1066 1602
rect 1399 1588 1449 1634
rect 1690 1588 1740 1667
rect 1850 1667 1856 1701
rect 1890 1667 1896 1701
rect 1850 1634 1896 1667
rect 2014 1666 2020 1718
rect 2072 1666 2078 1718
rect 2182 1701 2228 1734
rect 2182 1667 2188 1701
rect 2222 1667 2228 1701
rect 2024 1634 2070 1666
rect 2182 1634 2228 1667
rect 2366 1701 2412 1734
rect 2524 1716 2570 1734
rect 2366 1667 2372 1701
rect 2406 1667 2412 1701
rect 2366 1634 2412 1667
rect 2516 1664 2522 1716
rect 2574 1664 2580 1716
rect 2524 1634 2570 1664
rect 2024 1602 2068 1634
rect 2612 1602 2656 1794
rect 994 1548 1066 1578
rect 1324 1533 1960 1588
rect 2024 1558 2656 1602
rect 2694 1794 2802 1838
rect 2832 1824 2904 1834
rect 2694 1596 2738 1794
rect 2832 1772 2842 1824
rect 2894 1772 2904 1824
rect 2832 1762 2904 1772
rect 2933 1734 2972 1872
rect 3118 1734 3157 1872
rect 3272 1828 3316 1872
rect 3268 1822 3320 1828
rect 3555 1797 3561 1849
rect 3613 1842 3619 1849
rect 3662 1842 3713 1854
rect 3613 1839 3713 1842
rect 3613 1805 3670 1839
rect 3704 1805 3713 1839
rect 3613 1803 3713 1805
rect 3613 1797 3619 1803
rect 3662 1791 3713 1803
rect 3897 1833 3936 1882
rect 3976 1840 4027 1845
rect 3970 1833 3976 1840
rect 3897 1794 3976 1833
rect 3268 1764 3320 1770
rect 3897 1744 3936 1794
rect 3970 1788 3976 1794
rect 4028 1788 4034 1840
rect 4206 1826 4245 1882
rect 4300 1826 4347 1837
rect 4206 1824 4347 1826
rect 4206 1791 4306 1824
rect 3976 1782 4027 1788
rect 4206 1744 4245 1791
rect 4300 1790 4306 1791
rect 4340 1790 4347 1824
rect 4300 1778 4347 1790
rect 2766 1728 2818 1734
rect 2766 1670 2776 1676
rect 2770 1667 2776 1670
rect 2810 1670 2818 1676
rect 2928 1701 2974 1734
rect 2810 1667 2816 1670
rect 2770 1634 2816 1667
rect 2928 1667 2934 1701
rect 2968 1667 2974 1701
rect 2928 1634 2974 1667
rect 3114 1701 3160 1734
rect 3114 1667 3120 1701
rect 3154 1667 3160 1701
rect 3114 1634 3160 1667
rect 3272 1701 3318 1734
rect 3272 1667 3278 1701
rect 3312 1667 3318 1701
rect 3272 1634 3318 1667
rect 3274 1596 3318 1634
rect 2694 1552 3318 1596
rect 3736 1711 3782 1744
rect 3736 1677 3742 1711
rect 3776 1677 3782 1711
rect 3736 1644 3782 1677
rect 3894 1711 3940 1744
rect 3894 1677 3900 1711
rect 3934 1677 3940 1711
rect 4044 1711 4090 1744
rect 4044 1682 4050 1711
rect 3894 1644 3940 1677
rect 4042 1677 4050 1682
rect 4084 1677 4090 1711
rect 4042 1644 4090 1677
rect 4202 1711 4248 1744
rect 4202 1677 4208 1711
rect 4242 1677 4248 1711
rect 4202 1644 4248 1677
rect 3736 1588 3780 1644
rect 4042 1588 4089 1644
rect 1324 1481 1360 1533
rect 1412 1481 1424 1533
rect 1476 1524 1488 1533
rect 1540 1524 1552 1533
rect 1604 1524 1616 1533
rect 1668 1524 1680 1533
rect 1732 1524 1744 1533
rect 1796 1524 1808 1533
rect 1479 1490 1488 1524
rect 1551 1490 1552 1524
rect 1732 1490 1733 1524
rect 1796 1490 1805 1524
rect 1476 1481 1488 1490
rect 1540 1481 1552 1490
rect 1604 1481 1616 1490
rect 1668 1481 1680 1490
rect 1732 1481 1744 1490
rect 1796 1481 1808 1490
rect 1860 1481 1872 1533
rect 1924 1481 1960 1533
rect 3704 1544 4244 1588
rect 3704 1535 3756 1544
rect 3808 1535 3820 1544
rect 1324 1448 1960 1481
rect 2346 1503 2426 1528
rect 2346 1499 3517 1503
rect 2346 1465 2369 1499
rect 2403 1465 3517 1499
rect 2346 1461 3517 1465
rect 2346 1436 2426 1461
rect 2636 1403 2702 1415
rect 272 1349 278 1403
rect 332 1349 2642 1403
rect 2696 1349 2702 1403
rect 2636 1337 2702 1349
rect 3475 1308 3517 1461
rect 3704 1501 3741 1535
rect 3808 1501 3813 1535
rect 3704 1492 3756 1501
rect 3808 1492 3820 1501
rect 3872 1492 3884 1544
rect 3936 1492 3948 1544
rect 4000 1492 4012 1544
rect 4064 1492 4076 1544
rect 4128 1535 4140 1544
rect 4192 1535 4244 1544
rect 4135 1501 4140 1535
rect 4207 1501 4244 1535
rect 4128 1492 4140 1501
rect 4192 1492 4244 1501
rect 3704 1448 4244 1492
rect 3559 1343 3565 1395
rect 3617 1388 3623 1395
rect 4306 1388 4345 1778
rect 4558 1746 4597 1882
rect 4628 1851 4680 1857
rect 4625 1802 4628 1848
rect 4680 1802 4683 1848
rect 4875 1806 4904 1882
rect 4628 1793 4680 1799
rect 4875 1778 4980 1806
rect 4396 1713 4442 1746
rect 4396 1679 4402 1713
rect 4436 1679 4442 1713
rect 4396 1646 4442 1679
rect 4554 1726 4600 1746
rect 4704 1726 4750 1746
rect 4862 1726 4908 1746
rect 4554 1713 4750 1726
rect 4554 1679 4560 1713
rect 4594 1679 4710 1713
rect 4744 1679 4750 1713
rect 4554 1660 4750 1679
rect 4856 1674 4862 1726
rect 4914 1674 4920 1726
rect 4554 1646 4600 1660
rect 4704 1646 4750 1660
rect 4862 1646 4908 1674
rect 4402 1496 4430 1646
rect 4558 1601 4597 1646
rect 4552 1595 4604 1601
rect 4552 1537 4604 1543
rect 4952 1496 4980 1778
rect 5026 1728 5056 1913
rect 5694 1882 5740 1930
rect 5852 2036 5898 2082
rect 5852 2002 5858 2036
rect 5892 2002 5898 2036
rect 5852 1964 5898 2002
rect 5852 1930 5858 1964
rect 5892 1930 5898 1964
rect 5852 1882 5898 1930
rect 6002 2036 6048 2138
rect 6516 2082 6556 2288
rect 6862 2282 6868 2288
rect 6920 2282 6926 2334
rect 6985 2322 7015 2375
rect 6985 2293 7016 2322
rect 6002 2002 6008 2036
rect 6042 2002 6048 2036
rect 6002 1964 6048 2002
rect 6002 1930 6008 1964
rect 6042 1930 6048 1964
rect 6002 1882 6048 1930
rect 6160 2036 6206 2082
rect 6160 2002 6166 2036
rect 6200 2002 6206 2036
rect 6354 2036 6400 2082
rect 6354 2010 6360 2036
rect 6160 1964 6206 2002
rect 6160 1930 6166 1964
rect 6200 1930 6206 1964
rect 6244 2008 6360 2010
rect 6244 1956 6250 2008
rect 6302 2002 6360 2008
rect 6394 2002 6400 2036
rect 6302 1964 6400 2002
rect 6302 1956 6360 1964
rect 6244 1954 6360 1956
rect 6160 1882 6206 1930
rect 6354 1930 6360 1954
rect 6394 1930 6400 1964
rect 6354 1882 6400 1930
rect 6512 2036 6558 2082
rect 6512 2002 6518 2036
rect 6552 2002 6558 2036
rect 6662 2036 6708 2082
rect 6662 2002 6668 2036
rect 6702 2002 6708 2036
rect 6512 1964 6708 2002
rect 6512 1930 6518 1964
rect 6552 1936 6668 1964
rect 6552 1930 6558 1936
rect 6512 1882 6558 1930
rect 6662 1930 6668 1936
rect 6702 1930 6708 1964
rect 6662 1882 6708 1930
rect 6820 2036 6866 2082
rect 6820 2002 6826 2036
rect 6860 2002 6866 2036
rect 6986 2006 7016 2293
rect 6820 1964 6866 2002
rect 6820 1930 6826 1964
rect 6860 1930 6866 1964
rect 6968 1954 6974 2006
rect 7026 1954 7032 2006
rect 6820 1882 6866 1930
rect 6984 1914 7016 1954
rect 5111 1797 5117 1849
rect 5169 1842 5175 1849
rect 5620 1842 5672 1854
rect 5169 1840 5672 1842
rect 5169 1806 5628 1840
rect 5662 1806 5672 1840
rect 5169 1803 5672 1806
rect 5169 1797 5175 1803
rect 5620 1792 5672 1803
rect 5856 1834 5894 1882
rect 5934 1840 5986 1846
rect 5928 1834 5934 1840
rect 5856 1794 5934 1834
rect 5856 1744 5894 1794
rect 5928 1788 5934 1794
rect 5986 1788 5992 1840
rect 6164 1826 6204 1882
rect 6258 1826 6306 1838
rect 6164 1824 6306 1826
rect 6164 1792 6264 1824
rect 5934 1782 5986 1788
rect 6164 1744 6204 1792
rect 6258 1790 6264 1792
rect 6298 1790 6306 1824
rect 6258 1778 6306 1790
rect 5009 1676 5015 1728
rect 5067 1676 5073 1728
rect 5694 1712 5740 1744
rect 5694 1678 5700 1712
rect 5734 1678 5740 1712
rect 4402 1468 4980 1496
rect 3617 1349 4345 1388
rect 3617 1343 3623 1349
rect 5021 1308 5063 1676
rect 5694 1644 5740 1678
rect 5852 1712 5898 1744
rect 5852 1678 5858 1712
rect 5892 1678 5898 1712
rect 6002 1712 6048 1744
rect 6002 1682 6008 1712
rect 5852 1644 5898 1678
rect 6000 1678 6008 1682
rect 6042 1678 6048 1712
rect 5694 1588 5738 1644
rect 6000 1588 6048 1678
rect 6160 1712 6206 1744
rect 6160 1678 6166 1712
rect 6200 1678 6206 1712
rect 6160 1644 6206 1678
rect 5662 1544 6202 1588
rect 5662 1536 5714 1544
rect 5766 1536 5778 1544
rect 5662 1502 5700 1536
rect 5766 1502 5772 1536
rect 5662 1492 5714 1502
rect 5766 1492 5778 1502
rect 5830 1492 5842 1544
rect 5894 1492 5906 1544
rect 5958 1492 5970 1544
rect 6022 1492 6034 1544
rect 6086 1536 6098 1544
rect 6150 1536 6202 1544
rect 6094 1502 6098 1536
rect 6166 1502 6202 1536
rect 6086 1492 6098 1502
rect 6150 1492 6202 1502
rect 5662 1448 6202 1492
rect 5111 1343 5117 1395
rect 5169 1388 5175 1395
rect 6264 1388 6304 1778
rect 6516 1746 6556 1882
rect 6586 1852 6638 1858
rect 6584 1802 6586 1848
rect 6638 1802 6642 1848
rect 6834 1806 6862 1882
rect 6586 1794 6638 1800
rect 6834 1778 6936 1806
rect 6354 1714 6400 1746
rect 6354 1680 6360 1714
rect 6394 1680 6400 1714
rect 6354 1646 6400 1680
rect 6512 1726 6558 1746
rect 6662 1726 6708 1746
rect 6820 1726 6866 1746
rect 6512 1714 6708 1726
rect 6512 1680 6518 1714
rect 6552 1680 6668 1714
rect 6702 1680 6708 1714
rect 6512 1660 6708 1680
rect 6814 1674 6820 1726
rect 6872 1674 6878 1726
rect 6512 1646 6558 1660
rect 6662 1646 6708 1660
rect 6820 1646 6866 1674
rect 6360 1496 6388 1646
rect 6516 1602 6556 1646
rect 6510 1596 6562 1602
rect 6510 1538 6562 1544
rect 6908 1496 6936 1778
rect 6984 1728 7014 1914
rect 6968 1676 6974 1728
rect 7026 1676 7032 1728
rect 6360 1468 6936 1496
rect 6908 1404 6936 1468
rect 5169 1350 6304 1388
rect 6346 1376 6936 1404
rect 5169 1349 5572 1350
rect 5169 1343 5175 1349
rect 3475 1266 5063 1308
rect 5035 1225 5087 1231
rect 3472 1141 4907 1180
rect 6346 1213 6374 1376
rect 6908 1374 6936 1376
rect 5087 1185 6374 1213
rect 5035 1167 5087 1173
rect 1348 1007 1880 1050
rect 1348 998 1398 1007
rect 1450 998 1462 1007
rect 1348 964 1383 998
rect 1450 964 1455 998
rect 1348 955 1398 964
rect 1450 955 1462 964
rect 1514 955 1526 1007
rect 1578 955 1590 1007
rect 1642 955 1654 1007
rect 1706 955 1718 1007
rect 1770 998 1782 1007
rect 1834 998 1880 1007
rect 1777 964 1782 998
rect 1849 964 1880 998
rect 3472 983 3511 1141
rect 4738 1099 4744 1106
rect 4558 1060 4744 1099
rect 1770 955 1782 964
rect 1834 955 1880 964
rect 550 936 622 940
rect 550 884 560 936
rect 612 884 622 936
rect 696 934 768 940
rect 550 872 566 884
rect 607 872 622 884
rect 682 932 768 934
rect 682 880 702 932
rect 754 880 768 932
rect 682 878 710 880
rect 550 842 622 872
rect 696 872 710 878
rect 751 872 768 880
rect 696 842 768 872
rect 840 917 912 946
rect 840 877 856 917
rect 897 877 912 917
rect 840 848 912 877
rect 994 917 1066 946
rect 994 877 1009 917
rect 1050 877 1066 917
rect 1348 910 1880 955
rect 994 848 1066 877
rect 564 802 608 842
rect 856 782 900 848
rect 378 774 433 780
rect 846 730 852 782
rect 904 730 910 782
rect 378 489 433 719
rect 856 690 900 730
rect 1008 690 1052 848
rect 1407 844 1448 910
rect 1693 844 1735 910
rect 1941 907 2687 952
rect 1404 797 1450 844
rect 1404 763 1410 797
rect 1444 763 1450 797
rect 1404 725 1450 763
rect 1404 691 1410 725
rect 1444 691 1450 725
rect 708 646 900 690
rect 372 434 378 489
rect 433 434 439 489
rect 708 412 752 646
rect 998 638 1004 690
rect 1056 638 1062 690
rect 1404 644 1450 691
rect 1562 797 1608 844
rect 1562 763 1568 797
rect 1602 763 1608 797
rect 1562 725 1608 763
rect 1562 691 1568 725
rect 1602 691 1608 725
rect 1562 644 1608 691
rect 1692 797 1738 844
rect 1692 763 1698 797
rect 1732 763 1738 797
rect 1692 725 1738 763
rect 1692 691 1698 725
rect 1732 691 1738 725
rect 1692 644 1738 691
rect 1850 841 1896 844
rect 1941 841 1986 907
rect 1850 797 1986 841
rect 1850 763 1856 797
rect 1890 796 1986 797
rect 2024 797 2070 844
rect 1890 763 1896 796
rect 1850 725 1896 763
rect 2024 763 2030 797
rect 2064 763 2070 797
rect 2024 728 2070 763
rect 1998 726 2070 728
rect 1850 691 1856 725
rect 1890 691 1896 725
rect 1850 644 1896 691
rect 1928 725 2070 726
rect 1928 701 2030 725
rect 1928 684 1935 701
rect 1929 649 1935 684
rect 1987 691 2030 701
rect 2064 691 2070 725
rect 1987 684 2070 691
rect 1987 649 1993 684
rect 2024 644 2070 684
rect 2182 800 2228 844
rect 2366 800 2412 844
rect 2182 797 2412 800
rect 2182 763 2188 797
rect 2222 763 2372 797
rect 2406 763 2412 797
rect 2182 725 2412 763
rect 2182 691 2188 725
rect 2222 691 2372 725
rect 2406 691 2412 725
rect 2182 674 2412 691
rect 2182 644 2228 674
rect 2366 644 2412 674
rect 2524 797 2570 844
rect 2524 763 2530 797
rect 2564 763 2570 797
rect 2642 773 2687 907
rect 3118 944 3511 983
rect 3724 1006 4264 1050
rect 3724 954 3776 1006
rect 3828 997 3840 1006
rect 3892 997 3904 1006
rect 3956 997 3968 1006
rect 4020 997 4032 1006
rect 4084 997 4096 1006
rect 4148 997 4160 1006
rect 3831 963 3840 997
rect 3903 963 3904 997
rect 4084 963 4085 997
rect 4148 963 4157 997
rect 3828 954 3840 963
rect 3892 954 3904 963
rect 3956 954 3968 963
rect 4020 954 4032 963
rect 4084 954 4096 963
rect 4148 954 4160 963
rect 4212 954 4264 1006
rect 2774 900 2816 901
rect 2758 892 2816 900
rect 2758 840 2769 892
rect 2821 840 2827 892
rect 3118 844 3157 944
rect 3724 910 4264 954
rect 3741 854 3787 910
rect 3736 853 3787 854
rect 2758 797 2816 840
rect 2524 725 2570 763
rect 2524 691 2530 725
rect 2564 691 2570 725
rect 2524 684 2570 691
rect 2613 745 2715 773
rect 2613 711 2647 745
rect 2681 711 2715 745
rect 2524 644 2574 684
rect 2613 683 2715 711
rect 2758 763 2776 797
rect 2810 763 2816 797
rect 2758 725 2816 763
rect 2758 691 2776 725
rect 2810 691 2816 725
rect 1008 584 1052 638
rect 1245 603 1328 622
rect 852 540 1052 584
rect 1148 601 1328 603
rect 1148 549 1155 601
rect 1207 591 1328 601
rect 1207 557 1269 591
rect 1303 557 1328 591
rect 1207 549 1328 557
rect 1148 548 1328 549
rect 852 418 896 540
rect 1245 527 1328 548
rect 1568 610 1602 644
rect 1568 600 1820 610
rect 1568 548 1758 600
rect 1810 548 1820 600
rect 1568 538 1820 548
rect 1568 506 1608 538
rect 1853 506 1892 644
rect 2185 506 2224 644
rect 2255 607 2325 613
rect 2255 598 2331 607
rect 2255 546 2270 598
rect 2322 546 2331 598
rect 2255 537 2331 546
rect 2255 531 2325 537
rect 2368 506 2407 644
rect 2530 610 2574 644
rect 2758 644 2816 691
rect 2928 797 2974 844
rect 2928 763 2934 797
rect 2968 784 2974 797
rect 3114 797 3160 844
rect 3114 784 3120 797
rect 2968 763 3120 784
rect 3154 763 3160 797
rect 3272 797 3318 844
rect 3272 787 3278 797
rect 3312 787 3318 797
rect 3736 807 3782 853
rect 2928 725 3160 763
rect 3262 735 3268 787
rect 3320 735 3326 787
rect 3736 773 3742 807
rect 3776 773 3782 807
rect 3736 735 3782 773
rect 2928 691 2934 725
rect 2968 691 3120 725
rect 3154 691 3160 725
rect 2928 674 3160 691
rect 2928 644 2974 674
rect 3114 644 3160 674
rect 3272 725 3318 735
rect 3272 691 3278 725
rect 3312 691 3318 725
rect 3272 644 3318 691
rect 3736 701 3742 735
rect 3776 701 3782 735
rect 3736 654 3782 701
rect 3894 807 3940 854
rect 3894 773 3900 807
rect 3934 773 3940 807
rect 3894 735 3940 773
rect 3894 701 3900 735
rect 3934 701 3940 735
rect 3894 654 3940 701
rect 4044 807 4090 910
rect 4558 854 4597 1060
rect 4738 1054 4744 1060
rect 4796 1054 4802 1106
rect 4868 854 4907 1141
rect 4044 773 4050 807
rect 4084 773 4090 807
rect 4044 735 4090 773
rect 4044 701 4050 735
rect 4084 701 4090 735
rect 4044 654 4090 701
rect 4202 807 4248 854
rect 4202 773 4208 807
rect 4242 773 4248 807
rect 4396 807 4442 854
rect 4396 781 4402 807
rect 4202 735 4248 773
rect 4202 701 4208 735
rect 4242 701 4248 735
rect 4285 779 4402 781
rect 4285 727 4292 779
rect 4344 773 4402 779
rect 4436 773 4442 807
rect 4344 735 4442 773
rect 4344 727 4402 735
rect 4285 726 4402 727
rect 4202 654 4248 701
rect 4396 701 4402 726
rect 4436 701 4442 735
rect 4396 654 4442 701
rect 4554 807 4600 854
rect 4554 773 4560 807
rect 4594 774 4600 807
rect 4704 807 4750 854
rect 4704 774 4710 807
rect 4594 773 4710 774
rect 4744 773 4750 807
rect 4554 735 4750 773
rect 4554 701 4560 735
rect 4594 708 4710 735
rect 4594 701 4600 708
rect 4554 654 4600 701
rect 4704 701 4710 708
rect 4744 701 4750 735
rect 4704 654 4750 701
rect 4862 807 4908 854
rect 4862 773 4868 807
rect 4902 773 4908 807
rect 5027 778 5057 787
rect 4862 735 4908 773
rect 4862 701 4868 735
rect 4902 701 4908 735
rect 5010 726 5016 778
rect 5068 726 5074 778
rect 4862 654 4908 701
rect 5026 685 5057 726
rect 2758 610 2802 644
rect 2530 566 2656 610
rect 1242 486 1248 490
rect 1138 442 1248 486
rect 1138 418 1182 442
rect 1242 438 1248 442
rect 1300 438 1306 490
rect 1404 473 1450 506
rect 1404 439 1410 473
rect 1444 439 1450 473
rect 1404 435 1450 439
rect 378 390 434 396
rect 550 390 622 412
rect 434 384 622 390
rect 434 344 565 384
rect 606 344 622 384
rect 434 334 622 344
rect 378 328 434 334
rect 550 314 622 334
rect 696 384 768 412
rect 696 344 712 384
rect 753 344 768 384
rect 696 314 768 344
rect 840 389 912 418
rect 840 349 856 389
rect 897 349 912 389
rect 840 320 912 349
rect 994 390 1182 418
rect 994 350 1010 390
rect 1051 374 1182 390
rect 1399 406 1450 435
rect 1562 473 1608 506
rect 1562 439 1568 473
rect 1602 439 1608 473
rect 1692 473 1738 506
rect 1692 444 1698 473
rect 1562 406 1608 439
rect 1690 439 1698 444
rect 1732 444 1738 473
rect 1850 473 1896 506
rect 2024 490 2070 506
rect 1732 439 1740 444
rect 1051 350 1066 374
rect 1399 360 1449 406
rect 1690 360 1740 439
rect 1850 439 1856 473
rect 1890 439 1896 473
rect 1850 406 1896 439
rect 2014 438 2020 490
rect 2072 438 2078 490
rect 2182 473 2228 506
rect 2182 439 2188 473
rect 2222 439 2228 473
rect 2024 406 2070 438
rect 2182 406 2228 439
rect 2366 473 2412 506
rect 2524 488 2570 506
rect 2366 439 2372 473
rect 2406 439 2412 473
rect 2366 406 2412 439
rect 2516 436 2522 488
rect 2574 436 2580 488
rect 2524 406 2570 436
rect 2024 374 2068 406
rect 2612 374 2656 566
rect 994 320 1066 350
rect 1324 305 1960 360
rect 2024 330 2656 374
rect 2694 566 2802 610
rect 2832 596 2904 606
rect 2694 368 2738 566
rect 2832 544 2842 596
rect 2894 544 2904 596
rect 2832 534 2904 544
rect 2933 506 2972 644
rect 3118 506 3157 644
rect 3272 600 3316 644
rect 3268 594 3320 600
rect 3555 569 3561 621
rect 3613 614 3619 621
rect 3662 614 3713 626
rect 3613 611 3713 614
rect 3613 577 3670 611
rect 3704 577 3713 611
rect 3613 575 3713 577
rect 3613 569 3619 575
rect 3662 563 3713 575
rect 3897 605 3936 654
rect 3976 612 4027 617
rect 3970 605 3976 612
rect 3897 566 3976 605
rect 3268 536 3320 542
rect 3897 516 3936 566
rect 3970 560 3976 566
rect 4028 560 4034 612
rect 4206 598 4245 654
rect 4300 598 4347 609
rect 4206 596 4347 598
rect 4206 563 4306 596
rect 3976 554 4027 560
rect 4206 516 4245 563
rect 4300 562 4306 563
rect 4340 562 4347 596
rect 4300 550 4347 562
rect 2766 500 2818 506
rect 2766 442 2776 448
rect 2770 439 2776 442
rect 2810 442 2818 448
rect 2928 473 2974 506
rect 2810 439 2816 442
rect 2770 406 2816 439
rect 2928 439 2934 473
rect 2968 439 2974 473
rect 2928 406 2974 439
rect 3114 473 3160 506
rect 3114 439 3120 473
rect 3154 439 3160 473
rect 3114 406 3160 439
rect 3272 473 3318 506
rect 3272 439 3278 473
rect 3312 439 3318 473
rect 3272 406 3318 439
rect 3274 368 3318 406
rect 2694 324 3318 368
rect 3736 483 3782 516
rect 3736 449 3742 483
rect 3776 449 3782 483
rect 3736 416 3782 449
rect 3894 483 3940 516
rect 3894 449 3900 483
rect 3934 449 3940 483
rect 4044 483 4090 516
rect 4044 454 4050 483
rect 3894 416 3940 449
rect 4042 449 4050 454
rect 4084 449 4090 483
rect 4042 416 4090 449
rect 4202 483 4248 516
rect 4202 449 4208 483
rect 4242 449 4248 483
rect 4202 416 4248 449
rect 3736 360 3780 416
rect 4042 360 4089 416
rect 1324 253 1360 305
rect 1412 253 1424 305
rect 1476 296 1488 305
rect 1540 296 1552 305
rect 1604 296 1616 305
rect 1668 296 1680 305
rect 1732 296 1744 305
rect 1796 296 1808 305
rect 1479 262 1488 296
rect 1551 262 1552 296
rect 1732 262 1733 296
rect 1796 262 1805 296
rect 1476 253 1488 262
rect 1540 253 1552 262
rect 1604 253 1616 262
rect 1668 253 1680 262
rect 1732 253 1744 262
rect 1796 253 1808 262
rect 1860 253 1872 305
rect 1924 253 1960 305
rect 3704 316 4244 360
rect 3704 307 3756 316
rect 3808 307 3820 316
rect 1324 220 1960 253
rect 2346 275 2426 300
rect 2346 271 3517 275
rect 2346 237 2369 271
rect 2403 237 3517 271
rect 2346 233 3517 237
rect 2346 208 2426 233
rect 2636 175 2702 187
rect 272 121 278 175
rect 332 121 2642 175
rect 2696 121 2702 175
rect 2636 109 2702 121
rect 3475 80 3517 233
rect 3704 273 3741 307
rect 3808 273 3813 307
rect 3704 264 3756 273
rect 3808 264 3820 273
rect 3872 264 3884 316
rect 3936 264 3948 316
rect 4000 264 4012 316
rect 4064 264 4076 316
rect 4128 307 4140 316
rect 4192 307 4244 316
rect 4135 273 4140 307
rect 4207 273 4244 307
rect 4128 264 4140 273
rect 4192 264 4244 273
rect 3704 220 4244 264
rect 3559 115 3565 167
rect 3617 160 3623 167
rect 4306 160 4345 550
rect 4558 518 4597 654
rect 4628 623 4680 629
rect 4625 574 4628 620
rect 4680 574 4683 620
rect 4875 578 4904 654
rect 4628 565 4680 571
rect 4875 550 4980 578
rect 4396 485 4442 518
rect 4396 451 4402 485
rect 4436 451 4442 485
rect 4396 418 4442 451
rect 4554 498 4600 518
rect 4704 498 4750 518
rect 4862 498 4908 518
rect 4554 485 4750 498
rect 4554 451 4560 485
rect 4594 451 4710 485
rect 4744 451 4750 485
rect 4554 432 4750 451
rect 4856 446 4862 498
rect 4914 446 4920 498
rect 4554 418 4600 432
rect 4704 418 4750 432
rect 4862 418 4908 446
rect 4402 268 4430 418
rect 4558 373 4597 418
rect 4552 367 4604 373
rect 4552 309 4604 315
rect 4952 268 4980 550
rect 5026 500 5056 685
rect 5009 448 5015 500
rect 5067 448 5073 500
rect 4402 240 4980 268
rect 3617 121 4345 160
rect 3617 115 3623 121
rect 5021 80 5063 448
rect 3475 38 5063 80
<< via1 >>
rect 1398 19418 1450 19427
rect 1462 19418 1514 19427
rect 1398 19384 1417 19418
rect 1417 19384 1450 19418
rect 1462 19384 1489 19418
rect 1489 19384 1514 19418
rect 1398 19375 1450 19384
rect 1462 19375 1514 19384
rect 1526 19418 1578 19427
rect 1526 19384 1527 19418
rect 1527 19384 1561 19418
rect 1561 19384 1578 19418
rect 1526 19375 1578 19384
rect 1590 19418 1642 19427
rect 1590 19384 1599 19418
rect 1599 19384 1633 19418
rect 1633 19384 1642 19418
rect 1590 19375 1642 19384
rect 1654 19418 1706 19427
rect 1654 19384 1671 19418
rect 1671 19384 1705 19418
rect 1705 19384 1706 19418
rect 1654 19375 1706 19384
rect 1718 19418 1770 19427
rect 1782 19418 1834 19427
rect 1718 19384 1743 19418
rect 1743 19384 1770 19418
rect 1782 19384 1815 19418
rect 1815 19384 1834 19418
rect 1718 19375 1770 19384
rect 1782 19375 1834 19384
rect 560 19332 612 19356
rect 560 19304 566 19332
rect 566 19304 607 19332
rect 607 19304 612 19332
rect 702 19332 754 19352
rect 702 19300 710 19332
rect 710 19300 751 19332
rect 751 19300 754 19332
rect 378 19139 433 19194
rect 852 19150 904 19202
rect 378 18854 433 18909
rect 1004 19058 1056 19110
rect 1935 19069 1987 19121
rect 3776 19417 3828 19426
rect 3840 19417 3892 19426
rect 3904 19417 3956 19426
rect 3968 19417 4020 19426
rect 4032 19417 4084 19426
rect 4096 19417 4148 19426
rect 4160 19417 4212 19426
rect 3776 19383 3797 19417
rect 3797 19383 3828 19417
rect 3840 19383 3869 19417
rect 3869 19383 3892 19417
rect 3904 19383 3941 19417
rect 3941 19383 3956 19417
rect 3968 19383 3975 19417
rect 3975 19383 4013 19417
rect 4013 19383 4020 19417
rect 4032 19383 4047 19417
rect 4047 19383 4084 19417
rect 4096 19383 4119 19417
rect 4119 19383 4148 19417
rect 4160 19383 4191 19417
rect 4191 19383 4212 19417
rect 3776 19374 3828 19383
rect 3840 19374 3892 19383
rect 3904 19374 3956 19383
rect 3968 19374 4020 19383
rect 4032 19374 4084 19383
rect 4096 19374 4148 19383
rect 4160 19374 4212 19383
rect 2769 19260 2821 19312
rect 1155 18969 1207 19021
rect 1758 19011 1810 19020
rect 1758 18977 1773 19011
rect 1773 18977 1807 19011
rect 1807 18977 1810 19011
rect 1758 18968 1810 18977
rect 2270 19009 2322 19018
rect 2270 18975 2273 19009
rect 2273 18975 2307 19009
rect 2307 18975 2322 19009
rect 2270 18966 2322 18975
rect 3268 19183 3278 19207
rect 3278 19183 3312 19207
rect 3312 19183 3320 19207
rect 3268 19155 3320 19183
rect 4744 19474 4796 19526
rect 5029 19556 5081 19608
rect 5734 19416 5786 19426
rect 5798 19416 5850 19426
rect 5862 19416 5914 19426
rect 5926 19416 5978 19426
rect 5990 19416 6042 19426
rect 6054 19416 6106 19426
rect 6118 19416 6170 19426
rect 5734 19382 5756 19416
rect 5756 19382 5786 19416
rect 5798 19382 5828 19416
rect 5828 19382 5850 19416
rect 5862 19382 5900 19416
rect 5900 19382 5914 19416
rect 5926 19382 5934 19416
rect 5934 19382 5972 19416
rect 5972 19382 5978 19416
rect 5990 19382 6006 19416
rect 6006 19382 6042 19416
rect 6054 19382 6078 19416
rect 6078 19382 6106 19416
rect 6118 19382 6150 19416
rect 6150 19382 6170 19416
rect 5734 19374 5786 19382
rect 5798 19374 5850 19382
rect 5862 19374 5914 19382
rect 5926 19374 5978 19382
rect 5990 19374 6042 19382
rect 6054 19374 6106 19382
rect 6118 19374 6170 19382
rect 4292 19147 4344 19199
rect 5016 19146 5068 19198
rect 1248 18858 1300 18910
rect 378 18754 434 18810
rect 2020 18893 2072 18910
rect 2020 18859 2030 18893
rect 2030 18859 2064 18893
rect 2064 18859 2072 18893
rect 2020 18858 2072 18859
rect 2522 18893 2574 18908
rect 2522 18859 2530 18893
rect 2530 18859 2564 18893
rect 2564 18859 2574 18893
rect 2522 18856 2574 18859
rect 2842 19007 2894 19016
rect 2842 18973 2857 19007
rect 2857 18973 2891 19007
rect 2891 18973 2894 19007
rect 2842 18964 2894 18973
rect 3268 18962 3320 19014
rect 3561 18989 3613 19041
rect 3976 19022 4028 19032
rect 3976 18988 3984 19022
rect 3984 18988 4018 19022
rect 4018 18988 4028 19022
rect 3976 18980 4028 18988
rect 2766 18893 2818 18920
rect 2766 18868 2776 18893
rect 2776 18868 2810 18893
rect 2810 18868 2818 18893
rect 1360 18716 1412 18725
rect 1360 18682 1373 18716
rect 1373 18682 1407 18716
rect 1407 18682 1412 18716
rect 1360 18673 1412 18682
rect 1424 18716 1476 18725
rect 1488 18716 1540 18725
rect 1552 18716 1604 18725
rect 1616 18716 1668 18725
rect 1680 18716 1732 18725
rect 1744 18716 1796 18725
rect 1808 18716 1860 18725
rect 1424 18682 1445 18716
rect 1445 18682 1476 18716
rect 1488 18682 1517 18716
rect 1517 18682 1540 18716
rect 1552 18682 1589 18716
rect 1589 18682 1604 18716
rect 1616 18682 1623 18716
rect 1623 18682 1661 18716
rect 1661 18682 1668 18716
rect 1680 18682 1695 18716
rect 1695 18682 1732 18716
rect 1744 18682 1767 18716
rect 1767 18682 1796 18716
rect 1808 18682 1839 18716
rect 1839 18682 1860 18716
rect 1424 18673 1476 18682
rect 1488 18673 1540 18682
rect 1552 18673 1604 18682
rect 1616 18673 1668 18682
rect 1680 18673 1732 18682
rect 1744 18673 1796 18682
rect 1808 18673 1860 18682
rect 1872 18716 1924 18725
rect 1872 18682 1877 18716
rect 1877 18682 1911 18716
rect 1911 18682 1924 18716
rect 1872 18673 1924 18682
rect 3756 18727 3808 18736
rect 3820 18727 3872 18736
rect 278 18541 332 18595
rect 3756 18693 3775 18727
rect 3775 18693 3808 18727
rect 3820 18693 3847 18727
rect 3847 18693 3872 18727
rect 3756 18684 3808 18693
rect 3820 18684 3872 18693
rect 3884 18727 3936 18736
rect 3884 18693 3885 18727
rect 3885 18693 3919 18727
rect 3919 18693 3936 18727
rect 3884 18684 3936 18693
rect 3948 18727 4000 18736
rect 3948 18693 3957 18727
rect 3957 18693 3991 18727
rect 3991 18693 4000 18727
rect 3948 18684 4000 18693
rect 4012 18727 4064 18736
rect 4012 18693 4029 18727
rect 4029 18693 4063 18727
rect 4063 18693 4064 18727
rect 4012 18684 4064 18693
rect 4076 18727 4128 18736
rect 4140 18727 4192 18736
rect 4076 18693 4101 18727
rect 4101 18693 4128 18727
rect 4140 18693 4173 18727
rect 4173 18693 4192 18727
rect 4076 18684 4128 18693
rect 4140 18684 4192 18693
rect 3565 18535 3617 18587
rect 4628 19034 4680 19043
rect 4628 19000 4637 19034
rect 4637 19000 4671 19034
rect 4671 19000 4680 19034
rect 4628 18991 4680 19000
rect 4862 18905 4914 18918
rect 4862 18871 4868 18905
rect 4868 18871 4902 18905
rect 4902 18871 4914 18905
rect 4862 18866 4914 18871
rect 4552 18735 4604 18787
rect 6868 19474 6920 19526
rect 6250 19148 6302 19200
rect 6974 19146 7026 19198
rect 5117 18989 5169 19041
rect 5934 19022 5986 19032
rect 5934 18988 5942 19022
rect 5942 18988 5976 19022
rect 5976 18988 5986 19022
rect 5934 18980 5986 18988
rect 5015 18868 5067 18920
rect 5714 18728 5766 18736
rect 5778 18728 5830 18736
rect 5714 18694 5734 18728
rect 5734 18694 5766 18728
rect 5778 18694 5806 18728
rect 5806 18694 5830 18728
rect 5714 18684 5766 18694
rect 5778 18684 5830 18694
rect 5842 18728 5894 18736
rect 5842 18694 5844 18728
rect 5844 18694 5878 18728
rect 5878 18694 5894 18728
rect 5842 18684 5894 18694
rect 5906 18728 5958 18736
rect 5906 18694 5916 18728
rect 5916 18694 5950 18728
rect 5950 18694 5958 18728
rect 5906 18684 5958 18694
rect 5970 18728 6022 18736
rect 5970 18694 5988 18728
rect 5988 18694 6022 18728
rect 5970 18684 6022 18694
rect 6034 18728 6086 18736
rect 6098 18728 6150 18736
rect 6034 18694 6060 18728
rect 6060 18694 6086 18728
rect 6098 18694 6132 18728
rect 6132 18694 6150 18728
rect 6034 18684 6086 18694
rect 6098 18684 6150 18694
rect 5117 18535 5169 18587
rect 6586 19034 6638 19044
rect 6586 19000 6596 19034
rect 6596 19000 6630 19034
rect 6630 19000 6638 19034
rect 6586 18992 6638 19000
rect 6820 18906 6872 18918
rect 6820 18872 6826 18906
rect 6826 18872 6860 18906
rect 6860 18872 6872 18906
rect 6820 18866 6872 18872
rect 6510 18736 6562 18788
rect 6974 18868 7026 18920
rect 5035 18365 5087 18417
rect 6512 18450 6564 18502
rect 1398 18190 1450 18199
rect 1462 18190 1514 18199
rect 1398 18156 1417 18190
rect 1417 18156 1450 18190
rect 1462 18156 1489 18190
rect 1489 18156 1514 18190
rect 1398 18147 1450 18156
rect 1462 18147 1514 18156
rect 1526 18190 1578 18199
rect 1526 18156 1527 18190
rect 1527 18156 1561 18190
rect 1561 18156 1578 18190
rect 1526 18147 1578 18156
rect 1590 18190 1642 18199
rect 1590 18156 1599 18190
rect 1599 18156 1633 18190
rect 1633 18156 1642 18190
rect 1590 18147 1642 18156
rect 1654 18190 1706 18199
rect 1654 18156 1671 18190
rect 1671 18156 1705 18190
rect 1705 18156 1706 18190
rect 1654 18147 1706 18156
rect 1718 18190 1770 18199
rect 1782 18190 1834 18199
rect 1718 18156 1743 18190
rect 1743 18156 1770 18190
rect 1782 18156 1815 18190
rect 1815 18156 1834 18190
rect 1718 18147 1770 18156
rect 1782 18147 1834 18156
rect 560 18104 612 18128
rect 560 18076 566 18104
rect 566 18076 607 18104
rect 607 18076 612 18104
rect 702 18104 754 18124
rect 702 18072 710 18104
rect 710 18072 751 18104
rect 751 18072 754 18104
rect 378 17911 433 17966
rect 852 17922 904 17974
rect 378 17626 433 17681
rect 1004 17830 1056 17882
rect 1935 17841 1987 17893
rect 3776 18189 3828 18198
rect 3840 18189 3892 18198
rect 3904 18189 3956 18198
rect 3968 18189 4020 18198
rect 4032 18189 4084 18198
rect 4096 18189 4148 18198
rect 4160 18189 4212 18198
rect 3776 18155 3797 18189
rect 3797 18155 3828 18189
rect 3840 18155 3869 18189
rect 3869 18155 3892 18189
rect 3904 18155 3941 18189
rect 3941 18155 3956 18189
rect 3968 18155 3975 18189
rect 3975 18155 4013 18189
rect 4013 18155 4020 18189
rect 4032 18155 4047 18189
rect 4047 18155 4084 18189
rect 4096 18155 4119 18189
rect 4119 18155 4148 18189
rect 4160 18155 4191 18189
rect 4191 18155 4212 18189
rect 3776 18146 3828 18155
rect 3840 18146 3892 18155
rect 3904 18146 3956 18155
rect 3968 18146 4020 18155
rect 4032 18146 4084 18155
rect 4096 18146 4148 18155
rect 4160 18146 4212 18155
rect 2769 18032 2821 18084
rect 1155 17741 1207 17793
rect 1758 17783 1810 17792
rect 1758 17749 1773 17783
rect 1773 17749 1807 17783
rect 1807 17749 1810 17783
rect 1758 17740 1810 17749
rect 2270 17781 2322 17790
rect 2270 17747 2273 17781
rect 2273 17747 2307 17781
rect 2307 17747 2322 17781
rect 2270 17738 2322 17747
rect 3268 17955 3278 17979
rect 3278 17955 3312 17979
rect 3312 17955 3320 17979
rect 3268 17927 3320 17955
rect 4744 18246 4796 18298
rect 5734 18188 5786 18198
rect 5798 18188 5850 18198
rect 5862 18188 5914 18198
rect 5926 18188 5978 18198
rect 5990 18188 6042 18198
rect 6054 18188 6106 18198
rect 6118 18188 6170 18198
rect 5734 18154 5756 18188
rect 5756 18154 5786 18188
rect 5798 18154 5828 18188
rect 5828 18154 5850 18188
rect 5862 18154 5900 18188
rect 5900 18154 5914 18188
rect 5926 18154 5934 18188
rect 5934 18154 5972 18188
rect 5972 18154 5978 18188
rect 5990 18154 6006 18188
rect 6006 18154 6042 18188
rect 6054 18154 6078 18188
rect 6078 18154 6106 18188
rect 6118 18154 6150 18188
rect 6150 18154 6170 18188
rect 5734 18146 5786 18154
rect 5798 18146 5850 18154
rect 5862 18146 5914 18154
rect 5926 18146 5978 18154
rect 5990 18146 6042 18154
rect 6054 18146 6106 18154
rect 6118 18146 6170 18154
rect 4292 17919 4344 17971
rect 5016 17918 5068 17970
rect 1248 17630 1300 17682
rect 378 17526 434 17582
rect 2020 17665 2072 17682
rect 2020 17631 2030 17665
rect 2030 17631 2064 17665
rect 2064 17631 2072 17665
rect 2020 17630 2072 17631
rect 2522 17665 2574 17680
rect 2522 17631 2530 17665
rect 2530 17631 2564 17665
rect 2564 17631 2574 17665
rect 2522 17628 2574 17631
rect 2842 17779 2894 17788
rect 2842 17745 2857 17779
rect 2857 17745 2891 17779
rect 2891 17745 2894 17779
rect 2842 17736 2894 17745
rect 3268 17734 3320 17786
rect 3561 17761 3613 17813
rect 3976 17794 4028 17804
rect 3976 17760 3984 17794
rect 3984 17760 4018 17794
rect 4018 17760 4028 17794
rect 3976 17752 4028 17760
rect 2766 17665 2818 17692
rect 2766 17640 2776 17665
rect 2776 17640 2810 17665
rect 2810 17640 2818 17665
rect 1360 17488 1412 17497
rect 1360 17454 1373 17488
rect 1373 17454 1407 17488
rect 1407 17454 1412 17488
rect 1360 17445 1412 17454
rect 1424 17488 1476 17497
rect 1488 17488 1540 17497
rect 1552 17488 1604 17497
rect 1616 17488 1668 17497
rect 1680 17488 1732 17497
rect 1744 17488 1796 17497
rect 1808 17488 1860 17497
rect 1424 17454 1445 17488
rect 1445 17454 1476 17488
rect 1488 17454 1517 17488
rect 1517 17454 1540 17488
rect 1552 17454 1589 17488
rect 1589 17454 1604 17488
rect 1616 17454 1623 17488
rect 1623 17454 1661 17488
rect 1661 17454 1668 17488
rect 1680 17454 1695 17488
rect 1695 17454 1732 17488
rect 1744 17454 1767 17488
rect 1767 17454 1796 17488
rect 1808 17454 1839 17488
rect 1839 17454 1860 17488
rect 1424 17445 1476 17454
rect 1488 17445 1540 17454
rect 1552 17445 1604 17454
rect 1616 17445 1668 17454
rect 1680 17445 1732 17454
rect 1744 17445 1796 17454
rect 1808 17445 1860 17454
rect 1872 17488 1924 17497
rect 1872 17454 1877 17488
rect 1877 17454 1911 17488
rect 1911 17454 1924 17488
rect 1872 17445 1924 17454
rect 3756 17499 3808 17508
rect 3820 17499 3872 17508
rect 278 17313 332 17367
rect 3756 17465 3775 17499
rect 3775 17465 3808 17499
rect 3820 17465 3847 17499
rect 3847 17465 3872 17499
rect 3756 17456 3808 17465
rect 3820 17456 3872 17465
rect 3884 17499 3936 17508
rect 3884 17465 3885 17499
rect 3885 17465 3919 17499
rect 3919 17465 3936 17499
rect 3884 17456 3936 17465
rect 3948 17499 4000 17508
rect 3948 17465 3957 17499
rect 3957 17465 3991 17499
rect 3991 17465 4000 17499
rect 3948 17456 4000 17465
rect 4012 17499 4064 17508
rect 4012 17465 4029 17499
rect 4029 17465 4063 17499
rect 4063 17465 4064 17499
rect 4012 17456 4064 17465
rect 4076 17499 4128 17508
rect 4140 17499 4192 17508
rect 4076 17465 4101 17499
rect 4101 17465 4128 17499
rect 4140 17465 4173 17499
rect 4173 17465 4192 17499
rect 4076 17456 4128 17465
rect 4140 17456 4192 17465
rect 3565 17307 3617 17359
rect 4628 17806 4680 17815
rect 4628 17772 4637 17806
rect 4637 17772 4671 17806
rect 4671 17772 4680 17806
rect 4628 17763 4680 17772
rect 4862 17677 4914 17690
rect 4862 17643 4868 17677
rect 4868 17643 4902 17677
rect 4902 17643 4914 17677
rect 4862 17638 4914 17643
rect 4552 17507 4604 17559
rect 6843 18246 6895 18298
rect 6250 17920 6302 17972
rect 6974 17918 7026 17970
rect 5197 17761 5249 17813
rect 5934 17794 5986 17804
rect 5934 17760 5942 17794
rect 5942 17760 5976 17794
rect 5976 17760 5986 17794
rect 5934 17752 5986 17760
rect 5015 17640 5067 17692
rect 5714 17500 5766 17508
rect 5778 17500 5830 17508
rect 5714 17466 5734 17500
rect 5734 17466 5766 17500
rect 5778 17466 5806 17500
rect 5806 17466 5830 17500
rect 5714 17456 5766 17466
rect 5778 17456 5830 17466
rect 5842 17500 5894 17508
rect 5842 17466 5844 17500
rect 5844 17466 5878 17500
rect 5878 17466 5894 17500
rect 5842 17456 5894 17466
rect 5906 17500 5958 17508
rect 5906 17466 5916 17500
rect 5916 17466 5950 17500
rect 5950 17466 5958 17500
rect 5906 17456 5958 17466
rect 5970 17500 6022 17508
rect 5970 17466 5988 17500
rect 5988 17466 6022 17500
rect 5970 17456 6022 17466
rect 6034 17500 6086 17508
rect 6098 17500 6150 17508
rect 6034 17466 6060 17500
rect 6060 17466 6086 17500
rect 6098 17466 6132 17500
rect 6132 17466 6150 17500
rect 6034 17456 6086 17466
rect 6098 17456 6150 17466
rect 5197 17307 5249 17359
rect 6586 17806 6638 17816
rect 6586 17772 6596 17806
rect 6596 17772 6630 17806
rect 6630 17772 6638 17806
rect 6586 17764 6638 17772
rect 6820 17678 6872 17690
rect 6820 17644 6826 17678
rect 6826 17644 6860 17678
rect 6860 17644 6872 17678
rect 6820 17638 6872 17644
rect 6510 17508 6562 17560
rect 6974 17640 7026 17692
rect 7107 17220 7159 17272
rect 1398 16962 1450 16971
rect 1462 16962 1514 16971
rect 1398 16928 1417 16962
rect 1417 16928 1450 16962
rect 1462 16928 1489 16962
rect 1489 16928 1514 16962
rect 1398 16919 1450 16928
rect 1462 16919 1514 16928
rect 1526 16962 1578 16971
rect 1526 16928 1527 16962
rect 1527 16928 1561 16962
rect 1561 16928 1578 16962
rect 1526 16919 1578 16928
rect 1590 16962 1642 16971
rect 1590 16928 1599 16962
rect 1599 16928 1633 16962
rect 1633 16928 1642 16962
rect 1590 16919 1642 16928
rect 1654 16962 1706 16971
rect 1654 16928 1671 16962
rect 1671 16928 1705 16962
rect 1705 16928 1706 16962
rect 1654 16919 1706 16928
rect 1718 16962 1770 16971
rect 1782 16962 1834 16971
rect 1718 16928 1743 16962
rect 1743 16928 1770 16962
rect 1782 16928 1815 16962
rect 1815 16928 1834 16962
rect 1718 16919 1770 16928
rect 1782 16919 1834 16928
rect 560 16876 612 16900
rect 560 16848 566 16876
rect 566 16848 607 16876
rect 607 16848 612 16876
rect 702 16876 754 16896
rect 702 16844 710 16876
rect 710 16844 751 16876
rect 751 16844 754 16876
rect 378 16683 433 16738
rect 852 16694 904 16746
rect 378 16398 433 16453
rect 1004 16602 1056 16654
rect 1935 16613 1987 16665
rect 3776 16961 3828 16970
rect 3840 16961 3892 16970
rect 3904 16961 3956 16970
rect 3968 16961 4020 16970
rect 4032 16961 4084 16970
rect 4096 16961 4148 16970
rect 4160 16961 4212 16970
rect 3776 16927 3797 16961
rect 3797 16927 3828 16961
rect 3840 16927 3869 16961
rect 3869 16927 3892 16961
rect 3904 16927 3941 16961
rect 3941 16927 3956 16961
rect 3968 16927 3975 16961
rect 3975 16927 4013 16961
rect 4013 16927 4020 16961
rect 4032 16927 4047 16961
rect 4047 16927 4084 16961
rect 4096 16927 4119 16961
rect 4119 16927 4148 16961
rect 4160 16927 4191 16961
rect 4191 16927 4212 16961
rect 3776 16918 3828 16927
rect 3840 16918 3892 16927
rect 3904 16918 3956 16927
rect 3968 16918 4020 16927
rect 4032 16918 4084 16927
rect 4096 16918 4148 16927
rect 4160 16918 4212 16927
rect 2769 16804 2821 16856
rect 1155 16513 1207 16565
rect 1758 16555 1810 16564
rect 1758 16521 1773 16555
rect 1773 16521 1807 16555
rect 1807 16521 1810 16555
rect 1758 16512 1810 16521
rect 2270 16553 2322 16562
rect 2270 16519 2273 16553
rect 2273 16519 2307 16553
rect 2307 16519 2322 16553
rect 2270 16510 2322 16519
rect 3268 16727 3278 16751
rect 3278 16727 3312 16751
rect 3312 16727 3320 16751
rect 3268 16699 3320 16727
rect 4744 17018 4796 17070
rect 5029 17100 5081 17152
rect 5734 16960 5786 16970
rect 5798 16960 5850 16970
rect 5862 16960 5914 16970
rect 5926 16960 5978 16970
rect 5990 16960 6042 16970
rect 6054 16960 6106 16970
rect 6118 16960 6170 16970
rect 5734 16926 5756 16960
rect 5756 16926 5786 16960
rect 5798 16926 5828 16960
rect 5828 16926 5850 16960
rect 5862 16926 5900 16960
rect 5900 16926 5914 16960
rect 5926 16926 5934 16960
rect 5934 16926 5972 16960
rect 5972 16926 5978 16960
rect 5990 16926 6006 16960
rect 6006 16926 6042 16960
rect 6054 16926 6078 16960
rect 6078 16926 6106 16960
rect 6118 16926 6150 16960
rect 6150 16926 6170 16960
rect 5734 16918 5786 16926
rect 5798 16918 5850 16926
rect 5862 16918 5914 16926
rect 5926 16918 5978 16926
rect 5990 16918 6042 16926
rect 6054 16918 6106 16926
rect 6118 16918 6170 16926
rect 4292 16691 4344 16743
rect 5016 16690 5068 16742
rect 1248 16402 1300 16454
rect 378 16298 434 16354
rect 2020 16437 2072 16454
rect 2020 16403 2030 16437
rect 2030 16403 2064 16437
rect 2064 16403 2072 16437
rect 2020 16402 2072 16403
rect 2522 16437 2574 16452
rect 2522 16403 2530 16437
rect 2530 16403 2564 16437
rect 2564 16403 2574 16437
rect 2522 16400 2574 16403
rect 2842 16551 2894 16560
rect 2842 16517 2857 16551
rect 2857 16517 2891 16551
rect 2891 16517 2894 16551
rect 2842 16508 2894 16517
rect 3268 16506 3320 16558
rect 3561 16533 3613 16585
rect 3976 16566 4028 16576
rect 3976 16532 3984 16566
rect 3984 16532 4018 16566
rect 4018 16532 4028 16566
rect 3976 16524 4028 16532
rect 2766 16437 2818 16464
rect 2766 16412 2776 16437
rect 2776 16412 2810 16437
rect 2810 16412 2818 16437
rect 1360 16260 1412 16269
rect 1360 16226 1373 16260
rect 1373 16226 1407 16260
rect 1407 16226 1412 16260
rect 1360 16217 1412 16226
rect 1424 16260 1476 16269
rect 1488 16260 1540 16269
rect 1552 16260 1604 16269
rect 1616 16260 1668 16269
rect 1680 16260 1732 16269
rect 1744 16260 1796 16269
rect 1808 16260 1860 16269
rect 1424 16226 1445 16260
rect 1445 16226 1476 16260
rect 1488 16226 1517 16260
rect 1517 16226 1540 16260
rect 1552 16226 1589 16260
rect 1589 16226 1604 16260
rect 1616 16226 1623 16260
rect 1623 16226 1661 16260
rect 1661 16226 1668 16260
rect 1680 16226 1695 16260
rect 1695 16226 1732 16260
rect 1744 16226 1767 16260
rect 1767 16226 1796 16260
rect 1808 16226 1839 16260
rect 1839 16226 1860 16260
rect 1424 16217 1476 16226
rect 1488 16217 1540 16226
rect 1552 16217 1604 16226
rect 1616 16217 1668 16226
rect 1680 16217 1732 16226
rect 1744 16217 1796 16226
rect 1808 16217 1860 16226
rect 1872 16260 1924 16269
rect 1872 16226 1877 16260
rect 1877 16226 1911 16260
rect 1911 16226 1924 16260
rect 1872 16217 1924 16226
rect 3756 16271 3808 16280
rect 3820 16271 3872 16280
rect 278 16085 332 16139
rect 3756 16237 3775 16271
rect 3775 16237 3808 16271
rect 3820 16237 3847 16271
rect 3847 16237 3872 16271
rect 3756 16228 3808 16237
rect 3820 16228 3872 16237
rect 3884 16271 3936 16280
rect 3884 16237 3885 16271
rect 3885 16237 3919 16271
rect 3919 16237 3936 16271
rect 3884 16228 3936 16237
rect 3948 16271 4000 16280
rect 3948 16237 3957 16271
rect 3957 16237 3991 16271
rect 3991 16237 4000 16271
rect 3948 16228 4000 16237
rect 4012 16271 4064 16280
rect 4012 16237 4029 16271
rect 4029 16237 4063 16271
rect 4063 16237 4064 16271
rect 4012 16228 4064 16237
rect 4076 16271 4128 16280
rect 4140 16271 4192 16280
rect 4076 16237 4101 16271
rect 4101 16237 4128 16271
rect 4140 16237 4173 16271
rect 4173 16237 4192 16271
rect 4076 16228 4128 16237
rect 4140 16228 4192 16237
rect 3565 16079 3617 16131
rect 4628 16578 4680 16587
rect 4628 16544 4637 16578
rect 4637 16544 4671 16578
rect 4671 16544 4680 16578
rect 4628 16535 4680 16544
rect 4862 16449 4914 16462
rect 4862 16415 4868 16449
rect 4868 16415 4902 16449
rect 4902 16415 4914 16449
rect 4862 16410 4914 16415
rect 4552 16279 4604 16331
rect 6868 17018 6920 17070
rect 6250 16692 6302 16744
rect 6974 16690 7026 16742
rect 5117 16533 5169 16585
rect 5934 16566 5986 16576
rect 5934 16532 5942 16566
rect 5942 16532 5976 16566
rect 5976 16532 5986 16566
rect 5934 16524 5986 16532
rect 5015 16412 5067 16464
rect 5714 16272 5766 16280
rect 5778 16272 5830 16280
rect 5714 16238 5734 16272
rect 5734 16238 5766 16272
rect 5778 16238 5806 16272
rect 5806 16238 5830 16272
rect 5714 16228 5766 16238
rect 5778 16228 5830 16238
rect 5842 16272 5894 16280
rect 5842 16238 5844 16272
rect 5844 16238 5878 16272
rect 5878 16238 5894 16272
rect 5842 16228 5894 16238
rect 5906 16272 5958 16280
rect 5906 16238 5916 16272
rect 5916 16238 5950 16272
rect 5950 16238 5958 16272
rect 5906 16228 5958 16238
rect 5970 16272 6022 16280
rect 5970 16238 5988 16272
rect 5988 16238 6022 16272
rect 5970 16228 6022 16238
rect 6034 16272 6086 16280
rect 6098 16272 6150 16280
rect 6034 16238 6060 16272
rect 6060 16238 6086 16272
rect 6098 16238 6132 16272
rect 6132 16238 6150 16272
rect 6034 16228 6086 16238
rect 6098 16228 6150 16238
rect 5117 16079 5169 16131
rect 6586 16578 6638 16588
rect 6586 16544 6596 16578
rect 6596 16544 6630 16578
rect 6630 16544 6638 16578
rect 6586 16536 6638 16544
rect 6820 16450 6872 16462
rect 6820 16416 6826 16450
rect 6826 16416 6860 16450
rect 6860 16416 6872 16450
rect 6820 16410 6872 16416
rect 6510 16280 6562 16332
rect 6974 16412 7026 16464
rect 5035 15909 5087 15961
rect 6974 15910 7026 15962
rect 1398 15734 1450 15743
rect 1462 15734 1514 15743
rect 1398 15700 1417 15734
rect 1417 15700 1450 15734
rect 1462 15700 1489 15734
rect 1489 15700 1514 15734
rect 1398 15691 1450 15700
rect 1462 15691 1514 15700
rect 1526 15734 1578 15743
rect 1526 15700 1527 15734
rect 1527 15700 1561 15734
rect 1561 15700 1578 15734
rect 1526 15691 1578 15700
rect 1590 15734 1642 15743
rect 1590 15700 1599 15734
rect 1599 15700 1633 15734
rect 1633 15700 1642 15734
rect 1590 15691 1642 15700
rect 1654 15734 1706 15743
rect 1654 15700 1671 15734
rect 1671 15700 1705 15734
rect 1705 15700 1706 15734
rect 1654 15691 1706 15700
rect 1718 15734 1770 15743
rect 1782 15734 1834 15743
rect 1718 15700 1743 15734
rect 1743 15700 1770 15734
rect 1782 15700 1815 15734
rect 1815 15700 1834 15734
rect 1718 15691 1770 15700
rect 1782 15691 1834 15700
rect 560 15648 612 15672
rect 560 15620 566 15648
rect 566 15620 607 15648
rect 607 15620 612 15648
rect 702 15648 754 15668
rect 702 15616 710 15648
rect 710 15616 751 15648
rect 751 15616 754 15648
rect 378 15455 433 15510
rect 852 15466 904 15518
rect 378 15170 433 15225
rect 1004 15374 1056 15426
rect 1935 15385 1987 15437
rect 3776 15733 3828 15742
rect 3840 15733 3892 15742
rect 3904 15733 3956 15742
rect 3968 15733 4020 15742
rect 4032 15733 4084 15742
rect 4096 15733 4148 15742
rect 4160 15733 4212 15742
rect 3776 15699 3797 15733
rect 3797 15699 3828 15733
rect 3840 15699 3869 15733
rect 3869 15699 3892 15733
rect 3904 15699 3941 15733
rect 3941 15699 3956 15733
rect 3968 15699 3975 15733
rect 3975 15699 4013 15733
rect 4013 15699 4020 15733
rect 4032 15699 4047 15733
rect 4047 15699 4084 15733
rect 4096 15699 4119 15733
rect 4119 15699 4148 15733
rect 4160 15699 4191 15733
rect 4191 15699 4212 15733
rect 3776 15690 3828 15699
rect 3840 15690 3892 15699
rect 3904 15690 3956 15699
rect 3968 15690 4020 15699
rect 4032 15690 4084 15699
rect 4096 15690 4148 15699
rect 4160 15690 4212 15699
rect 2769 15576 2821 15628
rect 1155 15285 1207 15337
rect 1758 15327 1810 15336
rect 1758 15293 1773 15327
rect 1773 15293 1807 15327
rect 1807 15293 1810 15327
rect 1758 15284 1810 15293
rect 2270 15325 2322 15334
rect 2270 15291 2273 15325
rect 2273 15291 2307 15325
rect 2307 15291 2322 15325
rect 2270 15282 2322 15291
rect 3268 15499 3278 15523
rect 3278 15499 3312 15523
rect 3312 15499 3320 15523
rect 3268 15471 3320 15499
rect 4744 15790 4796 15842
rect 5734 15732 5786 15742
rect 5798 15732 5850 15742
rect 5862 15732 5914 15742
rect 5926 15732 5978 15742
rect 5990 15732 6042 15742
rect 6054 15732 6106 15742
rect 6118 15732 6170 15742
rect 5734 15698 5756 15732
rect 5756 15698 5786 15732
rect 5798 15698 5828 15732
rect 5828 15698 5850 15732
rect 5862 15698 5900 15732
rect 5900 15698 5914 15732
rect 5926 15698 5934 15732
rect 5934 15698 5972 15732
rect 5972 15698 5978 15732
rect 5990 15698 6006 15732
rect 6006 15698 6042 15732
rect 6054 15698 6078 15732
rect 6078 15698 6106 15732
rect 6118 15698 6150 15732
rect 6150 15698 6170 15732
rect 5734 15690 5786 15698
rect 5798 15690 5850 15698
rect 5862 15690 5914 15698
rect 5926 15690 5978 15698
rect 5990 15690 6042 15698
rect 6054 15690 6106 15698
rect 6118 15690 6170 15698
rect 4292 15463 4344 15515
rect 5016 15462 5068 15514
rect 1248 15174 1300 15226
rect 378 15070 434 15126
rect 2020 15209 2072 15226
rect 2020 15175 2030 15209
rect 2030 15175 2064 15209
rect 2064 15175 2072 15209
rect 2020 15174 2072 15175
rect 2522 15209 2574 15224
rect 2522 15175 2530 15209
rect 2530 15175 2564 15209
rect 2564 15175 2574 15209
rect 2522 15172 2574 15175
rect 2842 15323 2894 15332
rect 2842 15289 2857 15323
rect 2857 15289 2891 15323
rect 2891 15289 2894 15323
rect 2842 15280 2894 15289
rect 3268 15278 3320 15330
rect 3561 15305 3613 15357
rect 3976 15338 4028 15348
rect 3976 15304 3984 15338
rect 3984 15304 4018 15338
rect 4018 15304 4028 15338
rect 3976 15296 4028 15304
rect 2766 15209 2818 15236
rect 2766 15184 2776 15209
rect 2776 15184 2810 15209
rect 2810 15184 2818 15209
rect 1360 15032 1412 15041
rect 1360 14998 1373 15032
rect 1373 14998 1407 15032
rect 1407 14998 1412 15032
rect 1360 14989 1412 14998
rect 1424 15032 1476 15041
rect 1488 15032 1540 15041
rect 1552 15032 1604 15041
rect 1616 15032 1668 15041
rect 1680 15032 1732 15041
rect 1744 15032 1796 15041
rect 1808 15032 1860 15041
rect 1424 14998 1445 15032
rect 1445 14998 1476 15032
rect 1488 14998 1517 15032
rect 1517 14998 1540 15032
rect 1552 14998 1589 15032
rect 1589 14998 1604 15032
rect 1616 14998 1623 15032
rect 1623 14998 1661 15032
rect 1661 14998 1668 15032
rect 1680 14998 1695 15032
rect 1695 14998 1732 15032
rect 1744 14998 1767 15032
rect 1767 14998 1796 15032
rect 1808 14998 1839 15032
rect 1839 14998 1860 15032
rect 1424 14989 1476 14998
rect 1488 14989 1540 14998
rect 1552 14989 1604 14998
rect 1616 14989 1668 14998
rect 1680 14989 1732 14998
rect 1744 14989 1796 14998
rect 1808 14989 1860 14998
rect 1872 15032 1924 15041
rect 1872 14998 1877 15032
rect 1877 14998 1911 15032
rect 1911 14998 1924 15032
rect 1872 14989 1924 14998
rect 3756 15043 3808 15052
rect 3820 15043 3872 15052
rect 278 14857 332 14911
rect 3756 15009 3775 15043
rect 3775 15009 3808 15043
rect 3820 15009 3847 15043
rect 3847 15009 3872 15043
rect 3756 15000 3808 15009
rect 3820 15000 3872 15009
rect 3884 15043 3936 15052
rect 3884 15009 3885 15043
rect 3885 15009 3919 15043
rect 3919 15009 3936 15043
rect 3884 15000 3936 15009
rect 3948 15043 4000 15052
rect 3948 15009 3957 15043
rect 3957 15009 3991 15043
rect 3991 15009 4000 15043
rect 3948 15000 4000 15009
rect 4012 15043 4064 15052
rect 4012 15009 4029 15043
rect 4029 15009 4063 15043
rect 4063 15009 4064 15043
rect 4012 15000 4064 15009
rect 4076 15043 4128 15052
rect 4140 15043 4192 15052
rect 4076 15009 4101 15043
rect 4101 15009 4128 15043
rect 4140 15009 4173 15043
rect 4173 15009 4192 15043
rect 4076 15000 4128 15009
rect 4140 15000 4192 15009
rect 3565 14851 3617 14903
rect 4628 15350 4680 15359
rect 4628 15316 4637 15350
rect 4637 15316 4671 15350
rect 4671 15316 4680 15350
rect 4628 15307 4680 15316
rect 4862 15221 4914 15234
rect 4862 15187 4868 15221
rect 4868 15187 4902 15221
rect 4902 15187 4914 15221
rect 4862 15182 4914 15187
rect 4552 15051 4604 15103
rect 6250 15464 6302 15516
rect 6974 15462 7026 15514
rect 5279 15305 5331 15357
rect 5934 15338 5986 15348
rect 5934 15304 5942 15338
rect 5942 15304 5976 15338
rect 5976 15304 5986 15338
rect 5934 15296 5986 15304
rect 5015 15184 5067 15236
rect 5714 15044 5766 15052
rect 5778 15044 5830 15052
rect 5714 15010 5734 15044
rect 5734 15010 5766 15044
rect 5778 15010 5806 15044
rect 5806 15010 5830 15044
rect 5714 15000 5766 15010
rect 5778 15000 5830 15010
rect 5842 15044 5894 15052
rect 5842 15010 5844 15044
rect 5844 15010 5878 15044
rect 5878 15010 5894 15044
rect 5842 15000 5894 15010
rect 5906 15044 5958 15052
rect 5906 15010 5916 15044
rect 5916 15010 5950 15044
rect 5950 15010 5958 15044
rect 5906 15000 5958 15010
rect 5970 15044 6022 15052
rect 5970 15010 5988 15044
rect 5988 15010 6022 15044
rect 5970 15000 6022 15010
rect 6034 15044 6086 15052
rect 6098 15044 6150 15052
rect 6034 15010 6060 15044
rect 6060 15010 6086 15044
rect 6098 15010 6132 15044
rect 6132 15010 6150 15044
rect 6034 15000 6086 15010
rect 6098 15000 6150 15010
rect 5279 14851 5331 14903
rect 6586 15350 6638 15360
rect 6586 15316 6596 15350
rect 6596 15316 6630 15350
rect 6630 15316 6638 15350
rect 6586 15308 6638 15316
rect 6820 15222 6872 15234
rect 6820 15188 6826 15222
rect 6826 15188 6860 15222
rect 6860 15188 6872 15222
rect 6820 15182 6872 15188
rect 6510 15052 6562 15104
rect 6974 15184 7026 15236
rect 1398 14506 1450 14515
rect 1462 14506 1514 14515
rect 1398 14472 1417 14506
rect 1417 14472 1450 14506
rect 1462 14472 1489 14506
rect 1489 14472 1514 14506
rect 1398 14463 1450 14472
rect 1462 14463 1514 14472
rect 1526 14506 1578 14515
rect 1526 14472 1527 14506
rect 1527 14472 1561 14506
rect 1561 14472 1578 14506
rect 1526 14463 1578 14472
rect 1590 14506 1642 14515
rect 1590 14472 1599 14506
rect 1599 14472 1633 14506
rect 1633 14472 1642 14506
rect 1590 14463 1642 14472
rect 1654 14506 1706 14515
rect 1654 14472 1671 14506
rect 1671 14472 1705 14506
rect 1705 14472 1706 14506
rect 1654 14463 1706 14472
rect 1718 14506 1770 14515
rect 1782 14506 1834 14515
rect 1718 14472 1743 14506
rect 1743 14472 1770 14506
rect 1782 14472 1815 14506
rect 1815 14472 1834 14506
rect 1718 14463 1770 14472
rect 1782 14463 1834 14472
rect 560 14420 612 14444
rect 560 14392 566 14420
rect 566 14392 607 14420
rect 607 14392 612 14420
rect 702 14420 754 14440
rect 702 14388 710 14420
rect 710 14388 751 14420
rect 751 14388 754 14420
rect 378 14227 433 14282
rect 852 14238 904 14290
rect 378 13942 433 13997
rect 1004 14146 1056 14198
rect 1935 14157 1987 14209
rect 3776 14505 3828 14514
rect 3840 14505 3892 14514
rect 3904 14505 3956 14514
rect 3968 14505 4020 14514
rect 4032 14505 4084 14514
rect 4096 14505 4148 14514
rect 4160 14505 4212 14514
rect 3776 14471 3797 14505
rect 3797 14471 3828 14505
rect 3840 14471 3869 14505
rect 3869 14471 3892 14505
rect 3904 14471 3941 14505
rect 3941 14471 3956 14505
rect 3968 14471 3975 14505
rect 3975 14471 4013 14505
rect 4013 14471 4020 14505
rect 4032 14471 4047 14505
rect 4047 14471 4084 14505
rect 4096 14471 4119 14505
rect 4119 14471 4148 14505
rect 4160 14471 4191 14505
rect 4191 14471 4212 14505
rect 3776 14462 3828 14471
rect 3840 14462 3892 14471
rect 3904 14462 3956 14471
rect 3968 14462 4020 14471
rect 4032 14462 4084 14471
rect 4096 14462 4148 14471
rect 4160 14462 4212 14471
rect 2769 14348 2821 14400
rect 1155 14057 1207 14109
rect 1758 14099 1810 14108
rect 1758 14065 1773 14099
rect 1773 14065 1807 14099
rect 1807 14065 1810 14099
rect 1758 14056 1810 14065
rect 2270 14097 2322 14106
rect 2270 14063 2273 14097
rect 2273 14063 2307 14097
rect 2307 14063 2322 14097
rect 2270 14054 2322 14063
rect 3268 14271 3278 14295
rect 3278 14271 3312 14295
rect 3312 14271 3320 14295
rect 3268 14243 3320 14271
rect 4744 14562 4796 14614
rect 5029 14644 5081 14696
rect 5734 14504 5786 14514
rect 5798 14504 5850 14514
rect 5862 14504 5914 14514
rect 5926 14504 5978 14514
rect 5990 14504 6042 14514
rect 6054 14504 6106 14514
rect 6118 14504 6170 14514
rect 5734 14470 5756 14504
rect 5756 14470 5786 14504
rect 5798 14470 5828 14504
rect 5828 14470 5850 14504
rect 5862 14470 5900 14504
rect 5900 14470 5914 14504
rect 5926 14470 5934 14504
rect 5934 14470 5972 14504
rect 5972 14470 5978 14504
rect 5990 14470 6006 14504
rect 6006 14470 6042 14504
rect 6054 14470 6078 14504
rect 6078 14470 6106 14504
rect 6118 14470 6150 14504
rect 6150 14470 6170 14504
rect 5734 14462 5786 14470
rect 5798 14462 5850 14470
rect 5862 14462 5914 14470
rect 5926 14462 5978 14470
rect 5990 14462 6042 14470
rect 6054 14462 6106 14470
rect 6118 14462 6170 14470
rect 4292 14235 4344 14287
rect 5016 14234 5068 14286
rect 1248 13946 1300 13998
rect 378 13842 434 13898
rect 2020 13981 2072 13998
rect 2020 13947 2030 13981
rect 2030 13947 2064 13981
rect 2064 13947 2072 13981
rect 2020 13946 2072 13947
rect 2522 13981 2574 13996
rect 2522 13947 2530 13981
rect 2530 13947 2564 13981
rect 2564 13947 2574 13981
rect 2522 13944 2574 13947
rect 2842 14095 2894 14104
rect 2842 14061 2857 14095
rect 2857 14061 2891 14095
rect 2891 14061 2894 14095
rect 2842 14052 2894 14061
rect 3268 14050 3320 14102
rect 3561 14077 3613 14129
rect 3976 14110 4028 14120
rect 3976 14076 3984 14110
rect 3984 14076 4018 14110
rect 4018 14076 4028 14110
rect 3976 14068 4028 14076
rect 2766 13981 2818 14008
rect 2766 13956 2776 13981
rect 2776 13956 2810 13981
rect 2810 13956 2818 13981
rect 1360 13804 1412 13813
rect 1360 13770 1373 13804
rect 1373 13770 1407 13804
rect 1407 13770 1412 13804
rect 1360 13761 1412 13770
rect 1424 13804 1476 13813
rect 1488 13804 1540 13813
rect 1552 13804 1604 13813
rect 1616 13804 1668 13813
rect 1680 13804 1732 13813
rect 1744 13804 1796 13813
rect 1808 13804 1860 13813
rect 1424 13770 1445 13804
rect 1445 13770 1476 13804
rect 1488 13770 1517 13804
rect 1517 13770 1540 13804
rect 1552 13770 1589 13804
rect 1589 13770 1604 13804
rect 1616 13770 1623 13804
rect 1623 13770 1661 13804
rect 1661 13770 1668 13804
rect 1680 13770 1695 13804
rect 1695 13770 1732 13804
rect 1744 13770 1767 13804
rect 1767 13770 1796 13804
rect 1808 13770 1839 13804
rect 1839 13770 1860 13804
rect 1424 13761 1476 13770
rect 1488 13761 1540 13770
rect 1552 13761 1604 13770
rect 1616 13761 1668 13770
rect 1680 13761 1732 13770
rect 1744 13761 1796 13770
rect 1808 13761 1860 13770
rect 1872 13804 1924 13813
rect 1872 13770 1877 13804
rect 1877 13770 1911 13804
rect 1911 13770 1924 13804
rect 1872 13761 1924 13770
rect 3756 13815 3808 13824
rect 3820 13815 3872 13824
rect 278 13629 332 13683
rect 3756 13781 3775 13815
rect 3775 13781 3808 13815
rect 3820 13781 3847 13815
rect 3847 13781 3872 13815
rect 3756 13772 3808 13781
rect 3820 13772 3872 13781
rect 3884 13815 3936 13824
rect 3884 13781 3885 13815
rect 3885 13781 3919 13815
rect 3919 13781 3936 13815
rect 3884 13772 3936 13781
rect 3948 13815 4000 13824
rect 3948 13781 3957 13815
rect 3957 13781 3991 13815
rect 3991 13781 4000 13815
rect 3948 13772 4000 13781
rect 4012 13815 4064 13824
rect 4012 13781 4029 13815
rect 4029 13781 4063 13815
rect 4063 13781 4064 13815
rect 4012 13772 4064 13781
rect 4076 13815 4128 13824
rect 4140 13815 4192 13824
rect 4076 13781 4101 13815
rect 4101 13781 4128 13815
rect 4140 13781 4173 13815
rect 4173 13781 4192 13815
rect 4076 13772 4128 13781
rect 4140 13772 4192 13781
rect 3565 13623 3617 13675
rect 4628 14122 4680 14131
rect 4628 14088 4637 14122
rect 4637 14088 4671 14122
rect 4671 14088 4680 14122
rect 4628 14079 4680 14088
rect 4862 13993 4914 14006
rect 4862 13959 4868 13993
rect 4868 13959 4902 13993
rect 4902 13959 4914 13993
rect 4862 13954 4914 13959
rect 4552 13823 4604 13875
rect 6868 14562 6920 14614
rect 6250 14236 6302 14288
rect 7194 14444 7246 14496
rect 6974 14234 7026 14286
rect 5117 14077 5169 14129
rect 5934 14110 5986 14120
rect 5934 14076 5942 14110
rect 5942 14076 5976 14110
rect 5976 14076 5986 14110
rect 5934 14068 5986 14076
rect 5015 13956 5067 14008
rect 5714 13816 5766 13824
rect 5778 13816 5830 13824
rect 5714 13782 5734 13816
rect 5734 13782 5766 13816
rect 5778 13782 5806 13816
rect 5806 13782 5830 13816
rect 5714 13772 5766 13782
rect 5778 13772 5830 13782
rect 5842 13816 5894 13824
rect 5842 13782 5844 13816
rect 5844 13782 5878 13816
rect 5878 13782 5894 13816
rect 5842 13772 5894 13782
rect 5906 13816 5958 13824
rect 5906 13782 5916 13816
rect 5916 13782 5950 13816
rect 5950 13782 5958 13816
rect 5906 13772 5958 13782
rect 5970 13816 6022 13824
rect 5970 13782 5988 13816
rect 5988 13782 6022 13816
rect 5970 13772 6022 13782
rect 6034 13816 6086 13824
rect 6098 13816 6150 13824
rect 6034 13782 6060 13816
rect 6060 13782 6086 13816
rect 6098 13782 6132 13816
rect 6132 13782 6150 13816
rect 6034 13772 6086 13782
rect 6098 13772 6150 13782
rect 5117 13623 5169 13675
rect 6586 14122 6638 14132
rect 6586 14088 6596 14122
rect 6596 14088 6630 14122
rect 6630 14088 6638 14122
rect 6586 14080 6638 14088
rect 6820 13994 6872 14006
rect 6820 13960 6826 13994
rect 6826 13960 6860 13994
rect 6860 13960 6872 13994
rect 6820 13954 6872 13960
rect 6510 13824 6562 13876
rect 6974 13956 7026 14008
rect 5035 13453 5087 13505
rect 6512 13538 6564 13590
rect 1398 13278 1450 13287
rect 1462 13278 1514 13287
rect 1398 13244 1417 13278
rect 1417 13244 1450 13278
rect 1462 13244 1489 13278
rect 1489 13244 1514 13278
rect 1398 13235 1450 13244
rect 1462 13235 1514 13244
rect 1526 13278 1578 13287
rect 1526 13244 1527 13278
rect 1527 13244 1561 13278
rect 1561 13244 1578 13278
rect 1526 13235 1578 13244
rect 1590 13278 1642 13287
rect 1590 13244 1599 13278
rect 1599 13244 1633 13278
rect 1633 13244 1642 13278
rect 1590 13235 1642 13244
rect 1654 13278 1706 13287
rect 1654 13244 1671 13278
rect 1671 13244 1705 13278
rect 1705 13244 1706 13278
rect 1654 13235 1706 13244
rect 1718 13278 1770 13287
rect 1782 13278 1834 13287
rect 1718 13244 1743 13278
rect 1743 13244 1770 13278
rect 1782 13244 1815 13278
rect 1815 13244 1834 13278
rect 1718 13235 1770 13244
rect 1782 13235 1834 13244
rect 560 13192 612 13216
rect 560 13164 566 13192
rect 566 13164 607 13192
rect 607 13164 612 13192
rect 702 13192 754 13212
rect 702 13160 710 13192
rect 710 13160 751 13192
rect 751 13160 754 13192
rect 378 12999 433 13054
rect 852 13010 904 13062
rect 378 12714 433 12769
rect 1004 12918 1056 12970
rect 1935 12929 1987 12981
rect 3776 13277 3828 13286
rect 3840 13277 3892 13286
rect 3904 13277 3956 13286
rect 3968 13277 4020 13286
rect 4032 13277 4084 13286
rect 4096 13277 4148 13286
rect 4160 13277 4212 13286
rect 3776 13243 3797 13277
rect 3797 13243 3828 13277
rect 3840 13243 3869 13277
rect 3869 13243 3892 13277
rect 3904 13243 3941 13277
rect 3941 13243 3956 13277
rect 3968 13243 3975 13277
rect 3975 13243 4013 13277
rect 4013 13243 4020 13277
rect 4032 13243 4047 13277
rect 4047 13243 4084 13277
rect 4096 13243 4119 13277
rect 4119 13243 4148 13277
rect 4160 13243 4191 13277
rect 4191 13243 4212 13277
rect 3776 13234 3828 13243
rect 3840 13234 3892 13243
rect 3904 13234 3956 13243
rect 3968 13234 4020 13243
rect 4032 13234 4084 13243
rect 4096 13234 4148 13243
rect 4160 13234 4212 13243
rect 2769 13120 2821 13172
rect 1155 12829 1207 12881
rect 1758 12871 1810 12880
rect 1758 12837 1773 12871
rect 1773 12837 1807 12871
rect 1807 12837 1810 12871
rect 1758 12828 1810 12837
rect 2270 12869 2322 12878
rect 2270 12835 2273 12869
rect 2273 12835 2307 12869
rect 2307 12835 2322 12869
rect 2270 12826 2322 12835
rect 3268 13043 3278 13067
rect 3278 13043 3312 13067
rect 3312 13043 3320 13067
rect 3268 13015 3320 13043
rect 4744 13334 4796 13386
rect 5734 13276 5786 13286
rect 5798 13276 5850 13286
rect 5862 13276 5914 13286
rect 5926 13276 5978 13286
rect 5990 13276 6042 13286
rect 6054 13276 6106 13286
rect 6118 13276 6170 13286
rect 5734 13242 5756 13276
rect 5756 13242 5786 13276
rect 5798 13242 5828 13276
rect 5828 13242 5850 13276
rect 5862 13242 5900 13276
rect 5900 13242 5914 13276
rect 5926 13242 5934 13276
rect 5934 13242 5972 13276
rect 5972 13242 5978 13276
rect 5990 13242 6006 13276
rect 6006 13242 6042 13276
rect 6054 13242 6078 13276
rect 6078 13242 6106 13276
rect 6118 13242 6150 13276
rect 6150 13242 6170 13276
rect 5734 13234 5786 13242
rect 5798 13234 5850 13242
rect 5862 13234 5914 13242
rect 5926 13234 5978 13242
rect 5990 13234 6042 13242
rect 6054 13234 6106 13242
rect 6118 13234 6170 13242
rect 4292 13007 4344 13059
rect 5016 13006 5068 13058
rect 1248 12718 1300 12770
rect 378 12614 434 12670
rect 2020 12753 2072 12770
rect 2020 12719 2030 12753
rect 2030 12719 2064 12753
rect 2064 12719 2072 12753
rect 2020 12718 2072 12719
rect 2522 12753 2574 12768
rect 2522 12719 2530 12753
rect 2530 12719 2564 12753
rect 2564 12719 2574 12753
rect 2522 12716 2574 12719
rect 2842 12867 2894 12876
rect 2842 12833 2857 12867
rect 2857 12833 2891 12867
rect 2891 12833 2894 12867
rect 2842 12824 2894 12833
rect 3268 12822 3320 12874
rect 3561 12849 3613 12901
rect 3976 12882 4028 12892
rect 3976 12848 3984 12882
rect 3984 12848 4018 12882
rect 4018 12848 4028 12882
rect 3976 12840 4028 12848
rect 2766 12753 2818 12780
rect 2766 12728 2776 12753
rect 2776 12728 2810 12753
rect 2810 12728 2818 12753
rect 1360 12576 1412 12585
rect 1360 12542 1373 12576
rect 1373 12542 1407 12576
rect 1407 12542 1412 12576
rect 1360 12533 1412 12542
rect 1424 12576 1476 12585
rect 1488 12576 1540 12585
rect 1552 12576 1604 12585
rect 1616 12576 1668 12585
rect 1680 12576 1732 12585
rect 1744 12576 1796 12585
rect 1808 12576 1860 12585
rect 1424 12542 1445 12576
rect 1445 12542 1476 12576
rect 1488 12542 1517 12576
rect 1517 12542 1540 12576
rect 1552 12542 1589 12576
rect 1589 12542 1604 12576
rect 1616 12542 1623 12576
rect 1623 12542 1661 12576
rect 1661 12542 1668 12576
rect 1680 12542 1695 12576
rect 1695 12542 1732 12576
rect 1744 12542 1767 12576
rect 1767 12542 1796 12576
rect 1808 12542 1839 12576
rect 1839 12542 1860 12576
rect 1424 12533 1476 12542
rect 1488 12533 1540 12542
rect 1552 12533 1604 12542
rect 1616 12533 1668 12542
rect 1680 12533 1732 12542
rect 1744 12533 1796 12542
rect 1808 12533 1860 12542
rect 1872 12576 1924 12585
rect 1872 12542 1877 12576
rect 1877 12542 1911 12576
rect 1911 12542 1924 12576
rect 1872 12533 1924 12542
rect 3756 12587 3808 12596
rect 3820 12587 3872 12596
rect 278 12401 332 12455
rect 3756 12553 3775 12587
rect 3775 12553 3808 12587
rect 3820 12553 3847 12587
rect 3847 12553 3872 12587
rect 3756 12544 3808 12553
rect 3820 12544 3872 12553
rect 3884 12587 3936 12596
rect 3884 12553 3885 12587
rect 3885 12553 3919 12587
rect 3919 12553 3936 12587
rect 3884 12544 3936 12553
rect 3948 12587 4000 12596
rect 3948 12553 3957 12587
rect 3957 12553 3991 12587
rect 3991 12553 4000 12587
rect 3948 12544 4000 12553
rect 4012 12587 4064 12596
rect 4012 12553 4029 12587
rect 4029 12553 4063 12587
rect 4063 12553 4064 12587
rect 4012 12544 4064 12553
rect 4076 12587 4128 12596
rect 4140 12587 4192 12596
rect 4076 12553 4101 12587
rect 4101 12553 4128 12587
rect 4140 12553 4173 12587
rect 4173 12553 4192 12587
rect 4076 12544 4128 12553
rect 4140 12544 4192 12553
rect 3565 12395 3617 12447
rect 4628 12894 4680 12903
rect 4628 12860 4637 12894
rect 4637 12860 4671 12894
rect 4671 12860 4680 12894
rect 4628 12851 4680 12860
rect 4862 12765 4914 12778
rect 4862 12731 4868 12765
rect 4868 12731 4902 12765
rect 4902 12731 4914 12765
rect 4862 12726 4914 12731
rect 4552 12595 4604 12647
rect 6843 13334 6895 13386
rect 6250 13008 6302 13060
rect 6974 13006 7026 13058
rect 5197 12849 5249 12901
rect 5934 12882 5986 12892
rect 5934 12848 5942 12882
rect 5942 12848 5976 12882
rect 5976 12848 5986 12882
rect 5934 12840 5986 12848
rect 5015 12728 5067 12780
rect 5714 12588 5766 12596
rect 5778 12588 5830 12596
rect 5714 12554 5734 12588
rect 5734 12554 5766 12588
rect 5778 12554 5806 12588
rect 5806 12554 5830 12588
rect 5714 12544 5766 12554
rect 5778 12544 5830 12554
rect 5842 12588 5894 12596
rect 5842 12554 5844 12588
rect 5844 12554 5878 12588
rect 5878 12554 5894 12588
rect 5842 12544 5894 12554
rect 5906 12588 5958 12596
rect 5906 12554 5916 12588
rect 5916 12554 5950 12588
rect 5950 12554 5958 12588
rect 5906 12544 5958 12554
rect 5970 12588 6022 12596
rect 5970 12554 5988 12588
rect 5988 12554 6022 12588
rect 5970 12544 6022 12554
rect 6034 12588 6086 12596
rect 6098 12588 6150 12596
rect 6034 12554 6060 12588
rect 6060 12554 6086 12588
rect 6098 12554 6132 12588
rect 6132 12554 6150 12588
rect 6034 12544 6086 12554
rect 6098 12544 6150 12554
rect 5197 12395 5249 12447
rect 6586 12894 6638 12904
rect 6586 12860 6596 12894
rect 6596 12860 6630 12894
rect 6630 12860 6638 12894
rect 6586 12852 6638 12860
rect 6820 12766 6872 12778
rect 6820 12732 6826 12766
rect 6826 12732 6860 12766
rect 6860 12732 6872 12766
rect 6820 12726 6872 12732
rect 6510 12596 6562 12648
rect 6974 12728 7026 12780
rect 7107 12308 7159 12360
rect 1398 12050 1450 12059
rect 1462 12050 1514 12059
rect 1398 12016 1417 12050
rect 1417 12016 1450 12050
rect 1462 12016 1489 12050
rect 1489 12016 1514 12050
rect 1398 12007 1450 12016
rect 1462 12007 1514 12016
rect 1526 12050 1578 12059
rect 1526 12016 1527 12050
rect 1527 12016 1561 12050
rect 1561 12016 1578 12050
rect 1526 12007 1578 12016
rect 1590 12050 1642 12059
rect 1590 12016 1599 12050
rect 1599 12016 1633 12050
rect 1633 12016 1642 12050
rect 1590 12007 1642 12016
rect 1654 12050 1706 12059
rect 1654 12016 1671 12050
rect 1671 12016 1705 12050
rect 1705 12016 1706 12050
rect 1654 12007 1706 12016
rect 1718 12050 1770 12059
rect 1782 12050 1834 12059
rect 1718 12016 1743 12050
rect 1743 12016 1770 12050
rect 1782 12016 1815 12050
rect 1815 12016 1834 12050
rect 1718 12007 1770 12016
rect 1782 12007 1834 12016
rect 560 11964 612 11988
rect 560 11936 566 11964
rect 566 11936 607 11964
rect 607 11936 612 11964
rect 702 11964 754 11984
rect 702 11932 710 11964
rect 710 11932 751 11964
rect 751 11932 754 11964
rect 378 11771 433 11826
rect 852 11782 904 11834
rect 378 11486 433 11541
rect 1004 11690 1056 11742
rect 1935 11701 1987 11753
rect 3776 12049 3828 12058
rect 3840 12049 3892 12058
rect 3904 12049 3956 12058
rect 3968 12049 4020 12058
rect 4032 12049 4084 12058
rect 4096 12049 4148 12058
rect 4160 12049 4212 12058
rect 3776 12015 3797 12049
rect 3797 12015 3828 12049
rect 3840 12015 3869 12049
rect 3869 12015 3892 12049
rect 3904 12015 3941 12049
rect 3941 12015 3956 12049
rect 3968 12015 3975 12049
rect 3975 12015 4013 12049
rect 4013 12015 4020 12049
rect 4032 12015 4047 12049
rect 4047 12015 4084 12049
rect 4096 12015 4119 12049
rect 4119 12015 4148 12049
rect 4160 12015 4191 12049
rect 4191 12015 4212 12049
rect 3776 12006 3828 12015
rect 3840 12006 3892 12015
rect 3904 12006 3956 12015
rect 3968 12006 4020 12015
rect 4032 12006 4084 12015
rect 4096 12006 4148 12015
rect 4160 12006 4212 12015
rect 2769 11892 2821 11944
rect 1155 11601 1207 11653
rect 1758 11643 1810 11652
rect 1758 11609 1773 11643
rect 1773 11609 1807 11643
rect 1807 11609 1810 11643
rect 1758 11600 1810 11609
rect 2270 11641 2322 11650
rect 2270 11607 2273 11641
rect 2273 11607 2307 11641
rect 2307 11607 2322 11641
rect 2270 11598 2322 11607
rect 3268 11815 3278 11839
rect 3278 11815 3312 11839
rect 3312 11815 3320 11839
rect 3268 11787 3320 11815
rect 4744 12106 4796 12158
rect 5029 12188 5081 12240
rect 5734 12048 5786 12058
rect 5798 12048 5850 12058
rect 5862 12048 5914 12058
rect 5926 12048 5978 12058
rect 5990 12048 6042 12058
rect 6054 12048 6106 12058
rect 6118 12048 6170 12058
rect 5734 12014 5756 12048
rect 5756 12014 5786 12048
rect 5798 12014 5828 12048
rect 5828 12014 5850 12048
rect 5862 12014 5900 12048
rect 5900 12014 5914 12048
rect 5926 12014 5934 12048
rect 5934 12014 5972 12048
rect 5972 12014 5978 12048
rect 5990 12014 6006 12048
rect 6006 12014 6042 12048
rect 6054 12014 6078 12048
rect 6078 12014 6106 12048
rect 6118 12014 6150 12048
rect 6150 12014 6170 12048
rect 5734 12006 5786 12014
rect 5798 12006 5850 12014
rect 5862 12006 5914 12014
rect 5926 12006 5978 12014
rect 5990 12006 6042 12014
rect 6054 12006 6106 12014
rect 6118 12006 6170 12014
rect 4292 11779 4344 11831
rect 5016 11778 5068 11830
rect 1248 11490 1300 11542
rect 378 11386 434 11442
rect 2020 11525 2072 11542
rect 2020 11491 2030 11525
rect 2030 11491 2064 11525
rect 2064 11491 2072 11525
rect 2020 11490 2072 11491
rect 2522 11525 2574 11540
rect 2522 11491 2530 11525
rect 2530 11491 2564 11525
rect 2564 11491 2574 11525
rect 2522 11488 2574 11491
rect 2842 11639 2894 11648
rect 2842 11605 2857 11639
rect 2857 11605 2891 11639
rect 2891 11605 2894 11639
rect 2842 11596 2894 11605
rect 3268 11594 3320 11646
rect 3561 11621 3613 11673
rect 3976 11654 4028 11664
rect 3976 11620 3984 11654
rect 3984 11620 4018 11654
rect 4018 11620 4028 11654
rect 3976 11612 4028 11620
rect 2766 11525 2818 11552
rect 2766 11500 2776 11525
rect 2776 11500 2810 11525
rect 2810 11500 2818 11525
rect 1360 11348 1412 11357
rect 1360 11314 1373 11348
rect 1373 11314 1407 11348
rect 1407 11314 1412 11348
rect 1360 11305 1412 11314
rect 1424 11348 1476 11357
rect 1488 11348 1540 11357
rect 1552 11348 1604 11357
rect 1616 11348 1668 11357
rect 1680 11348 1732 11357
rect 1744 11348 1796 11357
rect 1808 11348 1860 11357
rect 1424 11314 1445 11348
rect 1445 11314 1476 11348
rect 1488 11314 1517 11348
rect 1517 11314 1540 11348
rect 1552 11314 1589 11348
rect 1589 11314 1604 11348
rect 1616 11314 1623 11348
rect 1623 11314 1661 11348
rect 1661 11314 1668 11348
rect 1680 11314 1695 11348
rect 1695 11314 1732 11348
rect 1744 11314 1767 11348
rect 1767 11314 1796 11348
rect 1808 11314 1839 11348
rect 1839 11314 1860 11348
rect 1424 11305 1476 11314
rect 1488 11305 1540 11314
rect 1552 11305 1604 11314
rect 1616 11305 1668 11314
rect 1680 11305 1732 11314
rect 1744 11305 1796 11314
rect 1808 11305 1860 11314
rect 1872 11348 1924 11357
rect 1872 11314 1877 11348
rect 1877 11314 1911 11348
rect 1911 11314 1924 11348
rect 1872 11305 1924 11314
rect 3756 11359 3808 11368
rect 3820 11359 3872 11368
rect 278 11173 332 11227
rect 3756 11325 3775 11359
rect 3775 11325 3808 11359
rect 3820 11325 3847 11359
rect 3847 11325 3872 11359
rect 3756 11316 3808 11325
rect 3820 11316 3872 11325
rect 3884 11359 3936 11368
rect 3884 11325 3885 11359
rect 3885 11325 3919 11359
rect 3919 11325 3936 11359
rect 3884 11316 3936 11325
rect 3948 11359 4000 11368
rect 3948 11325 3957 11359
rect 3957 11325 3991 11359
rect 3991 11325 4000 11359
rect 3948 11316 4000 11325
rect 4012 11359 4064 11368
rect 4012 11325 4029 11359
rect 4029 11325 4063 11359
rect 4063 11325 4064 11359
rect 4012 11316 4064 11325
rect 4076 11359 4128 11368
rect 4140 11359 4192 11368
rect 4076 11325 4101 11359
rect 4101 11325 4128 11359
rect 4140 11325 4173 11359
rect 4173 11325 4192 11359
rect 4076 11316 4128 11325
rect 4140 11316 4192 11325
rect 3565 11167 3617 11219
rect 4628 11666 4680 11675
rect 4628 11632 4637 11666
rect 4637 11632 4671 11666
rect 4671 11632 4680 11666
rect 4628 11623 4680 11632
rect 4862 11537 4914 11550
rect 4862 11503 4868 11537
rect 4868 11503 4902 11537
rect 4902 11503 4914 11537
rect 4862 11498 4914 11503
rect 4552 11367 4604 11419
rect 6868 12106 6920 12158
rect 6250 11780 6302 11832
rect 6974 11778 7026 11830
rect 5117 11621 5169 11673
rect 5934 11654 5986 11664
rect 5934 11620 5942 11654
rect 5942 11620 5976 11654
rect 5976 11620 5986 11654
rect 5934 11612 5986 11620
rect 5015 11500 5067 11552
rect 5714 11360 5766 11368
rect 5778 11360 5830 11368
rect 5714 11326 5734 11360
rect 5734 11326 5766 11360
rect 5778 11326 5806 11360
rect 5806 11326 5830 11360
rect 5714 11316 5766 11326
rect 5778 11316 5830 11326
rect 5842 11360 5894 11368
rect 5842 11326 5844 11360
rect 5844 11326 5878 11360
rect 5878 11326 5894 11360
rect 5842 11316 5894 11326
rect 5906 11360 5958 11368
rect 5906 11326 5916 11360
rect 5916 11326 5950 11360
rect 5950 11326 5958 11360
rect 5906 11316 5958 11326
rect 5970 11360 6022 11368
rect 5970 11326 5988 11360
rect 5988 11326 6022 11360
rect 5970 11316 6022 11326
rect 6034 11360 6086 11368
rect 6098 11360 6150 11368
rect 6034 11326 6060 11360
rect 6060 11326 6086 11360
rect 6098 11326 6132 11360
rect 6132 11326 6150 11360
rect 6034 11316 6086 11326
rect 6098 11316 6150 11326
rect 5117 11167 5169 11219
rect 6586 11666 6638 11676
rect 6586 11632 6596 11666
rect 6596 11632 6630 11666
rect 6630 11632 6638 11666
rect 6586 11624 6638 11632
rect 6820 11538 6872 11550
rect 6820 11504 6826 11538
rect 6826 11504 6860 11538
rect 6860 11504 6872 11538
rect 6820 11498 6872 11504
rect 6510 11368 6562 11420
rect 6974 11500 7026 11552
rect 5035 10997 5087 11049
rect 6974 10970 7026 11022
rect 1398 10822 1450 10831
rect 1462 10822 1514 10831
rect 1398 10788 1417 10822
rect 1417 10788 1450 10822
rect 1462 10788 1489 10822
rect 1489 10788 1514 10822
rect 1398 10779 1450 10788
rect 1462 10779 1514 10788
rect 1526 10822 1578 10831
rect 1526 10788 1527 10822
rect 1527 10788 1561 10822
rect 1561 10788 1578 10822
rect 1526 10779 1578 10788
rect 1590 10822 1642 10831
rect 1590 10788 1599 10822
rect 1599 10788 1633 10822
rect 1633 10788 1642 10822
rect 1590 10779 1642 10788
rect 1654 10822 1706 10831
rect 1654 10788 1671 10822
rect 1671 10788 1705 10822
rect 1705 10788 1706 10822
rect 1654 10779 1706 10788
rect 1718 10822 1770 10831
rect 1782 10822 1834 10831
rect 1718 10788 1743 10822
rect 1743 10788 1770 10822
rect 1782 10788 1815 10822
rect 1815 10788 1834 10822
rect 1718 10779 1770 10788
rect 1782 10779 1834 10788
rect 560 10736 612 10760
rect 560 10708 566 10736
rect 566 10708 607 10736
rect 607 10708 612 10736
rect 702 10736 754 10756
rect 702 10704 710 10736
rect 710 10704 751 10736
rect 751 10704 754 10736
rect 378 10543 433 10598
rect 852 10554 904 10606
rect 378 10258 433 10313
rect 1004 10462 1056 10514
rect 1935 10473 1987 10525
rect 3776 10821 3828 10830
rect 3840 10821 3892 10830
rect 3904 10821 3956 10830
rect 3968 10821 4020 10830
rect 4032 10821 4084 10830
rect 4096 10821 4148 10830
rect 4160 10821 4212 10830
rect 3776 10787 3797 10821
rect 3797 10787 3828 10821
rect 3840 10787 3869 10821
rect 3869 10787 3892 10821
rect 3904 10787 3941 10821
rect 3941 10787 3956 10821
rect 3968 10787 3975 10821
rect 3975 10787 4013 10821
rect 4013 10787 4020 10821
rect 4032 10787 4047 10821
rect 4047 10787 4084 10821
rect 4096 10787 4119 10821
rect 4119 10787 4148 10821
rect 4160 10787 4191 10821
rect 4191 10787 4212 10821
rect 3776 10778 3828 10787
rect 3840 10778 3892 10787
rect 3904 10778 3956 10787
rect 3968 10778 4020 10787
rect 4032 10778 4084 10787
rect 4096 10778 4148 10787
rect 4160 10778 4212 10787
rect 2769 10664 2821 10716
rect 1155 10373 1207 10425
rect 1758 10415 1810 10424
rect 1758 10381 1773 10415
rect 1773 10381 1807 10415
rect 1807 10381 1810 10415
rect 1758 10372 1810 10381
rect 2270 10413 2322 10422
rect 2270 10379 2273 10413
rect 2273 10379 2307 10413
rect 2307 10379 2322 10413
rect 2270 10370 2322 10379
rect 3268 10587 3278 10611
rect 3278 10587 3312 10611
rect 3312 10587 3320 10611
rect 3268 10559 3320 10587
rect 4744 10878 4796 10930
rect 5734 10820 5786 10830
rect 5798 10820 5850 10830
rect 5862 10820 5914 10830
rect 5926 10820 5978 10830
rect 5990 10820 6042 10830
rect 6054 10820 6106 10830
rect 6118 10820 6170 10830
rect 5734 10786 5756 10820
rect 5756 10786 5786 10820
rect 5798 10786 5828 10820
rect 5828 10786 5850 10820
rect 5862 10786 5900 10820
rect 5900 10786 5914 10820
rect 5926 10786 5934 10820
rect 5934 10786 5972 10820
rect 5972 10786 5978 10820
rect 5990 10786 6006 10820
rect 6006 10786 6042 10820
rect 6054 10786 6078 10820
rect 6078 10786 6106 10820
rect 6118 10786 6150 10820
rect 6150 10786 6170 10820
rect 5734 10778 5786 10786
rect 5798 10778 5850 10786
rect 5862 10778 5914 10786
rect 5926 10778 5978 10786
rect 5990 10778 6042 10786
rect 6054 10778 6106 10786
rect 6118 10778 6170 10786
rect 4292 10551 4344 10603
rect 5016 10550 5068 10602
rect 1248 10262 1300 10314
rect 378 10158 434 10214
rect 2020 10297 2072 10314
rect 2020 10263 2030 10297
rect 2030 10263 2064 10297
rect 2064 10263 2072 10297
rect 2020 10262 2072 10263
rect 2522 10297 2574 10312
rect 2522 10263 2530 10297
rect 2530 10263 2564 10297
rect 2564 10263 2574 10297
rect 2522 10260 2574 10263
rect 2842 10411 2894 10420
rect 2842 10377 2857 10411
rect 2857 10377 2891 10411
rect 2891 10377 2894 10411
rect 2842 10368 2894 10377
rect 3268 10366 3320 10418
rect 3561 10393 3613 10445
rect 3976 10426 4028 10436
rect 3976 10392 3984 10426
rect 3984 10392 4018 10426
rect 4018 10392 4028 10426
rect 3976 10384 4028 10392
rect 2766 10297 2818 10324
rect 2766 10272 2776 10297
rect 2776 10272 2810 10297
rect 2810 10272 2818 10297
rect 1360 10120 1412 10129
rect 1360 10086 1373 10120
rect 1373 10086 1407 10120
rect 1407 10086 1412 10120
rect 1360 10077 1412 10086
rect 1424 10120 1476 10129
rect 1488 10120 1540 10129
rect 1552 10120 1604 10129
rect 1616 10120 1668 10129
rect 1680 10120 1732 10129
rect 1744 10120 1796 10129
rect 1808 10120 1860 10129
rect 1424 10086 1445 10120
rect 1445 10086 1476 10120
rect 1488 10086 1517 10120
rect 1517 10086 1540 10120
rect 1552 10086 1589 10120
rect 1589 10086 1604 10120
rect 1616 10086 1623 10120
rect 1623 10086 1661 10120
rect 1661 10086 1668 10120
rect 1680 10086 1695 10120
rect 1695 10086 1732 10120
rect 1744 10086 1767 10120
rect 1767 10086 1796 10120
rect 1808 10086 1839 10120
rect 1839 10086 1860 10120
rect 1424 10077 1476 10086
rect 1488 10077 1540 10086
rect 1552 10077 1604 10086
rect 1616 10077 1668 10086
rect 1680 10077 1732 10086
rect 1744 10077 1796 10086
rect 1808 10077 1860 10086
rect 1872 10120 1924 10129
rect 1872 10086 1877 10120
rect 1877 10086 1911 10120
rect 1911 10086 1924 10120
rect 1872 10077 1924 10086
rect 3756 10131 3808 10140
rect 3820 10131 3872 10140
rect 278 9945 332 9999
rect 3756 10097 3775 10131
rect 3775 10097 3808 10131
rect 3820 10097 3847 10131
rect 3847 10097 3872 10131
rect 3756 10088 3808 10097
rect 3820 10088 3872 10097
rect 3884 10131 3936 10140
rect 3884 10097 3885 10131
rect 3885 10097 3919 10131
rect 3919 10097 3936 10131
rect 3884 10088 3936 10097
rect 3948 10131 4000 10140
rect 3948 10097 3957 10131
rect 3957 10097 3991 10131
rect 3991 10097 4000 10131
rect 3948 10088 4000 10097
rect 4012 10131 4064 10140
rect 4012 10097 4029 10131
rect 4029 10097 4063 10131
rect 4063 10097 4064 10131
rect 4012 10088 4064 10097
rect 4076 10131 4128 10140
rect 4140 10131 4192 10140
rect 4076 10097 4101 10131
rect 4101 10097 4128 10131
rect 4140 10097 4173 10131
rect 4173 10097 4192 10131
rect 4076 10088 4128 10097
rect 4140 10088 4192 10097
rect 3565 9939 3617 9991
rect 4628 10438 4680 10447
rect 4628 10404 4637 10438
rect 4637 10404 4671 10438
rect 4671 10404 4680 10438
rect 4628 10395 4680 10404
rect 4862 10309 4914 10322
rect 4862 10275 4868 10309
rect 4868 10275 4902 10309
rect 4902 10275 4914 10309
rect 4862 10270 4914 10275
rect 4552 10139 4604 10191
rect 6835 10878 6887 10930
rect 6250 10552 6302 10604
rect 6974 10550 7026 10602
rect 5356 10393 5408 10445
rect 5934 10426 5986 10436
rect 5934 10392 5942 10426
rect 5942 10392 5976 10426
rect 5976 10392 5986 10426
rect 5934 10384 5986 10392
rect 5015 10272 5067 10324
rect 5714 10132 5766 10140
rect 5778 10132 5830 10140
rect 5714 10098 5734 10132
rect 5734 10098 5766 10132
rect 5778 10098 5806 10132
rect 5806 10098 5830 10132
rect 5714 10088 5766 10098
rect 5778 10088 5830 10098
rect 5842 10132 5894 10140
rect 5842 10098 5844 10132
rect 5844 10098 5878 10132
rect 5878 10098 5894 10132
rect 5842 10088 5894 10098
rect 5906 10132 5958 10140
rect 5906 10098 5916 10132
rect 5916 10098 5950 10132
rect 5950 10098 5958 10132
rect 5906 10088 5958 10098
rect 5970 10132 6022 10140
rect 5970 10098 5988 10132
rect 5988 10098 6022 10132
rect 5970 10088 6022 10098
rect 6034 10132 6086 10140
rect 6098 10132 6150 10140
rect 6034 10098 6060 10132
rect 6060 10098 6086 10132
rect 6098 10098 6132 10132
rect 6132 10098 6150 10132
rect 6034 10088 6086 10098
rect 6098 10088 6150 10098
rect 5354 9939 5406 9991
rect 6586 10438 6638 10448
rect 6586 10404 6596 10438
rect 6596 10404 6630 10438
rect 6630 10404 6638 10438
rect 6586 10396 6638 10404
rect 6820 10310 6872 10322
rect 6820 10276 6826 10310
rect 6826 10276 6860 10310
rect 6860 10276 6872 10310
rect 6820 10270 6872 10276
rect 6510 10140 6562 10192
rect 6974 10272 7026 10324
rect 7085 9958 7137 10010
rect 1398 9594 1450 9603
rect 1462 9594 1514 9603
rect 1398 9560 1417 9594
rect 1417 9560 1450 9594
rect 1462 9560 1489 9594
rect 1489 9560 1514 9594
rect 1398 9551 1450 9560
rect 1462 9551 1514 9560
rect 1526 9594 1578 9603
rect 1526 9560 1527 9594
rect 1527 9560 1561 9594
rect 1561 9560 1578 9594
rect 1526 9551 1578 9560
rect 1590 9594 1642 9603
rect 1590 9560 1599 9594
rect 1599 9560 1633 9594
rect 1633 9560 1642 9594
rect 1590 9551 1642 9560
rect 1654 9594 1706 9603
rect 1654 9560 1671 9594
rect 1671 9560 1705 9594
rect 1705 9560 1706 9594
rect 1654 9551 1706 9560
rect 1718 9594 1770 9603
rect 1782 9594 1834 9603
rect 1718 9560 1743 9594
rect 1743 9560 1770 9594
rect 1782 9560 1815 9594
rect 1815 9560 1834 9594
rect 1718 9551 1770 9560
rect 1782 9551 1834 9560
rect 560 9508 612 9532
rect 560 9480 566 9508
rect 566 9480 607 9508
rect 607 9480 612 9508
rect 702 9508 754 9528
rect 702 9476 710 9508
rect 710 9476 751 9508
rect 751 9476 754 9508
rect 378 9315 433 9370
rect 852 9326 904 9378
rect 378 9030 433 9085
rect 1004 9234 1056 9286
rect 1935 9245 1987 9297
rect 3776 9593 3828 9602
rect 3840 9593 3892 9602
rect 3904 9593 3956 9602
rect 3968 9593 4020 9602
rect 4032 9593 4084 9602
rect 4096 9593 4148 9602
rect 4160 9593 4212 9602
rect 3776 9559 3797 9593
rect 3797 9559 3828 9593
rect 3840 9559 3869 9593
rect 3869 9559 3892 9593
rect 3904 9559 3941 9593
rect 3941 9559 3956 9593
rect 3968 9559 3975 9593
rect 3975 9559 4013 9593
rect 4013 9559 4020 9593
rect 4032 9559 4047 9593
rect 4047 9559 4084 9593
rect 4096 9559 4119 9593
rect 4119 9559 4148 9593
rect 4160 9559 4191 9593
rect 4191 9559 4212 9593
rect 3776 9550 3828 9559
rect 3840 9550 3892 9559
rect 3904 9550 3956 9559
rect 3968 9550 4020 9559
rect 4032 9550 4084 9559
rect 4096 9550 4148 9559
rect 4160 9550 4212 9559
rect 2769 9436 2821 9488
rect 1155 9145 1207 9197
rect 1758 9187 1810 9196
rect 1758 9153 1773 9187
rect 1773 9153 1807 9187
rect 1807 9153 1810 9187
rect 1758 9144 1810 9153
rect 2270 9185 2322 9194
rect 2270 9151 2273 9185
rect 2273 9151 2307 9185
rect 2307 9151 2322 9185
rect 2270 9142 2322 9151
rect 3268 9359 3278 9383
rect 3278 9359 3312 9383
rect 3312 9359 3320 9383
rect 3268 9331 3320 9359
rect 4744 9650 4796 9702
rect 5029 9732 5081 9784
rect 5734 9592 5786 9602
rect 5798 9592 5850 9602
rect 5862 9592 5914 9602
rect 5926 9592 5978 9602
rect 5990 9592 6042 9602
rect 6054 9592 6106 9602
rect 6118 9592 6170 9602
rect 5734 9558 5756 9592
rect 5756 9558 5786 9592
rect 5798 9558 5828 9592
rect 5828 9558 5850 9592
rect 5862 9558 5900 9592
rect 5900 9558 5914 9592
rect 5926 9558 5934 9592
rect 5934 9558 5972 9592
rect 5972 9558 5978 9592
rect 5990 9558 6006 9592
rect 6006 9558 6042 9592
rect 6054 9558 6078 9592
rect 6078 9558 6106 9592
rect 6118 9558 6150 9592
rect 6150 9558 6170 9592
rect 5734 9550 5786 9558
rect 5798 9550 5850 9558
rect 5862 9550 5914 9558
rect 5926 9550 5978 9558
rect 5990 9550 6042 9558
rect 6054 9550 6106 9558
rect 6118 9550 6170 9558
rect 4292 9323 4344 9375
rect 5016 9322 5068 9374
rect 1248 9034 1300 9086
rect 378 8930 434 8986
rect 2020 9069 2072 9086
rect 2020 9035 2030 9069
rect 2030 9035 2064 9069
rect 2064 9035 2072 9069
rect 2020 9034 2072 9035
rect 2522 9069 2574 9084
rect 2522 9035 2530 9069
rect 2530 9035 2564 9069
rect 2564 9035 2574 9069
rect 2522 9032 2574 9035
rect 2842 9183 2894 9192
rect 2842 9149 2857 9183
rect 2857 9149 2891 9183
rect 2891 9149 2894 9183
rect 2842 9140 2894 9149
rect 3268 9138 3320 9190
rect 3561 9165 3613 9217
rect 3976 9198 4028 9208
rect 3976 9164 3984 9198
rect 3984 9164 4018 9198
rect 4018 9164 4028 9198
rect 3976 9156 4028 9164
rect 2766 9069 2818 9096
rect 2766 9044 2776 9069
rect 2776 9044 2810 9069
rect 2810 9044 2818 9069
rect 1360 8892 1412 8901
rect 1360 8858 1373 8892
rect 1373 8858 1407 8892
rect 1407 8858 1412 8892
rect 1360 8849 1412 8858
rect 1424 8892 1476 8901
rect 1488 8892 1540 8901
rect 1552 8892 1604 8901
rect 1616 8892 1668 8901
rect 1680 8892 1732 8901
rect 1744 8892 1796 8901
rect 1808 8892 1860 8901
rect 1424 8858 1445 8892
rect 1445 8858 1476 8892
rect 1488 8858 1517 8892
rect 1517 8858 1540 8892
rect 1552 8858 1589 8892
rect 1589 8858 1604 8892
rect 1616 8858 1623 8892
rect 1623 8858 1661 8892
rect 1661 8858 1668 8892
rect 1680 8858 1695 8892
rect 1695 8858 1732 8892
rect 1744 8858 1767 8892
rect 1767 8858 1796 8892
rect 1808 8858 1839 8892
rect 1839 8858 1860 8892
rect 1424 8849 1476 8858
rect 1488 8849 1540 8858
rect 1552 8849 1604 8858
rect 1616 8849 1668 8858
rect 1680 8849 1732 8858
rect 1744 8849 1796 8858
rect 1808 8849 1860 8858
rect 1872 8892 1924 8901
rect 1872 8858 1877 8892
rect 1877 8858 1911 8892
rect 1911 8858 1924 8892
rect 1872 8849 1924 8858
rect 3756 8903 3808 8912
rect 3820 8903 3872 8912
rect 278 8717 332 8771
rect 3756 8869 3775 8903
rect 3775 8869 3808 8903
rect 3820 8869 3847 8903
rect 3847 8869 3872 8903
rect 3756 8860 3808 8869
rect 3820 8860 3872 8869
rect 3884 8903 3936 8912
rect 3884 8869 3885 8903
rect 3885 8869 3919 8903
rect 3919 8869 3936 8903
rect 3884 8860 3936 8869
rect 3948 8903 4000 8912
rect 3948 8869 3957 8903
rect 3957 8869 3991 8903
rect 3991 8869 4000 8903
rect 3948 8860 4000 8869
rect 4012 8903 4064 8912
rect 4012 8869 4029 8903
rect 4029 8869 4063 8903
rect 4063 8869 4064 8903
rect 4012 8860 4064 8869
rect 4076 8903 4128 8912
rect 4140 8903 4192 8912
rect 4076 8869 4101 8903
rect 4101 8869 4128 8903
rect 4140 8869 4173 8903
rect 4173 8869 4192 8903
rect 4076 8860 4128 8869
rect 4140 8860 4192 8869
rect 3565 8711 3617 8763
rect 4628 9210 4680 9219
rect 4628 9176 4637 9210
rect 4637 9176 4671 9210
rect 4671 9176 4680 9210
rect 4628 9167 4680 9176
rect 4862 9081 4914 9094
rect 4862 9047 4868 9081
rect 4868 9047 4902 9081
rect 4902 9047 4914 9081
rect 4862 9042 4914 9047
rect 4552 8911 4604 8963
rect 6868 9650 6920 9702
rect 6250 9324 6302 9376
rect 6974 9322 7026 9374
rect 5117 9165 5169 9217
rect 5934 9198 5986 9208
rect 5934 9164 5942 9198
rect 5942 9164 5976 9198
rect 5976 9164 5986 9198
rect 5934 9156 5986 9164
rect 5015 9044 5067 9096
rect 5714 8904 5766 8912
rect 5778 8904 5830 8912
rect 5714 8870 5734 8904
rect 5734 8870 5766 8904
rect 5778 8870 5806 8904
rect 5806 8870 5830 8904
rect 5714 8860 5766 8870
rect 5778 8860 5830 8870
rect 5842 8904 5894 8912
rect 5842 8870 5844 8904
rect 5844 8870 5878 8904
rect 5878 8870 5894 8904
rect 5842 8860 5894 8870
rect 5906 8904 5958 8912
rect 5906 8870 5916 8904
rect 5916 8870 5950 8904
rect 5950 8870 5958 8904
rect 5906 8860 5958 8870
rect 5970 8904 6022 8912
rect 5970 8870 5988 8904
rect 5988 8870 6022 8904
rect 5970 8860 6022 8870
rect 6034 8904 6086 8912
rect 6098 8904 6150 8912
rect 6034 8870 6060 8904
rect 6060 8870 6086 8904
rect 6098 8870 6132 8904
rect 6132 8870 6150 8904
rect 6034 8860 6086 8870
rect 6098 8860 6150 8870
rect 5117 8711 5169 8763
rect 6586 9210 6638 9220
rect 6586 9176 6596 9210
rect 6596 9176 6630 9210
rect 6630 9176 6638 9210
rect 6586 9168 6638 9176
rect 6820 9082 6872 9094
rect 6820 9048 6826 9082
rect 6826 9048 6860 9082
rect 6860 9048 6872 9082
rect 6820 9042 6872 9048
rect 6510 8912 6562 8964
rect 6974 9044 7026 9096
rect 5035 8541 5087 8593
rect 6512 8626 6564 8678
rect 1398 8366 1450 8375
rect 1462 8366 1514 8375
rect 1398 8332 1417 8366
rect 1417 8332 1450 8366
rect 1462 8332 1489 8366
rect 1489 8332 1514 8366
rect 1398 8323 1450 8332
rect 1462 8323 1514 8332
rect 1526 8366 1578 8375
rect 1526 8332 1527 8366
rect 1527 8332 1561 8366
rect 1561 8332 1578 8366
rect 1526 8323 1578 8332
rect 1590 8366 1642 8375
rect 1590 8332 1599 8366
rect 1599 8332 1633 8366
rect 1633 8332 1642 8366
rect 1590 8323 1642 8332
rect 1654 8366 1706 8375
rect 1654 8332 1671 8366
rect 1671 8332 1705 8366
rect 1705 8332 1706 8366
rect 1654 8323 1706 8332
rect 1718 8366 1770 8375
rect 1782 8366 1834 8375
rect 1718 8332 1743 8366
rect 1743 8332 1770 8366
rect 1782 8332 1815 8366
rect 1815 8332 1834 8366
rect 1718 8323 1770 8332
rect 1782 8323 1834 8332
rect 560 8280 612 8304
rect 560 8252 566 8280
rect 566 8252 607 8280
rect 607 8252 612 8280
rect 702 8280 754 8300
rect 702 8248 710 8280
rect 710 8248 751 8280
rect 751 8248 754 8280
rect 378 8087 433 8142
rect 852 8098 904 8150
rect 378 7802 433 7857
rect 1004 8006 1056 8058
rect 1935 8017 1987 8069
rect 3776 8365 3828 8374
rect 3840 8365 3892 8374
rect 3904 8365 3956 8374
rect 3968 8365 4020 8374
rect 4032 8365 4084 8374
rect 4096 8365 4148 8374
rect 4160 8365 4212 8374
rect 3776 8331 3797 8365
rect 3797 8331 3828 8365
rect 3840 8331 3869 8365
rect 3869 8331 3892 8365
rect 3904 8331 3941 8365
rect 3941 8331 3956 8365
rect 3968 8331 3975 8365
rect 3975 8331 4013 8365
rect 4013 8331 4020 8365
rect 4032 8331 4047 8365
rect 4047 8331 4084 8365
rect 4096 8331 4119 8365
rect 4119 8331 4148 8365
rect 4160 8331 4191 8365
rect 4191 8331 4212 8365
rect 3776 8322 3828 8331
rect 3840 8322 3892 8331
rect 3904 8322 3956 8331
rect 3968 8322 4020 8331
rect 4032 8322 4084 8331
rect 4096 8322 4148 8331
rect 4160 8322 4212 8331
rect 2769 8208 2821 8260
rect 1155 7917 1207 7969
rect 1758 7959 1810 7968
rect 1758 7925 1773 7959
rect 1773 7925 1807 7959
rect 1807 7925 1810 7959
rect 1758 7916 1810 7925
rect 2270 7957 2322 7966
rect 2270 7923 2273 7957
rect 2273 7923 2307 7957
rect 2307 7923 2322 7957
rect 2270 7914 2322 7923
rect 3268 8131 3278 8155
rect 3278 8131 3312 8155
rect 3312 8131 3320 8155
rect 3268 8103 3320 8131
rect 4744 8422 4796 8474
rect 5734 8364 5786 8374
rect 5798 8364 5850 8374
rect 5862 8364 5914 8374
rect 5926 8364 5978 8374
rect 5990 8364 6042 8374
rect 6054 8364 6106 8374
rect 6118 8364 6170 8374
rect 5734 8330 5756 8364
rect 5756 8330 5786 8364
rect 5798 8330 5828 8364
rect 5828 8330 5850 8364
rect 5862 8330 5900 8364
rect 5900 8330 5914 8364
rect 5926 8330 5934 8364
rect 5934 8330 5972 8364
rect 5972 8330 5978 8364
rect 5990 8330 6006 8364
rect 6006 8330 6042 8364
rect 6054 8330 6078 8364
rect 6078 8330 6106 8364
rect 6118 8330 6150 8364
rect 6150 8330 6170 8364
rect 5734 8322 5786 8330
rect 5798 8322 5850 8330
rect 5862 8322 5914 8330
rect 5926 8322 5978 8330
rect 5990 8322 6042 8330
rect 6054 8322 6106 8330
rect 6118 8322 6170 8330
rect 4292 8095 4344 8147
rect 5016 8094 5068 8146
rect 1248 7806 1300 7858
rect 378 7702 434 7758
rect 2020 7841 2072 7858
rect 2020 7807 2030 7841
rect 2030 7807 2064 7841
rect 2064 7807 2072 7841
rect 2020 7806 2072 7807
rect 2522 7841 2574 7856
rect 2522 7807 2530 7841
rect 2530 7807 2564 7841
rect 2564 7807 2574 7841
rect 2522 7804 2574 7807
rect 2842 7955 2894 7964
rect 2842 7921 2857 7955
rect 2857 7921 2891 7955
rect 2891 7921 2894 7955
rect 2842 7912 2894 7921
rect 3268 7910 3320 7962
rect 3561 7937 3613 7989
rect 3976 7970 4028 7980
rect 3976 7936 3984 7970
rect 3984 7936 4018 7970
rect 4018 7936 4028 7970
rect 3976 7928 4028 7936
rect 2766 7841 2818 7868
rect 2766 7816 2776 7841
rect 2776 7816 2810 7841
rect 2810 7816 2818 7841
rect 1360 7664 1412 7673
rect 1360 7630 1373 7664
rect 1373 7630 1407 7664
rect 1407 7630 1412 7664
rect 1360 7621 1412 7630
rect 1424 7664 1476 7673
rect 1488 7664 1540 7673
rect 1552 7664 1604 7673
rect 1616 7664 1668 7673
rect 1680 7664 1732 7673
rect 1744 7664 1796 7673
rect 1808 7664 1860 7673
rect 1424 7630 1445 7664
rect 1445 7630 1476 7664
rect 1488 7630 1517 7664
rect 1517 7630 1540 7664
rect 1552 7630 1589 7664
rect 1589 7630 1604 7664
rect 1616 7630 1623 7664
rect 1623 7630 1661 7664
rect 1661 7630 1668 7664
rect 1680 7630 1695 7664
rect 1695 7630 1732 7664
rect 1744 7630 1767 7664
rect 1767 7630 1796 7664
rect 1808 7630 1839 7664
rect 1839 7630 1860 7664
rect 1424 7621 1476 7630
rect 1488 7621 1540 7630
rect 1552 7621 1604 7630
rect 1616 7621 1668 7630
rect 1680 7621 1732 7630
rect 1744 7621 1796 7630
rect 1808 7621 1860 7630
rect 1872 7664 1924 7673
rect 1872 7630 1877 7664
rect 1877 7630 1911 7664
rect 1911 7630 1924 7664
rect 1872 7621 1924 7630
rect 3756 7675 3808 7684
rect 3820 7675 3872 7684
rect 278 7489 332 7543
rect 3756 7641 3775 7675
rect 3775 7641 3808 7675
rect 3820 7641 3847 7675
rect 3847 7641 3872 7675
rect 3756 7632 3808 7641
rect 3820 7632 3872 7641
rect 3884 7675 3936 7684
rect 3884 7641 3885 7675
rect 3885 7641 3919 7675
rect 3919 7641 3936 7675
rect 3884 7632 3936 7641
rect 3948 7675 4000 7684
rect 3948 7641 3957 7675
rect 3957 7641 3991 7675
rect 3991 7641 4000 7675
rect 3948 7632 4000 7641
rect 4012 7675 4064 7684
rect 4012 7641 4029 7675
rect 4029 7641 4063 7675
rect 4063 7641 4064 7675
rect 4012 7632 4064 7641
rect 4076 7675 4128 7684
rect 4140 7675 4192 7684
rect 4076 7641 4101 7675
rect 4101 7641 4128 7675
rect 4140 7641 4173 7675
rect 4173 7641 4192 7675
rect 4076 7632 4128 7641
rect 4140 7632 4192 7641
rect 3565 7483 3617 7535
rect 4628 7982 4680 7991
rect 4628 7948 4637 7982
rect 4637 7948 4671 7982
rect 4671 7948 4680 7982
rect 4628 7939 4680 7948
rect 4862 7853 4914 7866
rect 4862 7819 4868 7853
rect 4868 7819 4902 7853
rect 4902 7819 4914 7853
rect 4862 7814 4914 7819
rect 4552 7683 4604 7735
rect 6843 8422 6895 8474
rect 6250 8096 6302 8148
rect 6974 8094 7026 8146
rect 5197 7937 5249 7989
rect 5934 7970 5986 7980
rect 5934 7936 5942 7970
rect 5942 7936 5976 7970
rect 5976 7936 5986 7970
rect 5934 7928 5986 7936
rect 5015 7816 5067 7868
rect 5714 7676 5766 7684
rect 5778 7676 5830 7684
rect 5714 7642 5734 7676
rect 5734 7642 5766 7676
rect 5778 7642 5806 7676
rect 5806 7642 5830 7676
rect 5714 7632 5766 7642
rect 5778 7632 5830 7642
rect 5842 7676 5894 7684
rect 5842 7642 5844 7676
rect 5844 7642 5878 7676
rect 5878 7642 5894 7676
rect 5842 7632 5894 7642
rect 5906 7676 5958 7684
rect 5906 7642 5916 7676
rect 5916 7642 5950 7676
rect 5950 7642 5958 7676
rect 5906 7632 5958 7642
rect 5970 7676 6022 7684
rect 5970 7642 5988 7676
rect 5988 7642 6022 7676
rect 5970 7632 6022 7642
rect 6034 7676 6086 7684
rect 6098 7676 6150 7684
rect 6034 7642 6060 7676
rect 6060 7642 6086 7676
rect 6098 7642 6132 7676
rect 6132 7642 6150 7676
rect 6034 7632 6086 7642
rect 6098 7632 6150 7642
rect 5197 7483 5249 7535
rect 6586 7982 6638 7992
rect 6586 7948 6596 7982
rect 6596 7948 6630 7982
rect 6630 7948 6638 7982
rect 6586 7940 6638 7948
rect 6820 7854 6872 7866
rect 6820 7820 6826 7854
rect 6826 7820 6860 7854
rect 6860 7820 6872 7854
rect 6820 7814 6872 7820
rect 6510 7684 6562 7736
rect 6974 7816 7026 7868
rect 7107 7396 7159 7448
rect 1398 7138 1450 7147
rect 1462 7138 1514 7147
rect 1398 7104 1417 7138
rect 1417 7104 1450 7138
rect 1462 7104 1489 7138
rect 1489 7104 1514 7138
rect 1398 7095 1450 7104
rect 1462 7095 1514 7104
rect 1526 7138 1578 7147
rect 1526 7104 1527 7138
rect 1527 7104 1561 7138
rect 1561 7104 1578 7138
rect 1526 7095 1578 7104
rect 1590 7138 1642 7147
rect 1590 7104 1599 7138
rect 1599 7104 1633 7138
rect 1633 7104 1642 7138
rect 1590 7095 1642 7104
rect 1654 7138 1706 7147
rect 1654 7104 1671 7138
rect 1671 7104 1705 7138
rect 1705 7104 1706 7138
rect 1654 7095 1706 7104
rect 1718 7138 1770 7147
rect 1782 7138 1834 7147
rect 1718 7104 1743 7138
rect 1743 7104 1770 7138
rect 1782 7104 1815 7138
rect 1815 7104 1834 7138
rect 1718 7095 1770 7104
rect 1782 7095 1834 7104
rect 560 7052 612 7076
rect 560 7024 566 7052
rect 566 7024 607 7052
rect 607 7024 612 7052
rect 702 7052 754 7072
rect 702 7020 710 7052
rect 710 7020 751 7052
rect 751 7020 754 7052
rect 378 6859 433 6914
rect 852 6870 904 6922
rect 378 6574 433 6629
rect 1004 6778 1056 6830
rect 1935 6789 1987 6841
rect 3776 7137 3828 7146
rect 3840 7137 3892 7146
rect 3904 7137 3956 7146
rect 3968 7137 4020 7146
rect 4032 7137 4084 7146
rect 4096 7137 4148 7146
rect 4160 7137 4212 7146
rect 3776 7103 3797 7137
rect 3797 7103 3828 7137
rect 3840 7103 3869 7137
rect 3869 7103 3892 7137
rect 3904 7103 3941 7137
rect 3941 7103 3956 7137
rect 3968 7103 3975 7137
rect 3975 7103 4013 7137
rect 4013 7103 4020 7137
rect 4032 7103 4047 7137
rect 4047 7103 4084 7137
rect 4096 7103 4119 7137
rect 4119 7103 4148 7137
rect 4160 7103 4191 7137
rect 4191 7103 4212 7137
rect 3776 7094 3828 7103
rect 3840 7094 3892 7103
rect 3904 7094 3956 7103
rect 3968 7094 4020 7103
rect 4032 7094 4084 7103
rect 4096 7094 4148 7103
rect 4160 7094 4212 7103
rect 2769 6980 2821 7032
rect 1155 6689 1207 6741
rect 1758 6731 1810 6740
rect 1758 6697 1773 6731
rect 1773 6697 1807 6731
rect 1807 6697 1810 6731
rect 1758 6688 1810 6697
rect 2270 6729 2322 6738
rect 2270 6695 2273 6729
rect 2273 6695 2307 6729
rect 2307 6695 2322 6729
rect 2270 6686 2322 6695
rect 3268 6903 3278 6927
rect 3278 6903 3312 6927
rect 3312 6903 3320 6927
rect 3268 6875 3320 6903
rect 4744 7194 4796 7246
rect 5029 7276 5081 7328
rect 5734 7136 5786 7146
rect 5798 7136 5850 7146
rect 5862 7136 5914 7146
rect 5926 7136 5978 7146
rect 5990 7136 6042 7146
rect 6054 7136 6106 7146
rect 6118 7136 6170 7146
rect 5734 7102 5756 7136
rect 5756 7102 5786 7136
rect 5798 7102 5828 7136
rect 5828 7102 5850 7136
rect 5862 7102 5900 7136
rect 5900 7102 5914 7136
rect 5926 7102 5934 7136
rect 5934 7102 5972 7136
rect 5972 7102 5978 7136
rect 5990 7102 6006 7136
rect 6006 7102 6042 7136
rect 6054 7102 6078 7136
rect 6078 7102 6106 7136
rect 6118 7102 6150 7136
rect 6150 7102 6170 7136
rect 5734 7094 5786 7102
rect 5798 7094 5850 7102
rect 5862 7094 5914 7102
rect 5926 7094 5978 7102
rect 5990 7094 6042 7102
rect 6054 7094 6106 7102
rect 6118 7094 6170 7102
rect 4292 6867 4344 6919
rect 5016 6866 5068 6918
rect 1248 6578 1300 6630
rect 378 6474 434 6530
rect 2020 6613 2072 6630
rect 2020 6579 2030 6613
rect 2030 6579 2064 6613
rect 2064 6579 2072 6613
rect 2020 6578 2072 6579
rect 2522 6613 2574 6628
rect 2522 6579 2530 6613
rect 2530 6579 2564 6613
rect 2564 6579 2574 6613
rect 2522 6576 2574 6579
rect 2842 6727 2894 6736
rect 2842 6693 2857 6727
rect 2857 6693 2891 6727
rect 2891 6693 2894 6727
rect 2842 6684 2894 6693
rect 3268 6682 3320 6734
rect 3561 6709 3613 6761
rect 3976 6742 4028 6752
rect 3976 6708 3984 6742
rect 3984 6708 4018 6742
rect 4018 6708 4028 6742
rect 3976 6700 4028 6708
rect 2766 6613 2818 6640
rect 2766 6588 2776 6613
rect 2776 6588 2810 6613
rect 2810 6588 2818 6613
rect 1360 6436 1412 6445
rect 1360 6402 1373 6436
rect 1373 6402 1407 6436
rect 1407 6402 1412 6436
rect 1360 6393 1412 6402
rect 1424 6436 1476 6445
rect 1488 6436 1540 6445
rect 1552 6436 1604 6445
rect 1616 6436 1668 6445
rect 1680 6436 1732 6445
rect 1744 6436 1796 6445
rect 1808 6436 1860 6445
rect 1424 6402 1445 6436
rect 1445 6402 1476 6436
rect 1488 6402 1517 6436
rect 1517 6402 1540 6436
rect 1552 6402 1589 6436
rect 1589 6402 1604 6436
rect 1616 6402 1623 6436
rect 1623 6402 1661 6436
rect 1661 6402 1668 6436
rect 1680 6402 1695 6436
rect 1695 6402 1732 6436
rect 1744 6402 1767 6436
rect 1767 6402 1796 6436
rect 1808 6402 1839 6436
rect 1839 6402 1860 6436
rect 1424 6393 1476 6402
rect 1488 6393 1540 6402
rect 1552 6393 1604 6402
rect 1616 6393 1668 6402
rect 1680 6393 1732 6402
rect 1744 6393 1796 6402
rect 1808 6393 1860 6402
rect 1872 6436 1924 6445
rect 1872 6402 1877 6436
rect 1877 6402 1911 6436
rect 1911 6402 1924 6436
rect 1872 6393 1924 6402
rect 3756 6447 3808 6456
rect 3820 6447 3872 6456
rect 278 6261 332 6315
rect 3756 6413 3775 6447
rect 3775 6413 3808 6447
rect 3820 6413 3847 6447
rect 3847 6413 3872 6447
rect 3756 6404 3808 6413
rect 3820 6404 3872 6413
rect 3884 6447 3936 6456
rect 3884 6413 3885 6447
rect 3885 6413 3919 6447
rect 3919 6413 3936 6447
rect 3884 6404 3936 6413
rect 3948 6447 4000 6456
rect 3948 6413 3957 6447
rect 3957 6413 3991 6447
rect 3991 6413 4000 6447
rect 3948 6404 4000 6413
rect 4012 6447 4064 6456
rect 4012 6413 4029 6447
rect 4029 6413 4063 6447
rect 4063 6413 4064 6447
rect 4012 6404 4064 6413
rect 4076 6447 4128 6456
rect 4140 6447 4192 6456
rect 4076 6413 4101 6447
rect 4101 6413 4128 6447
rect 4140 6413 4173 6447
rect 4173 6413 4192 6447
rect 4076 6404 4128 6413
rect 4140 6404 4192 6413
rect 3565 6255 3617 6307
rect 4628 6754 4680 6763
rect 4628 6720 4637 6754
rect 4637 6720 4671 6754
rect 4671 6720 4680 6754
rect 4628 6711 4680 6720
rect 4862 6625 4914 6638
rect 4862 6591 4868 6625
rect 4868 6591 4902 6625
rect 4902 6591 4914 6625
rect 4862 6586 4914 6591
rect 4552 6455 4604 6507
rect 6868 7194 6920 7246
rect 6250 6868 6302 6920
rect 6974 6866 7026 6918
rect 5117 6709 5169 6761
rect 5934 6742 5986 6752
rect 5934 6708 5942 6742
rect 5942 6708 5976 6742
rect 5976 6708 5986 6742
rect 5934 6700 5986 6708
rect 5015 6588 5067 6640
rect 5714 6448 5766 6456
rect 5778 6448 5830 6456
rect 5714 6414 5734 6448
rect 5734 6414 5766 6448
rect 5778 6414 5806 6448
rect 5806 6414 5830 6448
rect 5714 6404 5766 6414
rect 5778 6404 5830 6414
rect 5842 6448 5894 6456
rect 5842 6414 5844 6448
rect 5844 6414 5878 6448
rect 5878 6414 5894 6448
rect 5842 6404 5894 6414
rect 5906 6448 5958 6456
rect 5906 6414 5916 6448
rect 5916 6414 5950 6448
rect 5950 6414 5958 6448
rect 5906 6404 5958 6414
rect 5970 6448 6022 6456
rect 5970 6414 5988 6448
rect 5988 6414 6022 6448
rect 5970 6404 6022 6414
rect 6034 6448 6086 6456
rect 6098 6448 6150 6456
rect 6034 6414 6060 6448
rect 6060 6414 6086 6448
rect 6098 6414 6132 6448
rect 6132 6414 6150 6448
rect 6034 6404 6086 6414
rect 6098 6404 6150 6414
rect 5117 6255 5169 6307
rect 6586 6754 6638 6764
rect 6586 6720 6596 6754
rect 6596 6720 6630 6754
rect 6630 6720 6638 6754
rect 6586 6712 6638 6720
rect 6820 6626 6872 6638
rect 6820 6592 6826 6626
rect 6826 6592 6860 6626
rect 6860 6592 6872 6626
rect 6820 6586 6872 6592
rect 6510 6456 6562 6508
rect 6974 6588 7026 6640
rect 5035 6085 5087 6137
rect 6974 6086 7026 6138
rect 1398 5910 1450 5919
rect 1462 5910 1514 5919
rect 1398 5876 1417 5910
rect 1417 5876 1450 5910
rect 1462 5876 1489 5910
rect 1489 5876 1514 5910
rect 1398 5867 1450 5876
rect 1462 5867 1514 5876
rect 1526 5910 1578 5919
rect 1526 5876 1527 5910
rect 1527 5876 1561 5910
rect 1561 5876 1578 5910
rect 1526 5867 1578 5876
rect 1590 5910 1642 5919
rect 1590 5876 1599 5910
rect 1599 5876 1633 5910
rect 1633 5876 1642 5910
rect 1590 5867 1642 5876
rect 1654 5910 1706 5919
rect 1654 5876 1671 5910
rect 1671 5876 1705 5910
rect 1705 5876 1706 5910
rect 1654 5867 1706 5876
rect 1718 5910 1770 5919
rect 1782 5910 1834 5919
rect 1718 5876 1743 5910
rect 1743 5876 1770 5910
rect 1782 5876 1815 5910
rect 1815 5876 1834 5910
rect 1718 5867 1770 5876
rect 1782 5867 1834 5876
rect 560 5824 612 5848
rect 560 5796 566 5824
rect 566 5796 607 5824
rect 607 5796 612 5824
rect 702 5824 754 5844
rect 702 5792 710 5824
rect 710 5792 751 5824
rect 751 5792 754 5824
rect 378 5631 433 5686
rect 852 5642 904 5694
rect 378 5346 433 5401
rect 1004 5550 1056 5602
rect 1935 5561 1987 5613
rect 3776 5909 3828 5918
rect 3840 5909 3892 5918
rect 3904 5909 3956 5918
rect 3968 5909 4020 5918
rect 4032 5909 4084 5918
rect 4096 5909 4148 5918
rect 4160 5909 4212 5918
rect 3776 5875 3797 5909
rect 3797 5875 3828 5909
rect 3840 5875 3869 5909
rect 3869 5875 3892 5909
rect 3904 5875 3941 5909
rect 3941 5875 3956 5909
rect 3968 5875 3975 5909
rect 3975 5875 4013 5909
rect 4013 5875 4020 5909
rect 4032 5875 4047 5909
rect 4047 5875 4084 5909
rect 4096 5875 4119 5909
rect 4119 5875 4148 5909
rect 4160 5875 4191 5909
rect 4191 5875 4212 5909
rect 3776 5866 3828 5875
rect 3840 5866 3892 5875
rect 3904 5866 3956 5875
rect 3968 5866 4020 5875
rect 4032 5866 4084 5875
rect 4096 5866 4148 5875
rect 4160 5866 4212 5875
rect 2769 5752 2821 5804
rect 1155 5461 1207 5513
rect 1758 5503 1810 5512
rect 1758 5469 1773 5503
rect 1773 5469 1807 5503
rect 1807 5469 1810 5503
rect 1758 5460 1810 5469
rect 2270 5501 2322 5510
rect 2270 5467 2273 5501
rect 2273 5467 2307 5501
rect 2307 5467 2322 5501
rect 2270 5458 2322 5467
rect 3268 5675 3278 5699
rect 3278 5675 3312 5699
rect 3312 5675 3320 5699
rect 3268 5647 3320 5675
rect 4744 5966 4796 6018
rect 5734 5908 5786 5918
rect 5798 5908 5850 5918
rect 5862 5908 5914 5918
rect 5926 5908 5978 5918
rect 5990 5908 6042 5918
rect 6054 5908 6106 5918
rect 6118 5908 6170 5918
rect 5734 5874 5756 5908
rect 5756 5874 5786 5908
rect 5798 5874 5828 5908
rect 5828 5874 5850 5908
rect 5862 5874 5900 5908
rect 5900 5874 5914 5908
rect 5926 5874 5934 5908
rect 5934 5874 5972 5908
rect 5972 5874 5978 5908
rect 5990 5874 6006 5908
rect 6006 5874 6042 5908
rect 6054 5874 6078 5908
rect 6078 5874 6106 5908
rect 6118 5874 6150 5908
rect 6150 5874 6170 5908
rect 5734 5866 5786 5874
rect 5798 5866 5850 5874
rect 5862 5866 5914 5874
rect 5926 5866 5978 5874
rect 5990 5866 6042 5874
rect 6054 5866 6106 5874
rect 6118 5866 6170 5874
rect 4292 5639 4344 5691
rect 5016 5638 5068 5690
rect 1248 5350 1300 5402
rect 378 5246 434 5302
rect 2020 5385 2072 5402
rect 2020 5351 2030 5385
rect 2030 5351 2064 5385
rect 2064 5351 2072 5385
rect 2020 5350 2072 5351
rect 2522 5385 2574 5400
rect 2522 5351 2530 5385
rect 2530 5351 2564 5385
rect 2564 5351 2574 5385
rect 2522 5348 2574 5351
rect 2842 5499 2894 5508
rect 2842 5465 2857 5499
rect 2857 5465 2891 5499
rect 2891 5465 2894 5499
rect 2842 5456 2894 5465
rect 3268 5454 3320 5506
rect 3561 5481 3613 5533
rect 3976 5514 4028 5524
rect 3976 5480 3984 5514
rect 3984 5480 4018 5514
rect 4018 5480 4028 5514
rect 3976 5472 4028 5480
rect 2766 5385 2818 5412
rect 2766 5360 2776 5385
rect 2776 5360 2810 5385
rect 2810 5360 2818 5385
rect 1360 5208 1412 5217
rect 1360 5174 1373 5208
rect 1373 5174 1407 5208
rect 1407 5174 1412 5208
rect 1360 5165 1412 5174
rect 1424 5208 1476 5217
rect 1488 5208 1540 5217
rect 1552 5208 1604 5217
rect 1616 5208 1668 5217
rect 1680 5208 1732 5217
rect 1744 5208 1796 5217
rect 1808 5208 1860 5217
rect 1424 5174 1445 5208
rect 1445 5174 1476 5208
rect 1488 5174 1517 5208
rect 1517 5174 1540 5208
rect 1552 5174 1589 5208
rect 1589 5174 1604 5208
rect 1616 5174 1623 5208
rect 1623 5174 1661 5208
rect 1661 5174 1668 5208
rect 1680 5174 1695 5208
rect 1695 5174 1732 5208
rect 1744 5174 1767 5208
rect 1767 5174 1796 5208
rect 1808 5174 1839 5208
rect 1839 5174 1860 5208
rect 1424 5165 1476 5174
rect 1488 5165 1540 5174
rect 1552 5165 1604 5174
rect 1616 5165 1668 5174
rect 1680 5165 1732 5174
rect 1744 5165 1796 5174
rect 1808 5165 1860 5174
rect 1872 5208 1924 5217
rect 1872 5174 1877 5208
rect 1877 5174 1911 5208
rect 1911 5174 1924 5208
rect 1872 5165 1924 5174
rect 3756 5219 3808 5228
rect 3820 5219 3872 5228
rect 278 5033 332 5087
rect 3756 5185 3775 5219
rect 3775 5185 3808 5219
rect 3820 5185 3847 5219
rect 3847 5185 3872 5219
rect 3756 5176 3808 5185
rect 3820 5176 3872 5185
rect 3884 5219 3936 5228
rect 3884 5185 3885 5219
rect 3885 5185 3919 5219
rect 3919 5185 3936 5219
rect 3884 5176 3936 5185
rect 3948 5219 4000 5228
rect 3948 5185 3957 5219
rect 3957 5185 3991 5219
rect 3991 5185 4000 5219
rect 3948 5176 4000 5185
rect 4012 5219 4064 5228
rect 4012 5185 4029 5219
rect 4029 5185 4063 5219
rect 4063 5185 4064 5219
rect 4012 5176 4064 5185
rect 4076 5219 4128 5228
rect 4140 5219 4192 5228
rect 4076 5185 4101 5219
rect 4101 5185 4128 5219
rect 4140 5185 4173 5219
rect 4173 5185 4192 5219
rect 4076 5176 4128 5185
rect 4140 5176 4192 5185
rect 3565 5027 3617 5079
rect 4628 5526 4680 5535
rect 4628 5492 4637 5526
rect 4637 5492 4671 5526
rect 4671 5492 4680 5526
rect 4628 5483 4680 5492
rect 4862 5397 4914 5410
rect 4862 5363 4868 5397
rect 4868 5363 4902 5397
rect 4902 5363 4914 5397
rect 4862 5358 4914 5363
rect 4552 5227 4604 5279
rect 6250 5640 6302 5692
rect 6974 5638 7026 5690
rect 5279 5481 5331 5533
rect 5934 5514 5986 5524
rect 5934 5480 5942 5514
rect 5942 5480 5976 5514
rect 5976 5480 5986 5514
rect 5934 5472 5986 5480
rect 5015 5360 5067 5412
rect 5714 5220 5766 5228
rect 5778 5220 5830 5228
rect 5714 5186 5734 5220
rect 5734 5186 5766 5220
rect 5778 5186 5806 5220
rect 5806 5186 5830 5220
rect 5714 5176 5766 5186
rect 5778 5176 5830 5186
rect 5842 5220 5894 5228
rect 5842 5186 5844 5220
rect 5844 5186 5878 5220
rect 5878 5186 5894 5220
rect 5842 5176 5894 5186
rect 5906 5220 5958 5228
rect 5906 5186 5916 5220
rect 5916 5186 5950 5220
rect 5950 5186 5958 5220
rect 5906 5176 5958 5186
rect 5970 5220 6022 5228
rect 5970 5186 5988 5220
rect 5988 5186 6022 5220
rect 5970 5176 6022 5186
rect 6034 5220 6086 5228
rect 6098 5220 6150 5228
rect 6034 5186 6060 5220
rect 6060 5186 6086 5220
rect 6098 5186 6132 5220
rect 6132 5186 6150 5220
rect 6034 5176 6086 5186
rect 6098 5176 6150 5186
rect 5279 5027 5331 5079
rect 6586 5526 6638 5536
rect 6586 5492 6596 5526
rect 6596 5492 6630 5526
rect 6630 5492 6638 5526
rect 6586 5484 6638 5492
rect 6820 5398 6872 5410
rect 6820 5364 6826 5398
rect 6826 5364 6860 5398
rect 6860 5364 6872 5398
rect 6820 5358 6872 5364
rect 6510 5228 6562 5280
rect 6974 5360 7026 5412
rect 1398 4682 1450 4691
rect 1462 4682 1514 4691
rect 1398 4648 1417 4682
rect 1417 4648 1450 4682
rect 1462 4648 1489 4682
rect 1489 4648 1514 4682
rect 1398 4639 1450 4648
rect 1462 4639 1514 4648
rect 1526 4682 1578 4691
rect 1526 4648 1527 4682
rect 1527 4648 1561 4682
rect 1561 4648 1578 4682
rect 1526 4639 1578 4648
rect 1590 4682 1642 4691
rect 1590 4648 1599 4682
rect 1599 4648 1633 4682
rect 1633 4648 1642 4682
rect 1590 4639 1642 4648
rect 1654 4682 1706 4691
rect 1654 4648 1671 4682
rect 1671 4648 1705 4682
rect 1705 4648 1706 4682
rect 1654 4639 1706 4648
rect 1718 4682 1770 4691
rect 1782 4682 1834 4691
rect 1718 4648 1743 4682
rect 1743 4648 1770 4682
rect 1782 4648 1815 4682
rect 1815 4648 1834 4682
rect 1718 4639 1770 4648
rect 1782 4639 1834 4648
rect 560 4596 612 4620
rect 560 4568 566 4596
rect 566 4568 607 4596
rect 607 4568 612 4596
rect 702 4596 754 4616
rect 702 4564 710 4596
rect 710 4564 751 4596
rect 751 4564 754 4596
rect 378 4403 433 4458
rect 852 4414 904 4466
rect 378 4118 433 4173
rect 1004 4322 1056 4374
rect 1935 4333 1987 4385
rect 3776 4681 3828 4690
rect 3840 4681 3892 4690
rect 3904 4681 3956 4690
rect 3968 4681 4020 4690
rect 4032 4681 4084 4690
rect 4096 4681 4148 4690
rect 4160 4681 4212 4690
rect 3776 4647 3797 4681
rect 3797 4647 3828 4681
rect 3840 4647 3869 4681
rect 3869 4647 3892 4681
rect 3904 4647 3941 4681
rect 3941 4647 3956 4681
rect 3968 4647 3975 4681
rect 3975 4647 4013 4681
rect 4013 4647 4020 4681
rect 4032 4647 4047 4681
rect 4047 4647 4084 4681
rect 4096 4647 4119 4681
rect 4119 4647 4148 4681
rect 4160 4647 4191 4681
rect 4191 4647 4212 4681
rect 3776 4638 3828 4647
rect 3840 4638 3892 4647
rect 3904 4638 3956 4647
rect 3968 4638 4020 4647
rect 4032 4638 4084 4647
rect 4096 4638 4148 4647
rect 4160 4638 4212 4647
rect 2769 4524 2821 4576
rect 1155 4233 1207 4285
rect 1758 4275 1810 4284
rect 1758 4241 1773 4275
rect 1773 4241 1807 4275
rect 1807 4241 1810 4275
rect 1758 4232 1810 4241
rect 2270 4273 2322 4282
rect 2270 4239 2273 4273
rect 2273 4239 2307 4273
rect 2307 4239 2322 4273
rect 2270 4230 2322 4239
rect 3268 4447 3278 4471
rect 3278 4447 3312 4471
rect 3312 4447 3320 4471
rect 3268 4419 3320 4447
rect 4744 4738 4796 4790
rect 5029 4820 5081 4872
rect 5734 4680 5786 4690
rect 5798 4680 5850 4690
rect 5862 4680 5914 4690
rect 5926 4680 5978 4690
rect 5990 4680 6042 4690
rect 6054 4680 6106 4690
rect 6118 4680 6170 4690
rect 5734 4646 5756 4680
rect 5756 4646 5786 4680
rect 5798 4646 5828 4680
rect 5828 4646 5850 4680
rect 5862 4646 5900 4680
rect 5900 4646 5914 4680
rect 5926 4646 5934 4680
rect 5934 4646 5972 4680
rect 5972 4646 5978 4680
rect 5990 4646 6006 4680
rect 6006 4646 6042 4680
rect 6054 4646 6078 4680
rect 6078 4646 6106 4680
rect 6118 4646 6150 4680
rect 6150 4646 6170 4680
rect 5734 4638 5786 4646
rect 5798 4638 5850 4646
rect 5862 4638 5914 4646
rect 5926 4638 5978 4646
rect 5990 4638 6042 4646
rect 6054 4638 6106 4646
rect 6118 4638 6170 4646
rect 4292 4411 4344 4463
rect 5016 4410 5068 4462
rect 1248 4122 1300 4174
rect 378 4018 434 4074
rect 2020 4157 2072 4174
rect 2020 4123 2030 4157
rect 2030 4123 2064 4157
rect 2064 4123 2072 4157
rect 2020 4122 2072 4123
rect 2522 4157 2574 4172
rect 2522 4123 2530 4157
rect 2530 4123 2564 4157
rect 2564 4123 2574 4157
rect 2522 4120 2574 4123
rect 2842 4271 2894 4280
rect 2842 4237 2857 4271
rect 2857 4237 2891 4271
rect 2891 4237 2894 4271
rect 2842 4228 2894 4237
rect 3268 4226 3320 4278
rect 3561 4253 3613 4305
rect 3976 4286 4028 4296
rect 3976 4252 3984 4286
rect 3984 4252 4018 4286
rect 4018 4252 4028 4286
rect 3976 4244 4028 4252
rect 2766 4157 2818 4184
rect 2766 4132 2776 4157
rect 2776 4132 2810 4157
rect 2810 4132 2818 4157
rect 1360 3980 1412 3989
rect 1360 3946 1373 3980
rect 1373 3946 1407 3980
rect 1407 3946 1412 3980
rect 1360 3937 1412 3946
rect 1424 3980 1476 3989
rect 1488 3980 1540 3989
rect 1552 3980 1604 3989
rect 1616 3980 1668 3989
rect 1680 3980 1732 3989
rect 1744 3980 1796 3989
rect 1808 3980 1860 3989
rect 1424 3946 1445 3980
rect 1445 3946 1476 3980
rect 1488 3946 1517 3980
rect 1517 3946 1540 3980
rect 1552 3946 1589 3980
rect 1589 3946 1604 3980
rect 1616 3946 1623 3980
rect 1623 3946 1661 3980
rect 1661 3946 1668 3980
rect 1680 3946 1695 3980
rect 1695 3946 1732 3980
rect 1744 3946 1767 3980
rect 1767 3946 1796 3980
rect 1808 3946 1839 3980
rect 1839 3946 1860 3980
rect 1424 3937 1476 3946
rect 1488 3937 1540 3946
rect 1552 3937 1604 3946
rect 1616 3937 1668 3946
rect 1680 3937 1732 3946
rect 1744 3937 1796 3946
rect 1808 3937 1860 3946
rect 1872 3980 1924 3989
rect 1872 3946 1877 3980
rect 1877 3946 1911 3980
rect 1911 3946 1924 3980
rect 1872 3937 1924 3946
rect 3756 3991 3808 4000
rect 3820 3991 3872 4000
rect 278 3805 332 3859
rect 3756 3957 3775 3991
rect 3775 3957 3808 3991
rect 3820 3957 3847 3991
rect 3847 3957 3872 3991
rect 3756 3948 3808 3957
rect 3820 3948 3872 3957
rect 3884 3991 3936 4000
rect 3884 3957 3885 3991
rect 3885 3957 3919 3991
rect 3919 3957 3936 3991
rect 3884 3948 3936 3957
rect 3948 3991 4000 4000
rect 3948 3957 3957 3991
rect 3957 3957 3991 3991
rect 3991 3957 4000 3991
rect 3948 3948 4000 3957
rect 4012 3991 4064 4000
rect 4012 3957 4029 3991
rect 4029 3957 4063 3991
rect 4063 3957 4064 3991
rect 4012 3948 4064 3957
rect 4076 3991 4128 4000
rect 4140 3991 4192 4000
rect 4076 3957 4101 3991
rect 4101 3957 4128 3991
rect 4140 3957 4173 3991
rect 4173 3957 4192 3991
rect 4076 3948 4128 3957
rect 4140 3948 4192 3957
rect 3565 3799 3617 3851
rect 4628 4298 4680 4307
rect 4628 4264 4637 4298
rect 4637 4264 4671 4298
rect 4671 4264 4680 4298
rect 4628 4255 4680 4264
rect 4862 4169 4914 4182
rect 4862 4135 4868 4169
rect 4868 4135 4902 4169
rect 4902 4135 4914 4169
rect 4862 4130 4914 4135
rect 4552 3999 4604 4051
rect 6868 4738 6920 4790
rect 6250 4412 6302 4464
rect 7194 4620 7246 4672
rect 6974 4410 7026 4462
rect 5117 4253 5169 4305
rect 5934 4286 5986 4296
rect 5934 4252 5942 4286
rect 5942 4252 5976 4286
rect 5976 4252 5986 4286
rect 5934 4244 5986 4252
rect 5015 4132 5067 4184
rect 5714 3992 5766 4000
rect 5778 3992 5830 4000
rect 5714 3958 5734 3992
rect 5734 3958 5766 3992
rect 5778 3958 5806 3992
rect 5806 3958 5830 3992
rect 5714 3948 5766 3958
rect 5778 3948 5830 3958
rect 5842 3992 5894 4000
rect 5842 3958 5844 3992
rect 5844 3958 5878 3992
rect 5878 3958 5894 3992
rect 5842 3948 5894 3958
rect 5906 3992 5958 4000
rect 5906 3958 5916 3992
rect 5916 3958 5950 3992
rect 5950 3958 5958 3992
rect 5906 3948 5958 3958
rect 5970 3992 6022 4000
rect 5970 3958 5988 3992
rect 5988 3958 6022 3992
rect 5970 3948 6022 3958
rect 6034 3992 6086 4000
rect 6098 3992 6150 4000
rect 6034 3958 6060 3992
rect 6060 3958 6086 3992
rect 6098 3958 6132 3992
rect 6132 3958 6150 3992
rect 6034 3948 6086 3958
rect 6098 3948 6150 3958
rect 5117 3799 5169 3851
rect 6586 4298 6638 4308
rect 6586 4264 6596 4298
rect 6596 4264 6630 4298
rect 6630 4264 6638 4298
rect 6586 4256 6638 4264
rect 6820 4170 6872 4182
rect 6820 4136 6826 4170
rect 6826 4136 6860 4170
rect 6860 4136 6872 4170
rect 6820 4130 6872 4136
rect 6510 4000 6562 4052
rect 6974 4132 7026 4184
rect 5035 3629 5087 3681
rect 6512 3714 6564 3766
rect 1398 3454 1450 3463
rect 1462 3454 1514 3463
rect 1398 3420 1417 3454
rect 1417 3420 1450 3454
rect 1462 3420 1489 3454
rect 1489 3420 1514 3454
rect 1398 3411 1450 3420
rect 1462 3411 1514 3420
rect 1526 3454 1578 3463
rect 1526 3420 1527 3454
rect 1527 3420 1561 3454
rect 1561 3420 1578 3454
rect 1526 3411 1578 3420
rect 1590 3454 1642 3463
rect 1590 3420 1599 3454
rect 1599 3420 1633 3454
rect 1633 3420 1642 3454
rect 1590 3411 1642 3420
rect 1654 3454 1706 3463
rect 1654 3420 1671 3454
rect 1671 3420 1705 3454
rect 1705 3420 1706 3454
rect 1654 3411 1706 3420
rect 1718 3454 1770 3463
rect 1782 3454 1834 3463
rect 1718 3420 1743 3454
rect 1743 3420 1770 3454
rect 1782 3420 1815 3454
rect 1815 3420 1834 3454
rect 1718 3411 1770 3420
rect 1782 3411 1834 3420
rect 560 3368 612 3392
rect 560 3340 566 3368
rect 566 3340 607 3368
rect 607 3340 612 3368
rect 702 3368 754 3388
rect 702 3336 710 3368
rect 710 3336 751 3368
rect 751 3336 754 3368
rect 378 3175 433 3230
rect 852 3186 904 3238
rect 378 2890 433 2945
rect 1004 3094 1056 3146
rect 1935 3105 1987 3157
rect 3776 3453 3828 3462
rect 3840 3453 3892 3462
rect 3904 3453 3956 3462
rect 3968 3453 4020 3462
rect 4032 3453 4084 3462
rect 4096 3453 4148 3462
rect 4160 3453 4212 3462
rect 3776 3419 3797 3453
rect 3797 3419 3828 3453
rect 3840 3419 3869 3453
rect 3869 3419 3892 3453
rect 3904 3419 3941 3453
rect 3941 3419 3956 3453
rect 3968 3419 3975 3453
rect 3975 3419 4013 3453
rect 4013 3419 4020 3453
rect 4032 3419 4047 3453
rect 4047 3419 4084 3453
rect 4096 3419 4119 3453
rect 4119 3419 4148 3453
rect 4160 3419 4191 3453
rect 4191 3419 4212 3453
rect 3776 3410 3828 3419
rect 3840 3410 3892 3419
rect 3904 3410 3956 3419
rect 3968 3410 4020 3419
rect 4032 3410 4084 3419
rect 4096 3410 4148 3419
rect 4160 3410 4212 3419
rect 2769 3296 2821 3348
rect 1155 3005 1207 3057
rect 1758 3047 1810 3056
rect 1758 3013 1773 3047
rect 1773 3013 1807 3047
rect 1807 3013 1810 3047
rect 1758 3004 1810 3013
rect 2270 3045 2322 3054
rect 2270 3011 2273 3045
rect 2273 3011 2307 3045
rect 2307 3011 2322 3045
rect 2270 3002 2322 3011
rect 3268 3219 3278 3243
rect 3278 3219 3312 3243
rect 3312 3219 3320 3243
rect 3268 3191 3320 3219
rect 4744 3510 4796 3562
rect 5734 3452 5786 3462
rect 5798 3452 5850 3462
rect 5862 3452 5914 3462
rect 5926 3452 5978 3462
rect 5990 3452 6042 3462
rect 6054 3452 6106 3462
rect 6118 3452 6170 3462
rect 5734 3418 5756 3452
rect 5756 3418 5786 3452
rect 5798 3418 5828 3452
rect 5828 3418 5850 3452
rect 5862 3418 5900 3452
rect 5900 3418 5914 3452
rect 5926 3418 5934 3452
rect 5934 3418 5972 3452
rect 5972 3418 5978 3452
rect 5990 3418 6006 3452
rect 6006 3418 6042 3452
rect 6054 3418 6078 3452
rect 6078 3418 6106 3452
rect 6118 3418 6150 3452
rect 6150 3418 6170 3452
rect 5734 3410 5786 3418
rect 5798 3410 5850 3418
rect 5862 3410 5914 3418
rect 5926 3410 5978 3418
rect 5990 3410 6042 3418
rect 6054 3410 6106 3418
rect 6118 3410 6170 3418
rect 4292 3183 4344 3235
rect 5016 3182 5068 3234
rect 1248 2894 1300 2946
rect 378 2790 434 2846
rect 2020 2929 2072 2946
rect 2020 2895 2030 2929
rect 2030 2895 2064 2929
rect 2064 2895 2072 2929
rect 2020 2894 2072 2895
rect 2522 2929 2574 2944
rect 2522 2895 2530 2929
rect 2530 2895 2564 2929
rect 2564 2895 2574 2929
rect 2522 2892 2574 2895
rect 2842 3043 2894 3052
rect 2842 3009 2857 3043
rect 2857 3009 2891 3043
rect 2891 3009 2894 3043
rect 2842 3000 2894 3009
rect 3268 2998 3320 3050
rect 3561 3025 3613 3077
rect 3976 3058 4028 3068
rect 3976 3024 3984 3058
rect 3984 3024 4018 3058
rect 4018 3024 4028 3058
rect 3976 3016 4028 3024
rect 2766 2929 2818 2956
rect 2766 2904 2776 2929
rect 2776 2904 2810 2929
rect 2810 2904 2818 2929
rect 1360 2752 1412 2761
rect 1360 2718 1373 2752
rect 1373 2718 1407 2752
rect 1407 2718 1412 2752
rect 1360 2709 1412 2718
rect 1424 2752 1476 2761
rect 1488 2752 1540 2761
rect 1552 2752 1604 2761
rect 1616 2752 1668 2761
rect 1680 2752 1732 2761
rect 1744 2752 1796 2761
rect 1808 2752 1860 2761
rect 1424 2718 1445 2752
rect 1445 2718 1476 2752
rect 1488 2718 1517 2752
rect 1517 2718 1540 2752
rect 1552 2718 1589 2752
rect 1589 2718 1604 2752
rect 1616 2718 1623 2752
rect 1623 2718 1661 2752
rect 1661 2718 1668 2752
rect 1680 2718 1695 2752
rect 1695 2718 1732 2752
rect 1744 2718 1767 2752
rect 1767 2718 1796 2752
rect 1808 2718 1839 2752
rect 1839 2718 1860 2752
rect 1424 2709 1476 2718
rect 1488 2709 1540 2718
rect 1552 2709 1604 2718
rect 1616 2709 1668 2718
rect 1680 2709 1732 2718
rect 1744 2709 1796 2718
rect 1808 2709 1860 2718
rect 1872 2752 1924 2761
rect 1872 2718 1877 2752
rect 1877 2718 1911 2752
rect 1911 2718 1924 2752
rect 1872 2709 1924 2718
rect 3756 2763 3808 2772
rect 3820 2763 3872 2772
rect 278 2577 332 2631
rect 3756 2729 3775 2763
rect 3775 2729 3808 2763
rect 3820 2729 3847 2763
rect 3847 2729 3872 2763
rect 3756 2720 3808 2729
rect 3820 2720 3872 2729
rect 3884 2763 3936 2772
rect 3884 2729 3885 2763
rect 3885 2729 3919 2763
rect 3919 2729 3936 2763
rect 3884 2720 3936 2729
rect 3948 2763 4000 2772
rect 3948 2729 3957 2763
rect 3957 2729 3991 2763
rect 3991 2729 4000 2763
rect 3948 2720 4000 2729
rect 4012 2763 4064 2772
rect 4012 2729 4029 2763
rect 4029 2729 4063 2763
rect 4063 2729 4064 2763
rect 4012 2720 4064 2729
rect 4076 2763 4128 2772
rect 4140 2763 4192 2772
rect 4076 2729 4101 2763
rect 4101 2729 4128 2763
rect 4140 2729 4173 2763
rect 4173 2729 4192 2763
rect 4076 2720 4128 2729
rect 4140 2720 4192 2729
rect 3565 2571 3617 2623
rect 4628 3070 4680 3079
rect 4628 3036 4637 3070
rect 4637 3036 4671 3070
rect 4671 3036 4680 3070
rect 4628 3027 4680 3036
rect 4862 2941 4914 2954
rect 4862 2907 4868 2941
rect 4868 2907 4902 2941
rect 4902 2907 4914 2941
rect 4862 2902 4914 2907
rect 4552 2771 4604 2823
rect 6843 3510 6895 3562
rect 6250 3184 6302 3236
rect 6974 3182 7026 3234
rect 5197 3025 5249 3077
rect 5934 3058 5986 3068
rect 5934 3024 5942 3058
rect 5942 3024 5976 3058
rect 5976 3024 5986 3058
rect 5934 3016 5986 3024
rect 5015 2904 5067 2956
rect 5714 2764 5766 2772
rect 5778 2764 5830 2772
rect 5714 2730 5734 2764
rect 5734 2730 5766 2764
rect 5778 2730 5806 2764
rect 5806 2730 5830 2764
rect 5714 2720 5766 2730
rect 5778 2720 5830 2730
rect 5842 2764 5894 2772
rect 5842 2730 5844 2764
rect 5844 2730 5878 2764
rect 5878 2730 5894 2764
rect 5842 2720 5894 2730
rect 5906 2764 5958 2772
rect 5906 2730 5916 2764
rect 5916 2730 5950 2764
rect 5950 2730 5958 2764
rect 5906 2720 5958 2730
rect 5970 2764 6022 2772
rect 5970 2730 5988 2764
rect 5988 2730 6022 2764
rect 5970 2720 6022 2730
rect 6034 2764 6086 2772
rect 6098 2764 6150 2772
rect 6034 2730 6060 2764
rect 6060 2730 6086 2764
rect 6098 2730 6132 2764
rect 6132 2730 6150 2764
rect 6034 2720 6086 2730
rect 6098 2720 6150 2730
rect 5197 2571 5249 2623
rect 6586 3070 6638 3080
rect 6586 3036 6596 3070
rect 6596 3036 6630 3070
rect 6630 3036 6638 3070
rect 6586 3028 6638 3036
rect 6820 2942 6872 2954
rect 6820 2908 6826 2942
rect 6826 2908 6860 2942
rect 6860 2908 6872 2942
rect 6820 2902 6872 2908
rect 6510 2772 6562 2824
rect 6974 2904 7026 2956
rect 7107 2484 7159 2536
rect 1398 2226 1450 2235
rect 1462 2226 1514 2235
rect 1398 2192 1417 2226
rect 1417 2192 1450 2226
rect 1462 2192 1489 2226
rect 1489 2192 1514 2226
rect 1398 2183 1450 2192
rect 1462 2183 1514 2192
rect 1526 2226 1578 2235
rect 1526 2192 1527 2226
rect 1527 2192 1561 2226
rect 1561 2192 1578 2226
rect 1526 2183 1578 2192
rect 1590 2226 1642 2235
rect 1590 2192 1599 2226
rect 1599 2192 1633 2226
rect 1633 2192 1642 2226
rect 1590 2183 1642 2192
rect 1654 2226 1706 2235
rect 1654 2192 1671 2226
rect 1671 2192 1705 2226
rect 1705 2192 1706 2226
rect 1654 2183 1706 2192
rect 1718 2226 1770 2235
rect 1782 2226 1834 2235
rect 1718 2192 1743 2226
rect 1743 2192 1770 2226
rect 1782 2192 1815 2226
rect 1815 2192 1834 2226
rect 1718 2183 1770 2192
rect 1782 2183 1834 2192
rect 560 2140 612 2164
rect 560 2112 566 2140
rect 566 2112 607 2140
rect 607 2112 612 2140
rect 702 2140 754 2160
rect 702 2108 710 2140
rect 710 2108 751 2140
rect 751 2108 754 2140
rect 378 1947 433 2002
rect 852 1958 904 2010
rect 378 1662 433 1717
rect 1004 1866 1056 1918
rect 1935 1877 1987 1929
rect 3776 2225 3828 2234
rect 3840 2225 3892 2234
rect 3904 2225 3956 2234
rect 3968 2225 4020 2234
rect 4032 2225 4084 2234
rect 4096 2225 4148 2234
rect 4160 2225 4212 2234
rect 3776 2191 3797 2225
rect 3797 2191 3828 2225
rect 3840 2191 3869 2225
rect 3869 2191 3892 2225
rect 3904 2191 3941 2225
rect 3941 2191 3956 2225
rect 3968 2191 3975 2225
rect 3975 2191 4013 2225
rect 4013 2191 4020 2225
rect 4032 2191 4047 2225
rect 4047 2191 4084 2225
rect 4096 2191 4119 2225
rect 4119 2191 4148 2225
rect 4160 2191 4191 2225
rect 4191 2191 4212 2225
rect 3776 2182 3828 2191
rect 3840 2182 3892 2191
rect 3904 2182 3956 2191
rect 3968 2182 4020 2191
rect 4032 2182 4084 2191
rect 4096 2182 4148 2191
rect 4160 2182 4212 2191
rect 2769 2068 2821 2120
rect 1155 1777 1207 1829
rect 1758 1819 1810 1828
rect 1758 1785 1773 1819
rect 1773 1785 1807 1819
rect 1807 1785 1810 1819
rect 1758 1776 1810 1785
rect 2270 1817 2322 1826
rect 2270 1783 2273 1817
rect 2273 1783 2307 1817
rect 2307 1783 2322 1817
rect 2270 1774 2322 1783
rect 3268 1991 3278 2015
rect 3278 1991 3312 2015
rect 3312 1991 3320 2015
rect 3268 1963 3320 1991
rect 4744 2282 4796 2334
rect 5029 2364 5081 2416
rect 5734 2224 5786 2234
rect 5798 2224 5850 2234
rect 5862 2224 5914 2234
rect 5926 2224 5978 2234
rect 5990 2224 6042 2234
rect 6054 2224 6106 2234
rect 6118 2224 6170 2234
rect 5734 2190 5756 2224
rect 5756 2190 5786 2224
rect 5798 2190 5828 2224
rect 5828 2190 5850 2224
rect 5862 2190 5900 2224
rect 5900 2190 5914 2224
rect 5926 2190 5934 2224
rect 5934 2190 5972 2224
rect 5972 2190 5978 2224
rect 5990 2190 6006 2224
rect 6006 2190 6042 2224
rect 6054 2190 6078 2224
rect 6078 2190 6106 2224
rect 6118 2190 6150 2224
rect 6150 2190 6170 2224
rect 5734 2182 5786 2190
rect 5798 2182 5850 2190
rect 5862 2182 5914 2190
rect 5926 2182 5978 2190
rect 5990 2182 6042 2190
rect 6054 2182 6106 2190
rect 6118 2182 6170 2190
rect 4292 1955 4344 2007
rect 5016 1954 5068 2006
rect 1248 1666 1300 1718
rect 378 1562 434 1618
rect 2020 1701 2072 1718
rect 2020 1667 2030 1701
rect 2030 1667 2064 1701
rect 2064 1667 2072 1701
rect 2020 1666 2072 1667
rect 2522 1701 2574 1716
rect 2522 1667 2530 1701
rect 2530 1667 2564 1701
rect 2564 1667 2574 1701
rect 2522 1664 2574 1667
rect 2842 1815 2894 1824
rect 2842 1781 2857 1815
rect 2857 1781 2891 1815
rect 2891 1781 2894 1815
rect 2842 1772 2894 1781
rect 3268 1770 3320 1822
rect 3561 1797 3613 1849
rect 3976 1830 4028 1840
rect 3976 1796 3984 1830
rect 3984 1796 4018 1830
rect 4018 1796 4028 1830
rect 3976 1788 4028 1796
rect 2766 1701 2818 1728
rect 2766 1676 2776 1701
rect 2776 1676 2810 1701
rect 2810 1676 2818 1701
rect 1360 1524 1412 1533
rect 1360 1490 1373 1524
rect 1373 1490 1407 1524
rect 1407 1490 1412 1524
rect 1360 1481 1412 1490
rect 1424 1524 1476 1533
rect 1488 1524 1540 1533
rect 1552 1524 1604 1533
rect 1616 1524 1668 1533
rect 1680 1524 1732 1533
rect 1744 1524 1796 1533
rect 1808 1524 1860 1533
rect 1424 1490 1445 1524
rect 1445 1490 1476 1524
rect 1488 1490 1517 1524
rect 1517 1490 1540 1524
rect 1552 1490 1589 1524
rect 1589 1490 1604 1524
rect 1616 1490 1623 1524
rect 1623 1490 1661 1524
rect 1661 1490 1668 1524
rect 1680 1490 1695 1524
rect 1695 1490 1732 1524
rect 1744 1490 1767 1524
rect 1767 1490 1796 1524
rect 1808 1490 1839 1524
rect 1839 1490 1860 1524
rect 1424 1481 1476 1490
rect 1488 1481 1540 1490
rect 1552 1481 1604 1490
rect 1616 1481 1668 1490
rect 1680 1481 1732 1490
rect 1744 1481 1796 1490
rect 1808 1481 1860 1490
rect 1872 1524 1924 1533
rect 1872 1490 1877 1524
rect 1877 1490 1911 1524
rect 1911 1490 1924 1524
rect 1872 1481 1924 1490
rect 3756 1535 3808 1544
rect 3820 1535 3872 1544
rect 278 1349 332 1403
rect 3756 1501 3775 1535
rect 3775 1501 3808 1535
rect 3820 1501 3847 1535
rect 3847 1501 3872 1535
rect 3756 1492 3808 1501
rect 3820 1492 3872 1501
rect 3884 1535 3936 1544
rect 3884 1501 3885 1535
rect 3885 1501 3919 1535
rect 3919 1501 3936 1535
rect 3884 1492 3936 1501
rect 3948 1535 4000 1544
rect 3948 1501 3957 1535
rect 3957 1501 3991 1535
rect 3991 1501 4000 1535
rect 3948 1492 4000 1501
rect 4012 1535 4064 1544
rect 4012 1501 4029 1535
rect 4029 1501 4063 1535
rect 4063 1501 4064 1535
rect 4012 1492 4064 1501
rect 4076 1535 4128 1544
rect 4140 1535 4192 1544
rect 4076 1501 4101 1535
rect 4101 1501 4128 1535
rect 4140 1501 4173 1535
rect 4173 1501 4192 1535
rect 4076 1492 4128 1501
rect 4140 1492 4192 1501
rect 3565 1343 3617 1395
rect 4628 1842 4680 1851
rect 4628 1808 4637 1842
rect 4637 1808 4671 1842
rect 4671 1808 4680 1842
rect 4628 1799 4680 1808
rect 4862 1713 4914 1726
rect 4862 1679 4868 1713
rect 4868 1679 4902 1713
rect 4902 1679 4914 1713
rect 4862 1674 4914 1679
rect 4552 1543 4604 1595
rect 6868 2282 6920 2334
rect 6250 1956 6302 2008
rect 6974 1954 7026 2006
rect 5117 1797 5169 1849
rect 5934 1830 5986 1840
rect 5934 1796 5942 1830
rect 5942 1796 5976 1830
rect 5976 1796 5986 1830
rect 5934 1788 5986 1796
rect 5015 1676 5067 1728
rect 5714 1536 5766 1544
rect 5778 1536 5830 1544
rect 5714 1502 5734 1536
rect 5734 1502 5766 1536
rect 5778 1502 5806 1536
rect 5806 1502 5830 1536
rect 5714 1492 5766 1502
rect 5778 1492 5830 1502
rect 5842 1536 5894 1544
rect 5842 1502 5844 1536
rect 5844 1502 5878 1536
rect 5878 1502 5894 1536
rect 5842 1492 5894 1502
rect 5906 1536 5958 1544
rect 5906 1502 5916 1536
rect 5916 1502 5950 1536
rect 5950 1502 5958 1536
rect 5906 1492 5958 1502
rect 5970 1536 6022 1544
rect 5970 1502 5988 1536
rect 5988 1502 6022 1536
rect 5970 1492 6022 1502
rect 6034 1536 6086 1544
rect 6098 1536 6150 1544
rect 6034 1502 6060 1536
rect 6060 1502 6086 1536
rect 6098 1502 6132 1536
rect 6132 1502 6150 1536
rect 6034 1492 6086 1502
rect 6098 1492 6150 1502
rect 5117 1343 5169 1395
rect 6586 1842 6638 1852
rect 6586 1808 6596 1842
rect 6596 1808 6630 1842
rect 6630 1808 6638 1842
rect 6586 1800 6638 1808
rect 6820 1714 6872 1726
rect 6820 1680 6826 1714
rect 6826 1680 6860 1714
rect 6860 1680 6872 1714
rect 6820 1674 6872 1680
rect 6510 1544 6562 1596
rect 6974 1676 7026 1728
rect 5035 1173 5087 1225
rect 1398 998 1450 1007
rect 1462 998 1514 1007
rect 1398 964 1417 998
rect 1417 964 1450 998
rect 1462 964 1489 998
rect 1489 964 1514 998
rect 1398 955 1450 964
rect 1462 955 1514 964
rect 1526 998 1578 1007
rect 1526 964 1527 998
rect 1527 964 1561 998
rect 1561 964 1578 998
rect 1526 955 1578 964
rect 1590 998 1642 1007
rect 1590 964 1599 998
rect 1599 964 1633 998
rect 1633 964 1642 998
rect 1590 955 1642 964
rect 1654 998 1706 1007
rect 1654 964 1671 998
rect 1671 964 1705 998
rect 1705 964 1706 998
rect 1654 955 1706 964
rect 1718 998 1770 1007
rect 1782 998 1834 1007
rect 1718 964 1743 998
rect 1743 964 1770 998
rect 1782 964 1815 998
rect 1815 964 1834 998
rect 1718 955 1770 964
rect 1782 955 1834 964
rect 560 912 612 936
rect 560 884 566 912
rect 566 884 607 912
rect 607 884 612 912
rect 702 912 754 932
rect 702 880 710 912
rect 710 880 751 912
rect 751 880 754 912
rect 378 719 433 774
rect 852 730 904 782
rect 378 434 433 489
rect 1004 638 1056 690
rect 1935 649 1987 701
rect 3776 997 3828 1006
rect 3840 997 3892 1006
rect 3904 997 3956 1006
rect 3968 997 4020 1006
rect 4032 997 4084 1006
rect 4096 997 4148 1006
rect 4160 997 4212 1006
rect 3776 963 3797 997
rect 3797 963 3828 997
rect 3840 963 3869 997
rect 3869 963 3892 997
rect 3904 963 3941 997
rect 3941 963 3956 997
rect 3968 963 3975 997
rect 3975 963 4013 997
rect 4013 963 4020 997
rect 4032 963 4047 997
rect 4047 963 4084 997
rect 4096 963 4119 997
rect 4119 963 4148 997
rect 4160 963 4191 997
rect 4191 963 4212 997
rect 3776 954 3828 963
rect 3840 954 3892 963
rect 3904 954 3956 963
rect 3968 954 4020 963
rect 4032 954 4084 963
rect 4096 954 4148 963
rect 4160 954 4212 963
rect 2769 840 2821 892
rect 1155 549 1207 601
rect 1758 591 1810 600
rect 1758 557 1773 591
rect 1773 557 1807 591
rect 1807 557 1810 591
rect 1758 548 1810 557
rect 2270 589 2322 598
rect 2270 555 2273 589
rect 2273 555 2307 589
rect 2307 555 2322 589
rect 2270 546 2322 555
rect 3268 763 3278 787
rect 3278 763 3312 787
rect 3312 763 3320 787
rect 3268 735 3320 763
rect 4744 1054 4796 1106
rect 4292 727 4344 779
rect 5016 726 5068 778
rect 1248 438 1300 490
rect 378 334 434 390
rect 2020 473 2072 490
rect 2020 439 2030 473
rect 2030 439 2064 473
rect 2064 439 2072 473
rect 2020 438 2072 439
rect 2522 473 2574 488
rect 2522 439 2530 473
rect 2530 439 2564 473
rect 2564 439 2574 473
rect 2522 436 2574 439
rect 2842 587 2894 596
rect 2842 553 2857 587
rect 2857 553 2891 587
rect 2891 553 2894 587
rect 2842 544 2894 553
rect 3268 542 3320 594
rect 3561 569 3613 621
rect 3976 602 4028 612
rect 3976 568 3984 602
rect 3984 568 4018 602
rect 4018 568 4028 602
rect 3976 560 4028 568
rect 2766 473 2818 500
rect 2766 448 2776 473
rect 2776 448 2810 473
rect 2810 448 2818 473
rect 1360 296 1412 305
rect 1360 262 1373 296
rect 1373 262 1407 296
rect 1407 262 1412 296
rect 1360 253 1412 262
rect 1424 296 1476 305
rect 1488 296 1540 305
rect 1552 296 1604 305
rect 1616 296 1668 305
rect 1680 296 1732 305
rect 1744 296 1796 305
rect 1808 296 1860 305
rect 1424 262 1445 296
rect 1445 262 1476 296
rect 1488 262 1517 296
rect 1517 262 1540 296
rect 1552 262 1589 296
rect 1589 262 1604 296
rect 1616 262 1623 296
rect 1623 262 1661 296
rect 1661 262 1668 296
rect 1680 262 1695 296
rect 1695 262 1732 296
rect 1744 262 1767 296
rect 1767 262 1796 296
rect 1808 262 1839 296
rect 1839 262 1860 296
rect 1424 253 1476 262
rect 1488 253 1540 262
rect 1552 253 1604 262
rect 1616 253 1668 262
rect 1680 253 1732 262
rect 1744 253 1796 262
rect 1808 253 1860 262
rect 1872 296 1924 305
rect 1872 262 1877 296
rect 1877 262 1911 296
rect 1911 262 1924 296
rect 1872 253 1924 262
rect 3756 307 3808 316
rect 3820 307 3872 316
rect 278 121 332 175
rect 3756 273 3775 307
rect 3775 273 3808 307
rect 3820 273 3847 307
rect 3847 273 3872 307
rect 3756 264 3808 273
rect 3820 264 3872 273
rect 3884 307 3936 316
rect 3884 273 3885 307
rect 3885 273 3919 307
rect 3919 273 3936 307
rect 3884 264 3936 273
rect 3948 307 4000 316
rect 3948 273 3957 307
rect 3957 273 3991 307
rect 3991 273 4000 307
rect 3948 264 4000 273
rect 4012 307 4064 316
rect 4012 273 4029 307
rect 4029 273 4063 307
rect 4063 273 4064 307
rect 4012 264 4064 273
rect 4076 307 4128 316
rect 4140 307 4192 316
rect 4076 273 4101 307
rect 4101 273 4128 307
rect 4140 273 4173 307
rect 4173 273 4192 307
rect 4076 264 4128 273
rect 4140 264 4192 273
rect 3565 115 3617 167
rect 4628 614 4680 623
rect 4628 580 4637 614
rect 4637 580 4671 614
rect 4671 580 4680 614
rect 4628 571 4680 580
rect 4862 485 4914 498
rect 4862 451 4868 485
rect 4868 451 4902 485
rect 4902 451 4914 485
rect 4862 446 4914 451
rect 4552 315 4604 367
rect 5015 448 5067 500
<< metal2 >>
rect 42 19426 110 19435
rect 42 18220 110 19358
rect 274 19023 329 19648
rect 378 19194 433 19648
rect 1348 19429 1880 19470
rect 1348 19373 1388 19429
rect 1444 19427 1468 19429
rect 1524 19427 1548 19429
rect 1604 19427 1628 19429
rect 1684 19427 1708 19429
rect 1764 19427 1788 19429
rect 1450 19375 1462 19427
rect 1524 19375 1526 19427
rect 1706 19375 1708 19427
rect 1770 19375 1782 19427
rect 1444 19373 1468 19375
rect 1524 19373 1548 19375
rect 1604 19373 1628 19375
rect 1684 19373 1708 19375
rect 1764 19373 1788 19375
rect 1844 19373 1880 19429
rect 560 19356 612 19362
rect 700 19354 756 19360
rect 612 19352 976 19354
rect 612 19304 702 19352
rect 560 19300 702 19304
rect 754 19300 976 19352
rect 1348 19330 1880 19373
rect 2759 19312 2827 19320
rect 560 19298 1268 19300
rect 700 19292 756 19298
rect 920 19292 1268 19298
rect 2759 19292 2769 19312
rect 920 19260 2769 19292
rect 2821 19260 2827 19312
rect 920 19248 2827 19260
rect 920 19244 1268 19248
rect 852 19202 904 19208
rect 372 19139 378 19194
rect 433 19139 439 19194
rect 1396 19203 2851 19212
rect 3268 19207 3320 19213
rect 1396 19198 3268 19203
rect 904 19168 3268 19198
rect 904 19154 1440 19168
rect 2851 19159 3268 19168
rect 852 19144 904 19150
rect 3268 19149 3320 19155
rect 1930 19122 1990 19133
rect 1004 19110 1056 19116
rect 1930 19111 1932 19122
rect 1056 19099 1242 19106
rect 1599 19099 1932 19111
rect 1056 19077 1932 19099
rect 1056 19065 1633 19077
rect 1930 19066 1932 19077
rect 1988 19111 1990 19122
rect 1988 19077 1991 19111
rect 1988 19066 1990 19077
rect 1056 19062 1242 19065
rect 1004 19052 1056 19058
rect 1930 19055 1990 19066
rect 3564 19047 3605 19648
rect 5023 19556 5029 19608
rect 5081 19556 5087 19608
rect 5122 19560 5163 19648
rect 5202 19560 5243 19648
rect 5282 19560 5323 19648
rect 5362 19560 5403 19648
rect 5442 19560 5483 19648
rect 5522 19560 5563 19648
rect 4744 19526 4796 19532
rect 5036 19520 5075 19556
rect 4796 19481 5075 19520
rect 3724 19428 4264 19470
rect 4744 19468 4796 19474
rect 3724 19372 3766 19428
rect 3822 19426 3846 19428
rect 3902 19426 3926 19428
rect 3982 19426 4006 19428
rect 4062 19426 4086 19428
rect 4142 19426 4166 19428
rect 3828 19374 3840 19426
rect 3902 19374 3904 19426
rect 4084 19374 4086 19426
rect 4148 19374 4160 19426
rect 3822 19372 3846 19374
rect 3902 19372 3926 19374
rect 3982 19372 4006 19374
rect 4062 19372 4086 19374
rect 4142 19372 4166 19374
rect 4222 19372 4264 19428
rect 3724 19330 4264 19372
rect 4291 19201 4346 19207
rect 5016 19201 5068 19204
rect 4291 19199 5084 19201
rect 4291 19147 4292 19199
rect 4344 19198 5084 19199
rect 4344 19147 5016 19198
rect 4291 19146 5016 19147
rect 5068 19146 5084 19198
rect 4291 19140 4346 19146
rect 5016 19140 5068 19146
rect 5122 19047 5164 19560
rect 3561 19041 3613 19047
rect 1154 19023 1209 19029
rect 274 19021 1209 19023
rect 274 18969 1155 19021
rect 1207 18969 1209 19021
rect 274 18968 1209 18969
rect 1154 18962 1209 18968
rect 1754 19024 1814 19030
rect 2267 19024 2325 19033
rect 1754 19021 2325 19024
rect 2838 19021 2898 19026
rect 1754 19020 2898 19021
rect 1754 18968 1758 19020
rect 1810 19018 2908 19020
rect 1810 18968 2270 19018
rect 1754 18966 2270 18968
rect 2322 19016 2908 19018
rect 2322 18966 2842 19016
rect 1754 18964 2842 18966
rect 2894 18964 2908 19016
rect 1754 18958 1814 18964
rect 2267 18963 2908 18964
rect 2267 18951 2325 18963
rect 2838 18960 2908 18963
rect 3262 18962 3268 19014
rect 3320 18962 3326 19014
rect 3976 19032 4028 19038
rect 3561 18983 3613 18989
rect 3975 18983 3976 19026
rect 2838 18954 2898 18960
rect 2768 18920 2816 18924
rect 378 18909 433 18915
rect 1248 18910 1300 18916
rect 433 18906 619 18909
rect 433 18862 1248 18906
rect 433 18854 619 18862
rect 2020 18910 2072 18916
rect 2522 18912 2574 18914
rect 1300 18862 2020 18906
rect 378 18848 433 18854
rect 1248 18852 1300 18858
rect 2020 18852 2072 18858
rect 2509 18910 2587 18912
rect 2509 18854 2520 18910
rect 2576 18854 2587 18910
rect 2760 18868 2766 18920
rect 2818 18916 2824 18920
rect 3270 18916 3314 18962
rect 3564 18944 3605 18983
rect 4622 18991 4628 19043
rect 4680 18991 4686 19043
rect 5117 19041 5169 19047
rect 3976 18974 4028 18980
rect 2818 18872 3314 18916
rect 3979 18927 4018 18974
rect 4637 18927 4671 18991
rect 5117 18983 5169 18989
rect 5122 18944 5164 18983
rect 5202 18944 5244 19560
rect 5282 18944 5324 19560
rect 5362 18944 5404 19560
rect 5442 18944 5484 19560
rect 5522 18944 5564 19560
rect 6868 19526 6920 19532
rect 6920 19481 7147 19520
rect 5682 19428 6222 19470
rect 6868 19468 6920 19474
rect 5682 19372 5724 19428
rect 5780 19426 5804 19428
rect 5860 19426 5884 19428
rect 5940 19426 5964 19428
rect 6020 19426 6044 19428
rect 6100 19426 6124 19428
rect 5786 19374 5798 19426
rect 5860 19374 5862 19426
rect 6042 19374 6044 19426
rect 6106 19374 6118 19426
rect 5780 19372 5804 19374
rect 5860 19372 5884 19374
rect 5940 19372 5964 19374
rect 6020 19372 6044 19374
rect 6100 19372 6124 19374
rect 6180 19372 6222 19428
rect 5682 19330 6222 19372
rect 6250 19202 6304 19208
rect 6974 19202 7026 19204
rect 6250 19200 7042 19202
rect 6302 19198 7042 19200
rect 6302 19148 6974 19198
rect 6250 19146 6974 19148
rect 7026 19146 7042 19198
rect 6250 19140 6304 19146
rect 6974 19140 7026 19146
rect 5934 19032 5986 19038
rect 6580 18992 6586 19044
rect 6638 18992 6644 19044
rect 5934 18974 5986 18980
rect 3979 18888 4673 18927
rect 4862 18918 4914 18924
rect 2818 18868 2824 18872
rect 2509 18852 2587 18854
rect 2522 18850 2574 18852
rect 2768 18828 2812 18868
rect 5015 18920 5067 18926
rect 4914 18878 5015 18907
rect 42 16970 110 18152
rect 42 15764 110 16902
rect 42 14514 110 15696
rect 42 13308 110 14446
rect 42 12058 110 13240
rect 42 10852 110 11990
rect 42 9602 110 10784
rect 42 8396 110 9534
rect 42 7146 110 8328
rect 42 5940 110 7078
rect 42 4690 110 5872
rect 42 3484 110 4622
rect 42 2234 110 3416
rect 42 1028 110 2166
rect 42 951 110 960
rect 144 18750 212 18759
rect 144 17514 212 18682
rect 274 18601 329 18790
rect 372 18754 378 18810
rect 434 18754 440 18810
rect 274 18595 332 18601
rect 274 18541 278 18595
rect 277 18420 332 18541
rect 378 18582 434 18754
rect 1324 18727 1960 18780
rect 1324 18725 1374 18727
rect 1430 18725 1454 18727
rect 1510 18725 1534 18727
rect 1590 18725 1614 18727
rect 1670 18725 1694 18727
rect 1750 18725 1774 18727
rect 1830 18725 1854 18727
rect 1910 18725 1960 18727
rect 1324 18673 1360 18725
rect 1604 18673 1614 18725
rect 1670 18673 1680 18725
rect 1924 18673 1960 18725
rect 1324 18671 1374 18673
rect 1430 18671 1454 18673
rect 1510 18671 1534 18673
rect 1590 18671 1614 18673
rect 1670 18671 1694 18673
rect 1750 18671 1774 18673
rect 1830 18671 1854 18673
rect 1910 18671 1960 18673
rect 1324 18640 1960 18671
rect 3564 18593 3605 18864
rect 4862 18860 4914 18866
rect 5015 18862 5067 18868
rect 5202 18864 5243 18944
rect 5282 18864 5323 18944
rect 5362 18864 5403 18944
rect 5442 18864 5483 18944
rect 5522 18864 5563 18944
rect 5938 18928 5976 18974
rect 6596 18928 6630 18992
rect 5938 18888 6632 18928
rect 6820 18918 6872 18924
rect 6974 18920 7026 18926
rect 6872 18878 6974 18908
rect 3704 18738 4244 18780
rect 3704 18682 3746 18738
rect 3802 18736 3826 18738
rect 3882 18736 3906 18738
rect 3962 18736 3986 18738
rect 4042 18736 4066 18738
rect 4122 18736 4146 18738
rect 3808 18684 3820 18736
rect 3882 18684 3884 18736
rect 4064 18684 4066 18736
rect 4128 18684 4140 18736
rect 3802 18682 3826 18684
rect 3882 18682 3906 18684
rect 3962 18682 3986 18684
rect 4042 18682 4066 18684
rect 4122 18682 4146 18684
rect 4202 18682 4244 18738
rect 4546 18735 4552 18787
rect 4604 18735 4610 18787
rect 3704 18640 4244 18682
rect 3564 18587 3617 18593
rect 274 17795 329 18420
rect 378 17966 433 18582
rect 3564 18535 3565 18587
rect 4559 18571 4598 18735
rect 5122 18593 5164 18864
rect 5117 18587 5169 18593
rect 3564 18529 3617 18535
rect 5117 18529 5169 18535
rect 1348 18201 1880 18242
rect 1348 18145 1388 18201
rect 1444 18199 1468 18201
rect 1524 18199 1548 18201
rect 1604 18199 1628 18201
rect 1684 18199 1708 18201
rect 1764 18199 1788 18201
rect 1450 18147 1462 18199
rect 1524 18147 1526 18199
rect 1706 18147 1708 18199
rect 1770 18147 1782 18199
rect 1444 18145 1468 18147
rect 1524 18145 1548 18147
rect 1604 18145 1628 18147
rect 1684 18145 1708 18147
rect 1764 18145 1788 18147
rect 1844 18145 1880 18201
rect 560 18128 612 18134
rect 700 18126 756 18132
rect 612 18124 976 18126
rect 612 18076 702 18124
rect 560 18072 702 18076
rect 754 18072 976 18124
rect 1348 18102 1880 18145
rect 2759 18084 2827 18092
rect 560 18070 1268 18072
rect 700 18064 756 18070
rect 920 18064 1268 18070
rect 2759 18064 2769 18084
rect 920 18032 2769 18064
rect 2821 18032 2827 18084
rect 920 18020 2827 18032
rect 920 18016 1268 18020
rect 852 17974 904 17980
rect 372 17911 378 17966
rect 433 17911 439 17966
rect 1396 17975 2851 17984
rect 3268 17979 3320 17985
rect 1396 17970 3268 17975
rect 904 17940 3268 17970
rect 904 17926 1440 17940
rect 2851 17931 3268 17940
rect 852 17916 904 17922
rect 3268 17921 3320 17927
rect 1930 17894 1990 17905
rect 1004 17882 1056 17888
rect 1930 17883 1932 17894
rect 1056 17871 1242 17878
rect 1599 17871 1932 17883
rect 1056 17849 1932 17871
rect 1056 17837 1633 17849
rect 1930 17838 1932 17849
rect 1988 17883 1990 17894
rect 1988 17849 1991 17883
rect 1988 17838 1990 17849
rect 1056 17834 1242 17837
rect 1004 17824 1056 17830
rect 1930 17827 1990 17838
rect 3564 17819 3605 18529
rect 5029 18365 5035 18417
rect 5087 18365 5093 18417
rect 4744 18298 4796 18304
rect 5047 18292 5075 18365
rect 4796 18253 5075 18292
rect 3724 18200 4264 18242
rect 4744 18240 4796 18246
rect 3724 18144 3766 18200
rect 3822 18198 3846 18200
rect 3902 18198 3926 18200
rect 3982 18198 4006 18200
rect 4062 18198 4086 18200
rect 4142 18198 4166 18200
rect 3828 18146 3840 18198
rect 3902 18146 3904 18198
rect 4084 18146 4086 18198
rect 4148 18146 4160 18198
rect 3822 18144 3846 18146
rect 3902 18144 3926 18146
rect 3982 18144 4006 18146
rect 4062 18144 4086 18146
rect 4142 18144 4166 18146
rect 4222 18144 4264 18200
rect 3724 18102 4264 18144
rect 4291 17973 4346 17979
rect 5016 17973 5068 17976
rect 4291 17971 5084 17973
rect 4291 17919 4292 17971
rect 4344 17970 5084 17971
rect 4344 17919 5016 17970
rect 4291 17918 5016 17919
rect 5068 17918 5084 17970
rect 4291 17912 4346 17918
rect 5016 17912 5068 17918
rect 3561 17813 3613 17819
rect 1154 17795 1209 17801
rect 274 17793 1209 17795
rect 274 17741 1155 17793
rect 1207 17741 1209 17793
rect 274 17740 1209 17741
rect 1154 17734 1209 17740
rect 1754 17796 1814 17802
rect 2267 17796 2325 17805
rect 1754 17793 2325 17796
rect 2838 17793 2898 17798
rect 1754 17792 2898 17793
rect 1754 17740 1758 17792
rect 1810 17790 2908 17792
rect 1810 17740 2270 17790
rect 1754 17738 2270 17740
rect 2322 17788 2908 17790
rect 2322 17738 2842 17788
rect 1754 17736 2842 17738
rect 2894 17736 2908 17788
rect 1754 17730 1814 17736
rect 2267 17735 2908 17736
rect 2267 17723 2325 17735
rect 2838 17732 2908 17735
rect 3262 17734 3268 17786
rect 3320 17734 3326 17786
rect 3976 17804 4028 17810
rect 3561 17755 3613 17761
rect 3975 17755 3976 17798
rect 2838 17726 2898 17732
rect 2768 17692 2816 17696
rect 378 17681 433 17687
rect 1248 17682 1300 17688
rect 433 17678 619 17681
rect 433 17634 1248 17678
rect 433 17626 619 17634
rect 2020 17682 2072 17688
rect 2522 17684 2574 17686
rect 1300 17634 2020 17678
rect 378 17620 433 17626
rect 1248 17624 1300 17630
rect 2020 17624 2072 17630
rect 2509 17682 2587 17684
rect 2509 17626 2520 17682
rect 2576 17626 2587 17682
rect 2760 17640 2766 17692
rect 2818 17688 2824 17692
rect 3270 17688 3314 17734
rect 3564 17716 3605 17755
rect 4622 17763 4628 17815
rect 4680 17763 4686 17815
rect 3976 17746 4028 17752
rect 2818 17644 3314 17688
rect 3979 17699 4018 17746
rect 4637 17699 4671 17763
rect 5122 17716 5164 18529
rect 5202 17819 5244 18864
rect 5197 17813 5249 17819
rect 5197 17755 5249 17761
rect 5202 17716 5244 17755
rect 5282 17716 5324 18864
rect 5362 17716 5404 18864
rect 5442 17716 5484 18864
rect 5522 17716 5564 18864
rect 6820 18860 6872 18866
rect 6974 18862 7026 18868
rect 5662 18738 6202 18780
rect 5662 18682 5704 18738
rect 5760 18736 5784 18738
rect 5840 18736 5864 18738
rect 5920 18736 5944 18738
rect 6000 18736 6024 18738
rect 6080 18736 6104 18738
rect 5766 18684 5778 18736
rect 5840 18684 5842 18736
rect 6022 18684 6024 18736
rect 6086 18684 6098 18736
rect 5760 18682 5784 18684
rect 5840 18682 5864 18684
rect 5920 18682 5944 18684
rect 6000 18682 6024 18684
rect 6080 18682 6104 18684
rect 6160 18682 6202 18738
rect 6504 18736 6510 18788
rect 6562 18736 6568 18788
rect 5662 18640 6202 18682
rect 6518 18572 6556 18736
rect 6523 18502 6553 18572
rect 6506 18450 6512 18502
rect 6564 18450 6570 18502
rect 6843 18298 6895 18304
rect 6895 18253 7241 18292
rect 5682 18200 6222 18242
rect 6843 18240 6895 18246
rect 5682 18144 5724 18200
rect 5780 18198 5804 18200
rect 5860 18198 5884 18200
rect 5940 18198 5964 18200
rect 6020 18198 6044 18200
rect 6100 18198 6124 18200
rect 5786 18146 5798 18198
rect 5860 18146 5862 18198
rect 6042 18146 6044 18198
rect 6106 18146 6118 18198
rect 5780 18144 5804 18146
rect 5860 18144 5884 18146
rect 5940 18144 5964 18146
rect 6020 18144 6044 18146
rect 6100 18144 6124 18146
rect 6180 18144 6222 18200
rect 5682 18102 6222 18144
rect 6250 17974 6304 17980
rect 6974 17974 7026 17976
rect 6250 17972 7042 17974
rect 6302 17970 7042 17972
rect 6302 17920 6974 17970
rect 6250 17918 6974 17920
rect 7026 17918 7042 17970
rect 6250 17912 6304 17918
rect 6974 17912 7026 17918
rect 5934 17804 5986 17810
rect 6580 17764 6586 17816
rect 6638 17764 6644 17816
rect 5934 17746 5986 17752
rect 3979 17660 4673 17699
rect 4862 17690 4914 17696
rect 2818 17640 2824 17644
rect 2509 17624 2587 17626
rect 2522 17622 2574 17624
rect 2768 17600 2812 17640
rect 5015 17692 5067 17698
rect 4914 17650 5015 17679
rect 144 16294 212 17446
rect 274 17373 329 17562
rect 372 17526 378 17582
rect 434 17526 440 17582
rect 274 17367 332 17373
rect 274 17313 278 17367
rect 277 17192 332 17313
rect 378 17354 434 17526
rect 1324 17499 1960 17552
rect 1324 17497 1374 17499
rect 1430 17497 1454 17499
rect 1510 17497 1534 17499
rect 1590 17497 1614 17499
rect 1670 17497 1694 17499
rect 1750 17497 1774 17499
rect 1830 17497 1854 17499
rect 1910 17497 1960 17499
rect 1324 17445 1360 17497
rect 1604 17445 1614 17497
rect 1670 17445 1680 17497
rect 1924 17445 1960 17497
rect 1324 17443 1374 17445
rect 1430 17443 1454 17445
rect 1510 17443 1534 17445
rect 1590 17443 1614 17445
rect 1670 17443 1694 17445
rect 1750 17443 1774 17445
rect 1830 17443 1854 17445
rect 1910 17443 1960 17445
rect 1324 17412 1960 17443
rect 3564 17365 3605 17636
rect 4862 17632 4914 17638
rect 5015 17634 5067 17640
rect 5122 17636 5163 17716
rect 5282 17636 5323 17716
rect 5362 17636 5403 17716
rect 5442 17636 5483 17716
rect 5522 17636 5563 17716
rect 5938 17700 5976 17746
rect 6596 17700 6630 17764
rect 5938 17660 6632 17700
rect 6820 17690 6872 17696
rect 6974 17692 7026 17698
rect 6872 17650 6974 17680
rect 3704 17510 4244 17552
rect 3704 17454 3746 17510
rect 3802 17508 3826 17510
rect 3882 17508 3906 17510
rect 3962 17508 3986 17510
rect 4042 17508 4066 17510
rect 4122 17508 4146 17510
rect 3808 17456 3820 17508
rect 3882 17456 3884 17508
rect 4064 17456 4066 17508
rect 4128 17456 4140 17508
rect 3802 17454 3826 17456
rect 3882 17454 3906 17456
rect 3962 17454 3986 17456
rect 4042 17454 4066 17456
rect 4122 17454 4146 17456
rect 4202 17454 4244 17510
rect 4546 17507 4552 17559
rect 4604 17507 4610 17559
rect 3704 17412 4244 17454
rect 3564 17359 3617 17365
rect 274 16567 329 17192
rect 378 16738 433 17354
rect 3564 17307 3565 17359
rect 4559 17343 4598 17507
rect 3564 17301 3617 17307
rect 1348 16973 1880 17014
rect 1348 16917 1388 16973
rect 1444 16971 1468 16973
rect 1524 16971 1548 16973
rect 1604 16971 1628 16973
rect 1684 16971 1708 16973
rect 1764 16971 1788 16973
rect 1450 16919 1462 16971
rect 1524 16919 1526 16971
rect 1706 16919 1708 16971
rect 1770 16919 1782 16971
rect 1444 16917 1468 16919
rect 1524 16917 1548 16919
rect 1604 16917 1628 16919
rect 1684 16917 1708 16919
rect 1764 16917 1788 16919
rect 1844 16917 1880 16973
rect 560 16900 612 16906
rect 700 16898 756 16904
rect 612 16896 976 16898
rect 612 16848 702 16896
rect 560 16844 702 16848
rect 754 16844 976 16896
rect 1348 16874 1880 16917
rect 2759 16856 2827 16864
rect 560 16842 1268 16844
rect 700 16836 756 16842
rect 920 16836 1268 16842
rect 2759 16836 2769 16856
rect 920 16804 2769 16836
rect 2821 16804 2827 16856
rect 920 16792 2827 16804
rect 920 16788 1268 16792
rect 852 16746 904 16752
rect 372 16683 378 16738
rect 433 16683 439 16738
rect 1396 16747 2851 16756
rect 3268 16751 3320 16757
rect 1396 16742 3268 16747
rect 904 16712 3268 16742
rect 904 16698 1440 16712
rect 2851 16703 3268 16712
rect 852 16688 904 16694
rect 3268 16693 3320 16699
rect 1930 16666 1990 16677
rect 1004 16654 1056 16660
rect 1930 16655 1932 16666
rect 1056 16643 1242 16650
rect 1599 16643 1932 16655
rect 1056 16621 1932 16643
rect 1056 16609 1633 16621
rect 1930 16610 1932 16621
rect 1988 16655 1990 16666
rect 1988 16621 1991 16655
rect 1988 16610 1990 16621
rect 1056 16606 1242 16609
rect 1004 16596 1056 16602
rect 1930 16599 1990 16610
rect 3564 16591 3605 17301
rect 5023 17100 5029 17152
rect 5081 17100 5087 17152
rect 4744 17070 4796 17076
rect 5036 17064 5075 17100
rect 4796 17025 5075 17064
rect 3724 16972 4264 17014
rect 4744 17012 4796 17018
rect 3724 16916 3766 16972
rect 3822 16970 3846 16972
rect 3902 16970 3926 16972
rect 3982 16970 4006 16972
rect 4062 16970 4086 16972
rect 4142 16970 4166 16972
rect 3828 16918 3840 16970
rect 3902 16918 3904 16970
rect 4084 16918 4086 16970
rect 4148 16918 4160 16970
rect 3822 16916 3846 16918
rect 3902 16916 3926 16918
rect 3982 16916 4006 16918
rect 4062 16916 4086 16918
rect 4142 16916 4166 16918
rect 4222 16916 4264 16972
rect 3724 16874 4264 16916
rect 4291 16745 4346 16751
rect 5016 16745 5068 16748
rect 4291 16743 5084 16745
rect 4291 16691 4292 16743
rect 4344 16742 5084 16743
rect 4344 16691 5016 16742
rect 4291 16690 5016 16691
rect 5068 16690 5084 16742
rect 4291 16684 4346 16690
rect 5016 16684 5068 16690
rect 5122 16591 5164 17636
rect 5202 17365 5244 17636
rect 5197 17359 5249 17365
rect 5197 17301 5249 17307
rect 3561 16585 3613 16591
rect 1154 16567 1209 16573
rect 274 16565 1209 16567
rect 274 16513 1155 16565
rect 1207 16513 1209 16565
rect 274 16512 1209 16513
rect 1154 16506 1209 16512
rect 1754 16568 1814 16574
rect 2267 16568 2325 16577
rect 1754 16565 2325 16568
rect 2838 16565 2898 16570
rect 1754 16564 2898 16565
rect 1754 16512 1758 16564
rect 1810 16562 2908 16564
rect 1810 16512 2270 16562
rect 1754 16510 2270 16512
rect 2322 16560 2908 16562
rect 2322 16510 2842 16560
rect 1754 16508 2842 16510
rect 2894 16508 2908 16560
rect 1754 16502 1814 16508
rect 2267 16507 2908 16508
rect 2267 16495 2325 16507
rect 2838 16504 2908 16507
rect 3262 16506 3268 16558
rect 3320 16506 3326 16558
rect 3976 16576 4028 16582
rect 3561 16527 3613 16533
rect 3975 16527 3976 16570
rect 2838 16498 2898 16504
rect 2768 16464 2816 16468
rect 378 16453 433 16459
rect 1248 16454 1300 16460
rect 433 16450 619 16453
rect 433 16406 1248 16450
rect 433 16398 619 16406
rect 2020 16454 2072 16460
rect 2522 16456 2574 16458
rect 1300 16406 2020 16450
rect 378 16392 433 16398
rect 1248 16396 1300 16402
rect 2020 16396 2072 16402
rect 2509 16454 2587 16456
rect 2509 16398 2520 16454
rect 2576 16398 2587 16454
rect 2760 16412 2766 16464
rect 2818 16460 2824 16464
rect 3270 16460 3314 16506
rect 3564 16488 3605 16527
rect 4622 16535 4628 16587
rect 4680 16535 4686 16587
rect 5117 16585 5169 16591
rect 3976 16518 4028 16524
rect 2818 16416 3314 16460
rect 3979 16471 4018 16518
rect 4637 16471 4671 16535
rect 5117 16527 5169 16533
rect 5122 16488 5164 16527
rect 5202 16488 5244 17301
rect 5282 16488 5324 17636
rect 5362 16488 5404 17636
rect 5442 16488 5484 17636
rect 5522 16488 5564 17636
rect 6820 17632 6872 17638
rect 6974 17634 7026 17640
rect 5662 17510 6202 17552
rect 5662 17454 5704 17510
rect 5760 17508 5784 17510
rect 5840 17508 5864 17510
rect 5920 17508 5944 17510
rect 6000 17508 6024 17510
rect 6080 17508 6104 17510
rect 5766 17456 5778 17508
rect 5840 17456 5842 17508
rect 6022 17456 6024 17508
rect 6086 17456 6098 17508
rect 5760 17454 5784 17456
rect 5840 17454 5864 17456
rect 5920 17454 5944 17456
rect 6000 17454 6024 17456
rect 6080 17454 6104 17456
rect 6160 17454 6202 17510
rect 6504 17508 6510 17560
rect 6562 17508 6568 17560
rect 5662 17412 6202 17454
rect 6518 17344 6556 17508
rect 7101 17220 7107 17272
rect 7159 17220 7165 17272
rect 6868 17070 6920 17076
rect 7119 17064 7147 17220
rect 6920 17025 7147 17064
rect 5682 16972 6222 17014
rect 6868 17012 6920 17018
rect 5682 16916 5724 16972
rect 5780 16970 5804 16972
rect 5860 16970 5884 16972
rect 5940 16970 5964 16972
rect 6020 16970 6044 16972
rect 6100 16970 6124 16972
rect 5786 16918 5798 16970
rect 5860 16918 5862 16970
rect 6042 16918 6044 16970
rect 6106 16918 6118 16970
rect 5780 16916 5804 16918
rect 5860 16916 5884 16918
rect 5940 16916 5964 16918
rect 6020 16916 6044 16918
rect 6100 16916 6124 16918
rect 6180 16916 6222 16972
rect 5682 16874 6222 16916
rect 6250 16746 6304 16752
rect 6974 16746 7026 16748
rect 6250 16744 7042 16746
rect 6302 16742 7042 16744
rect 6302 16692 6974 16742
rect 6250 16690 6974 16692
rect 7026 16690 7042 16742
rect 6250 16684 6304 16690
rect 6974 16684 7026 16690
rect 5934 16576 5986 16582
rect 6580 16536 6586 16588
rect 6638 16536 6644 16588
rect 5934 16518 5986 16524
rect 3979 16432 4673 16471
rect 4862 16462 4914 16468
rect 2818 16412 2824 16416
rect 2509 16396 2587 16398
rect 2522 16394 2574 16396
rect 2768 16372 2812 16412
rect 5015 16464 5067 16470
rect 4914 16422 5015 16451
rect 144 15058 212 16226
rect 274 16145 329 16334
rect 372 16298 378 16354
rect 434 16298 440 16354
rect 274 16139 332 16145
rect 274 16085 278 16139
rect 277 15964 332 16085
rect 378 16126 434 16298
rect 1324 16271 1960 16324
rect 1324 16269 1374 16271
rect 1430 16269 1454 16271
rect 1510 16269 1534 16271
rect 1590 16269 1614 16271
rect 1670 16269 1694 16271
rect 1750 16269 1774 16271
rect 1830 16269 1854 16271
rect 1910 16269 1960 16271
rect 1324 16217 1360 16269
rect 1604 16217 1614 16269
rect 1670 16217 1680 16269
rect 1924 16217 1960 16269
rect 1324 16215 1374 16217
rect 1430 16215 1454 16217
rect 1510 16215 1534 16217
rect 1590 16215 1614 16217
rect 1670 16215 1694 16217
rect 1750 16215 1774 16217
rect 1830 16215 1854 16217
rect 1910 16215 1960 16217
rect 1324 16184 1960 16215
rect 3564 16137 3605 16408
rect 4862 16404 4914 16410
rect 5015 16406 5067 16412
rect 5202 16408 5243 16488
rect 5282 16408 5323 16488
rect 5362 16408 5403 16488
rect 5442 16408 5483 16488
rect 5522 16408 5563 16488
rect 5938 16472 5976 16518
rect 6596 16472 6630 16536
rect 5938 16432 6632 16472
rect 6820 16462 6872 16468
rect 6974 16464 7026 16470
rect 6872 16422 6974 16452
rect 3704 16282 4244 16324
rect 3704 16226 3746 16282
rect 3802 16280 3826 16282
rect 3882 16280 3906 16282
rect 3962 16280 3986 16282
rect 4042 16280 4066 16282
rect 4122 16280 4146 16282
rect 3808 16228 3820 16280
rect 3882 16228 3884 16280
rect 4064 16228 4066 16280
rect 4128 16228 4140 16280
rect 3802 16226 3826 16228
rect 3882 16226 3906 16228
rect 3962 16226 3986 16228
rect 4042 16226 4066 16228
rect 4122 16226 4146 16228
rect 4202 16226 4244 16282
rect 4546 16279 4552 16331
rect 4604 16279 4610 16331
rect 3704 16184 4244 16226
rect 3564 16131 3617 16137
rect 274 15339 329 15964
rect 378 15510 433 16126
rect 3564 16079 3565 16131
rect 4559 16115 4598 16279
rect 5122 16137 5164 16408
rect 5117 16131 5169 16137
rect 3564 16073 3617 16079
rect 5117 16073 5169 16079
rect 1348 15745 1880 15786
rect 1348 15689 1388 15745
rect 1444 15743 1468 15745
rect 1524 15743 1548 15745
rect 1604 15743 1628 15745
rect 1684 15743 1708 15745
rect 1764 15743 1788 15745
rect 1450 15691 1462 15743
rect 1524 15691 1526 15743
rect 1706 15691 1708 15743
rect 1770 15691 1782 15743
rect 1444 15689 1468 15691
rect 1524 15689 1548 15691
rect 1604 15689 1628 15691
rect 1684 15689 1708 15691
rect 1764 15689 1788 15691
rect 1844 15689 1880 15745
rect 560 15672 612 15678
rect 700 15670 756 15676
rect 612 15668 976 15670
rect 612 15620 702 15668
rect 560 15616 702 15620
rect 754 15616 976 15668
rect 1348 15646 1880 15689
rect 2759 15628 2827 15636
rect 560 15614 1268 15616
rect 700 15608 756 15614
rect 920 15608 1268 15614
rect 2759 15608 2769 15628
rect 920 15576 2769 15608
rect 2821 15576 2827 15628
rect 920 15564 2827 15576
rect 920 15560 1268 15564
rect 852 15518 904 15524
rect 372 15455 378 15510
rect 433 15455 439 15510
rect 1396 15519 2851 15528
rect 3268 15523 3320 15529
rect 1396 15514 3268 15519
rect 904 15484 3268 15514
rect 904 15470 1440 15484
rect 2851 15475 3268 15484
rect 852 15460 904 15466
rect 3268 15465 3320 15471
rect 1930 15438 1990 15449
rect 1004 15426 1056 15432
rect 1930 15427 1932 15438
rect 1056 15415 1242 15422
rect 1599 15415 1932 15427
rect 1056 15393 1932 15415
rect 1056 15381 1633 15393
rect 1930 15382 1932 15393
rect 1988 15427 1990 15438
rect 1988 15393 1991 15427
rect 1988 15382 1990 15393
rect 1056 15378 1242 15381
rect 1004 15368 1056 15374
rect 1930 15371 1990 15382
rect 3564 15363 3605 16073
rect 5029 15909 5035 15961
rect 5087 15909 5093 15961
rect 4744 15842 4796 15848
rect 5047 15836 5075 15909
rect 4796 15797 5075 15836
rect 3724 15744 4264 15786
rect 4744 15784 4796 15790
rect 3724 15688 3766 15744
rect 3822 15742 3846 15744
rect 3902 15742 3926 15744
rect 3982 15742 4006 15744
rect 4062 15742 4086 15744
rect 4142 15742 4166 15744
rect 3828 15690 3840 15742
rect 3902 15690 3904 15742
rect 4084 15690 4086 15742
rect 4148 15690 4160 15742
rect 3822 15688 3846 15690
rect 3902 15688 3926 15690
rect 3982 15688 4006 15690
rect 4062 15688 4086 15690
rect 4142 15688 4166 15690
rect 4222 15688 4264 15744
rect 3724 15646 4264 15688
rect 4291 15517 4346 15523
rect 5016 15517 5068 15520
rect 4291 15515 5084 15517
rect 4291 15463 4292 15515
rect 4344 15514 5084 15515
rect 4344 15463 5016 15514
rect 4291 15462 5016 15463
rect 5068 15462 5084 15514
rect 4291 15456 4346 15462
rect 5016 15456 5068 15462
rect 3561 15357 3613 15363
rect 1154 15339 1209 15345
rect 274 15337 1209 15339
rect 274 15285 1155 15337
rect 1207 15285 1209 15337
rect 274 15284 1209 15285
rect 1154 15278 1209 15284
rect 1754 15340 1814 15346
rect 2267 15340 2325 15349
rect 1754 15337 2325 15340
rect 2838 15337 2898 15342
rect 1754 15336 2898 15337
rect 1754 15284 1758 15336
rect 1810 15334 2908 15336
rect 1810 15284 2270 15334
rect 1754 15282 2270 15284
rect 2322 15332 2908 15334
rect 2322 15282 2842 15332
rect 1754 15280 2842 15282
rect 2894 15280 2908 15332
rect 1754 15274 1814 15280
rect 2267 15279 2908 15280
rect 2267 15267 2325 15279
rect 2838 15276 2908 15279
rect 3262 15278 3268 15330
rect 3320 15278 3326 15330
rect 3976 15348 4028 15354
rect 3561 15299 3613 15305
rect 3975 15299 3976 15342
rect 2838 15270 2898 15276
rect 2768 15236 2816 15240
rect 378 15225 433 15231
rect 1248 15226 1300 15232
rect 433 15222 619 15225
rect 433 15178 1248 15222
rect 433 15170 619 15178
rect 2020 15226 2072 15232
rect 2522 15228 2574 15230
rect 1300 15178 2020 15222
rect 378 15164 433 15170
rect 1248 15168 1300 15174
rect 2020 15168 2072 15174
rect 2509 15226 2587 15228
rect 2509 15170 2520 15226
rect 2576 15170 2587 15226
rect 2760 15184 2766 15236
rect 2818 15232 2824 15236
rect 3270 15232 3314 15278
rect 3564 15260 3605 15299
rect 4622 15307 4628 15359
rect 4680 15307 4686 15359
rect 3976 15290 4028 15296
rect 2818 15188 3314 15232
rect 3979 15243 4018 15290
rect 4637 15243 4671 15307
rect 5122 15260 5164 16073
rect 5202 15260 5244 16408
rect 5282 15363 5324 16408
rect 5279 15357 5331 15363
rect 5279 15299 5331 15305
rect 5282 15260 5324 15299
rect 5362 15260 5404 16408
rect 5442 15260 5484 16408
rect 5522 15260 5564 16408
rect 6820 16404 6872 16410
rect 6974 16406 7026 16412
rect 5662 16282 6202 16324
rect 5662 16226 5704 16282
rect 5760 16280 5784 16282
rect 5840 16280 5864 16282
rect 5920 16280 5944 16282
rect 6000 16280 6024 16282
rect 6080 16280 6104 16282
rect 5766 16228 5778 16280
rect 5840 16228 5842 16280
rect 6022 16228 6024 16280
rect 6086 16228 6098 16280
rect 5760 16226 5784 16228
rect 5840 16226 5864 16228
rect 5920 16226 5944 16228
rect 6000 16226 6024 16228
rect 6080 16226 6104 16228
rect 6160 16226 6202 16282
rect 6504 16280 6510 16332
rect 6562 16280 6568 16332
rect 5662 16184 6202 16226
rect 6518 16116 6556 16280
rect 6974 15962 7026 15968
rect 7202 15951 7241 18253
rect 7026 15921 7241 15951
rect 6974 15904 7026 15910
rect 5682 15744 6222 15786
rect 5682 15688 5724 15744
rect 5780 15742 5804 15744
rect 5860 15742 5884 15744
rect 5940 15742 5964 15744
rect 6020 15742 6044 15744
rect 6100 15742 6124 15744
rect 5786 15690 5798 15742
rect 5860 15690 5862 15742
rect 6042 15690 6044 15742
rect 6106 15690 6118 15742
rect 5780 15688 5804 15690
rect 5860 15688 5884 15690
rect 5940 15688 5964 15690
rect 6020 15688 6044 15690
rect 6100 15688 6124 15690
rect 6180 15688 6222 15744
rect 5682 15646 6222 15688
rect 6250 15518 6304 15524
rect 6974 15518 7026 15520
rect 6250 15516 7042 15518
rect 6302 15514 7042 15516
rect 6302 15464 6974 15514
rect 6250 15462 6974 15464
rect 7026 15462 7042 15514
rect 6250 15456 6304 15462
rect 6974 15456 7026 15462
rect 5934 15348 5986 15354
rect 6580 15308 6586 15360
rect 6638 15308 6644 15360
rect 5934 15290 5986 15296
rect 3979 15204 4673 15243
rect 4862 15234 4914 15240
rect 2818 15184 2824 15188
rect 2509 15168 2587 15170
rect 2522 15166 2574 15168
rect 2768 15144 2812 15184
rect 5015 15236 5067 15242
rect 4914 15194 5015 15223
rect 144 13838 212 14990
rect 274 14917 329 15106
rect 372 15070 378 15126
rect 434 15070 440 15126
rect 274 14911 332 14917
rect 274 14857 278 14911
rect 277 14736 332 14857
rect 378 14898 434 15070
rect 1324 15043 1960 15096
rect 1324 15041 1374 15043
rect 1430 15041 1454 15043
rect 1510 15041 1534 15043
rect 1590 15041 1614 15043
rect 1670 15041 1694 15043
rect 1750 15041 1774 15043
rect 1830 15041 1854 15043
rect 1910 15041 1960 15043
rect 1324 14989 1360 15041
rect 1604 14989 1614 15041
rect 1670 14989 1680 15041
rect 1924 14989 1960 15041
rect 1324 14987 1374 14989
rect 1430 14987 1454 14989
rect 1510 14987 1534 14989
rect 1590 14987 1614 14989
rect 1670 14987 1694 14989
rect 1750 14987 1774 14989
rect 1830 14987 1854 14989
rect 1910 14987 1960 14989
rect 1324 14956 1960 14987
rect 3564 14909 3605 15180
rect 4862 15176 4914 15182
rect 5015 15178 5067 15184
rect 5122 15180 5163 15260
rect 5202 15180 5243 15260
rect 5362 15180 5403 15260
rect 5442 15180 5483 15260
rect 5522 15180 5563 15260
rect 5938 15244 5976 15290
rect 6596 15244 6630 15308
rect 5938 15204 6632 15244
rect 6820 15234 6872 15240
rect 6974 15236 7026 15242
rect 6872 15194 6974 15224
rect 3704 15054 4244 15096
rect 3704 14998 3746 15054
rect 3802 15052 3826 15054
rect 3882 15052 3906 15054
rect 3962 15052 3986 15054
rect 4042 15052 4066 15054
rect 4122 15052 4146 15054
rect 3808 15000 3820 15052
rect 3882 15000 3884 15052
rect 4064 15000 4066 15052
rect 4128 15000 4140 15052
rect 3802 14998 3826 15000
rect 3882 14998 3906 15000
rect 3962 14998 3986 15000
rect 4042 14998 4066 15000
rect 4122 14998 4146 15000
rect 4202 14998 4244 15054
rect 4546 15051 4552 15103
rect 4604 15051 4610 15103
rect 3704 14956 4244 14998
rect 3564 14903 3617 14909
rect 274 14111 329 14736
rect 378 14282 433 14898
rect 3564 14851 3565 14903
rect 4559 14887 4598 15051
rect 3564 14845 3617 14851
rect 1348 14517 1880 14558
rect 1348 14461 1388 14517
rect 1444 14515 1468 14517
rect 1524 14515 1548 14517
rect 1604 14515 1628 14517
rect 1684 14515 1708 14517
rect 1764 14515 1788 14517
rect 1450 14463 1462 14515
rect 1524 14463 1526 14515
rect 1706 14463 1708 14515
rect 1770 14463 1782 14515
rect 1444 14461 1468 14463
rect 1524 14461 1548 14463
rect 1604 14461 1628 14463
rect 1684 14461 1708 14463
rect 1764 14461 1788 14463
rect 1844 14461 1880 14517
rect 560 14444 612 14450
rect 700 14442 756 14448
rect 612 14440 976 14442
rect 612 14392 702 14440
rect 560 14388 702 14392
rect 754 14388 976 14440
rect 1348 14418 1880 14461
rect 2759 14400 2827 14408
rect 560 14386 1268 14388
rect 700 14380 756 14386
rect 920 14380 1268 14386
rect 2759 14380 2769 14400
rect 920 14348 2769 14380
rect 2821 14348 2827 14400
rect 920 14336 2827 14348
rect 920 14332 1268 14336
rect 852 14290 904 14296
rect 372 14227 378 14282
rect 433 14227 439 14282
rect 1396 14291 2851 14300
rect 3268 14295 3320 14301
rect 1396 14286 3268 14291
rect 904 14256 3268 14286
rect 904 14242 1440 14256
rect 2851 14247 3268 14256
rect 852 14232 904 14238
rect 3268 14237 3320 14243
rect 1930 14210 1990 14221
rect 1004 14198 1056 14204
rect 1930 14199 1932 14210
rect 1056 14187 1242 14194
rect 1599 14187 1932 14199
rect 1056 14165 1932 14187
rect 1056 14153 1633 14165
rect 1930 14154 1932 14165
rect 1988 14199 1990 14210
rect 1988 14165 1991 14199
rect 1988 14154 1990 14165
rect 1056 14150 1242 14153
rect 1004 14140 1056 14146
rect 1930 14143 1990 14154
rect 3564 14135 3605 14845
rect 5023 14644 5029 14696
rect 5081 14644 5087 14696
rect 4744 14614 4796 14620
rect 5036 14608 5075 14644
rect 4796 14569 5075 14608
rect 3724 14516 4264 14558
rect 4744 14556 4796 14562
rect 3724 14460 3766 14516
rect 3822 14514 3846 14516
rect 3902 14514 3926 14516
rect 3982 14514 4006 14516
rect 4062 14514 4086 14516
rect 4142 14514 4166 14516
rect 3828 14462 3840 14514
rect 3902 14462 3904 14514
rect 4084 14462 4086 14514
rect 4148 14462 4160 14514
rect 3822 14460 3846 14462
rect 3902 14460 3926 14462
rect 3982 14460 4006 14462
rect 4062 14460 4086 14462
rect 4142 14460 4166 14462
rect 4222 14460 4264 14516
rect 3724 14418 4264 14460
rect 4291 14289 4346 14295
rect 5016 14289 5068 14292
rect 4291 14287 5084 14289
rect 4291 14235 4292 14287
rect 4344 14286 5084 14287
rect 4344 14235 5016 14286
rect 4291 14234 5016 14235
rect 5068 14234 5084 14286
rect 4291 14228 4346 14234
rect 5016 14228 5068 14234
rect 5122 14135 5164 15180
rect 3561 14129 3613 14135
rect 1154 14111 1209 14117
rect 274 14109 1209 14111
rect 274 14057 1155 14109
rect 1207 14057 1209 14109
rect 274 14056 1209 14057
rect 1154 14050 1209 14056
rect 1754 14112 1814 14118
rect 2267 14112 2325 14121
rect 1754 14109 2325 14112
rect 2838 14109 2898 14114
rect 1754 14108 2898 14109
rect 1754 14056 1758 14108
rect 1810 14106 2908 14108
rect 1810 14056 2270 14106
rect 1754 14054 2270 14056
rect 2322 14104 2908 14106
rect 2322 14054 2842 14104
rect 1754 14052 2842 14054
rect 2894 14052 2908 14104
rect 1754 14046 1814 14052
rect 2267 14051 2908 14052
rect 2267 14039 2325 14051
rect 2838 14048 2908 14051
rect 3262 14050 3268 14102
rect 3320 14050 3326 14102
rect 3976 14120 4028 14126
rect 3561 14071 3613 14077
rect 3975 14071 3976 14114
rect 2838 14042 2898 14048
rect 2768 14008 2816 14012
rect 378 13997 433 14003
rect 1248 13998 1300 14004
rect 433 13994 619 13997
rect 433 13950 1248 13994
rect 433 13942 619 13950
rect 2020 13998 2072 14004
rect 2522 14000 2574 14002
rect 1300 13950 2020 13994
rect 378 13936 433 13942
rect 1248 13940 1300 13946
rect 2020 13940 2072 13946
rect 2509 13998 2587 14000
rect 2509 13942 2520 13998
rect 2576 13942 2587 13998
rect 2760 13956 2766 14008
rect 2818 14004 2824 14008
rect 3270 14004 3314 14050
rect 3564 14032 3605 14071
rect 4622 14079 4628 14131
rect 4680 14079 4686 14131
rect 5117 14129 5169 14135
rect 3976 14062 4028 14068
rect 2818 13960 3314 14004
rect 3979 14015 4018 14062
rect 4637 14015 4671 14079
rect 5117 14071 5169 14077
rect 5122 14032 5164 14071
rect 5202 14032 5244 15180
rect 5282 14909 5324 15180
rect 5279 14903 5331 14909
rect 5279 14845 5331 14851
rect 5282 14032 5324 14845
rect 5362 14032 5404 15180
rect 5442 14032 5484 15180
rect 5522 14032 5564 15180
rect 6820 15176 6872 15182
rect 6974 15178 7026 15184
rect 5662 15054 6202 15096
rect 5662 14998 5704 15054
rect 5760 15052 5784 15054
rect 5840 15052 5864 15054
rect 5920 15052 5944 15054
rect 6000 15052 6024 15054
rect 6080 15052 6104 15054
rect 5766 15000 5778 15052
rect 5840 15000 5842 15052
rect 6022 15000 6024 15052
rect 6086 15000 6098 15052
rect 5760 14998 5784 15000
rect 5840 14998 5864 15000
rect 5920 14998 5944 15000
rect 6000 14998 6024 15000
rect 6080 14998 6104 15000
rect 6160 14998 6202 15054
rect 6504 15052 6510 15104
rect 6562 15052 6568 15104
rect 5662 14956 6202 14998
rect 6518 14926 6556 15052
rect 6517 14887 7337 14926
rect 6868 14614 6920 14620
rect 6920 14569 7147 14608
rect 5682 14516 6222 14558
rect 6868 14556 6920 14562
rect 5682 14460 5724 14516
rect 5780 14514 5804 14516
rect 5860 14514 5884 14516
rect 5940 14514 5964 14516
rect 6020 14514 6044 14516
rect 6100 14514 6124 14516
rect 5786 14462 5798 14514
rect 5860 14462 5862 14514
rect 6042 14462 6044 14514
rect 6106 14462 6118 14514
rect 5780 14460 5804 14462
rect 5860 14460 5884 14462
rect 5940 14460 5964 14462
rect 6020 14460 6044 14462
rect 6100 14460 6124 14462
rect 6180 14460 6222 14516
rect 5682 14418 6222 14460
rect 7188 14444 7194 14496
rect 7246 14444 7252 14496
rect 6250 14290 6304 14296
rect 6974 14290 7026 14292
rect 6250 14288 7042 14290
rect 6302 14286 7042 14288
rect 6302 14236 6974 14286
rect 6250 14234 6974 14236
rect 7026 14234 7042 14286
rect 6250 14228 6304 14234
rect 6974 14228 7026 14234
rect 5934 14120 5986 14126
rect 6580 14080 6586 14132
rect 6638 14080 6644 14132
rect 5934 14062 5986 14068
rect 3979 13976 4673 14015
rect 4862 14006 4914 14012
rect 2818 13956 2824 13960
rect 2509 13940 2587 13942
rect 2522 13938 2574 13940
rect 2768 13916 2812 13956
rect 5015 14008 5067 14014
rect 4914 13966 5015 13995
rect 144 12602 212 13770
rect 274 13689 329 13878
rect 372 13842 378 13898
rect 434 13842 440 13898
rect 274 13683 332 13689
rect 274 13629 278 13683
rect 277 13508 332 13629
rect 378 13670 434 13842
rect 1324 13815 1960 13868
rect 1324 13813 1374 13815
rect 1430 13813 1454 13815
rect 1510 13813 1534 13815
rect 1590 13813 1614 13815
rect 1670 13813 1694 13815
rect 1750 13813 1774 13815
rect 1830 13813 1854 13815
rect 1910 13813 1960 13815
rect 1324 13761 1360 13813
rect 1604 13761 1614 13813
rect 1670 13761 1680 13813
rect 1924 13761 1960 13813
rect 1324 13759 1374 13761
rect 1430 13759 1454 13761
rect 1510 13759 1534 13761
rect 1590 13759 1614 13761
rect 1670 13759 1694 13761
rect 1750 13759 1774 13761
rect 1830 13759 1854 13761
rect 1910 13759 1960 13761
rect 1324 13728 1960 13759
rect 3564 13681 3605 13952
rect 4862 13948 4914 13954
rect 5015 13950 5067 13956
rect 5202 13952 5243 14032
rect 5282 13952 5323 14032
rect 5362 13952 5403 14032
rect 5442 13952 5483 14032
rect 5522 13952 5563 14032
rect 5938 14016 5976 14062
rect 6596 14016 6630 14080
rect 5938 13976 6632 14016
rect 6820 14006 6872 14012
rect 6974 14008 7026 14014
rect 6872 13966 6974 13996
rect 3704 13826 4244 13868
rect 3704 13770 3746 13826
rect 3802 13824 3826 13826
rect 3882 13824 3906 13826
rect 3962 13824 3986 13826
rect 4042 13824 4066 13826
rect 4122 13824 4146 13826
rect 3808 13772 3820 13824
rect 3882 13772 3884 13824
rect 4064 13772 4066 13824
rect 4128 13772 4140 13824
rect 3802 13770 3826 13772
rect 3882 13770 3906 13772
rect 3962 13770 3986 13772
rect 4042 13770 4066 13772
rect 4122 13770 4146 13772
rect 4202 13770 4244 13826
rect 4546 13823 4552 13875
rect 4604 13823 4610 13875
rect 3704 13728 4244 13770
rect 3564 13675 3617 13681
rect 274 12883 329 13508
rect 378 13054 433 13670
rect 3564 13623 3565 13675
rect 4559 13659 4598 13823
rect 5122 13681 5164 13952
rect 5117 13675 5169 13681
rect 3564 13617 3617 13623
rect 5117 13617 5169 13623
rect 1348 13289 1880 13330
rect 1348 13233 1388 13289
rect 1444 13287 1468 13289
rect 1524 13287 1548 13289
rect 1604 13287 1628 13289
rect 1684 13287 1708 13289
rect 1764 13287 1788 13289
rect 1450 13235 1462 13287
rect 1524 13235 1526 13287
rect 1706 13235 1708 13287
rect 1770 13235 1782 13287
rect 1444 13233 1468 13235
rect 1524 13233 1548 13235
rect 1604 13233 1628 13235
rect 1684 13233 1708 13235
rect 1764 13233 1788 13235
rect 1844 13233 1880 13289
rect 560 13216 612 13222
rect 700 13214 756 13220
rect 612 13212 976 13214
rect 612 13164 702 13212
rect 560 13160 702 13164
rect 754 13160 976 13212
rect 1348 13190 1880 13233
rect 2759 13172 2827 13180
rect 560 13158 1268 13160
rect 700 13152 756 13158
rect 920 13152 1268 13158
rect 2759 13152 2769 13172
rect 920 13120 2769 13152
rect 2821 13120 2827 13172
rect 920 13108 2827 13120
rect 920 13104 1268 13108
rect 852 13062 904 13068
rect 372 12999 378 13054
rect 433 12999 439 13054
rect 1396 13063 2851 13072
rect 3268 13067 3320 13073
rect 1396 13058 3268 13063
rect 904 13028 3268 13058
rect 904 13014 1440 13028
rect 2851 13019 3268 13028
rect 852 13004 904 13010
rect 3268 13009 3320 13015
rect 1930 12982 1990 12993
rect 1004 12970 1056 12976
rect 1930 12971 1932 12982
rect 1056 12959 1242 12966
rect 1599 12959 1932 12971
rect 1056 12937 1932 12959
rect 1056 12925 1633 12937
rect 1930 12926 1932 12937
rect 1988 12971 1990 12982
rect 1988 12937 1991 12971
rect 1988 12926 1990 12937
rect 1056 12922 1242 12925
rect 1004 12912 1056 12918
rect 1930 12915 1990 12926
rect 3564 12907 3605 13617
rect 5029 13453 5035 13505
rect 5087 13453 5093 13505
rect 4744 13386 4796 13392
rect 5047 13380 5075 13453
rect 4796 13341 5075 13380
rect 3724 13288 4264 13330
rect 4744 13328 4796 13334
rect 3724 13232 3766 13288
rect 3822 13286 3846 13288
rect 3902 13286 3926 13288
rect 3982 13286 4006 13288
rect 4062 13286 4086 13288
rect 4142 13286 4166 13288
rect 3828 13234 3840 13286
rect 3902 13234 3904 13286
rect 4084 13234 4086 13286
rect 4148 13234 4160 13286
rect 3822 13232 3846 13234
rect 3902 13232 3926 13234
rect 3982 13232 4006 13234
rect 4062 13232 4086 13234
rect 4142 13232 4166 13234
rect 4222 13232 4264 13288
rect 3724 13190 4264 13232
rect 4291 13061 4346 13067
rect 5016 13061 5068 13064
rect 4291 13059 5084 13061
rect 4291 13007 4292 13059
rect 4344 13058 5084 13059
rect 4344 13007 5016 13058
rect 4291 13006 5016 13007
rect 5068 13006 5084 13058
rect 4291 13000 4346 13006
rect 5016 13000 5068 13006
rect 3561 12901 3613 12907
rect 1154 12883 1209 12889
rect 274 12881 1209 12883
rect 274 12829 1155 12881
rect 1207 12829 1209 12881
rect 274 12828 1209 12829
rect 1154 12822 1209 12828
rect 1754 12884 1814 12890
rect 2267 12884 2325 12893
rect 1754 12881 2325 12884
rect 2838 12881 2898 12886
rect 1754 12880 2898 12881
rect 1754 12828 1758 12880
rect 1810 12878 2908 12880
rect 1810 12828 2270 12878
rect 1754 12826 2270 12828
rect 2322 12876 2908 12878
rect 2322 12826 2842 12876
rect 1754 12824 2842 12826
rect 2894 12824 2908 12876
rect 1754 12818 1814 12824
rect 2267 12823 2908 12824
rect 2267 12811 2325 12823
rect 2838 12820 2908 12823
rect 3262 12822 3268 12874
rect 3320 12822 3326 12874
rect 3976 12892 4028 12898
rect 3561 12843 3613 12849
rect 3975 12843 3976 12886
rect 2838 12814 2898 12820
rect 2768 12780 2816 12784
rect 378 12769 433 12775
rect 1248 12770 1300 12776
rect 433 12766 619 12769
rect 433 12722 1248 12766
rect 433 12714 619 12722
rect 2020 12770 2072 12776
rect 2522 12772 2574 12774
rect 1300 12722 2020 12766
rect 378 12708 433 12714
rect 1248 12712 1300 12718
rect 2020 12712 2072 12718
rect 2509 12770 2587 12772
rect 2509 12714 2520 12770
rect 2576 12714 2587 12770
rect 2760 12728 2766 12780
rect 2818 12776 2824 12780
rect 3270 12776 3314 12822
rect 3564 12804 3605 12843
rect 4622 12851 4628 12903
rect 4680 12851 4686 12903
rect 3976 12834 4028 12840
rect 2818 12732 3314 12776
rect 3979 12787 4018 12834
rect 4637 12787 4671 12851
rect 5122 12804 5164 13617
rect 5202 12907 5244 13952
rect 5197 12901 5249 12907
rect 5197 12843 5249 12849
rect 5202 12804 5244 12843
rect 5282 12804 5324 13952
rect 5362 12804 5404 13952
rect 5442 12804 5484 13952
rect 5522 12804 5564 13952
rect 6820 13948 6872 13954
rect 6974 13950 7026 13956
rect 5662 13826 6202 13868
rect 5662 13770 5704 13826
rect 5760 13824 5784 13826
rect 5840 13824 5864 13826
rect 5920 13824 5944 13826
rect 6000 13824 6024 13826
rect 6080 13824 6104 13826
rect 5766 13772 5778 13824
rect 5840 13772 5842 13824
rect 6022 13772 6024 13824
rect 6086 13772 6098 13824
rect 5760 13770 5784 13772
rect 5840 13770 5864 13772
rect 5920 13770 5944 13772
rect 6000 13770 6024 13772
rect 6080 13770 6104 13772
rect 6160 13770 6202 13826
rect 6504 13824 6510 13876
rect 6562 13824 6568 13876
rect 5662 13728 6202 13770
rect 6518 13660 6556 13824
rect 6523 13590 6553 13660
rect 6506 13538 6512 13590
rect 6564 13538 6570 13590
rect 6843 13386 6895 13392
rect 7196 13380 7235 14444
rect 6895 13341 7235 13380
rect 5682 13288 6222 13330
rect 6843 13328 6895 13334
rect 5682 13232 5724 13288
rect 5780 13286 5804 13288
rect 5860 13286 5884 13288
rect 5940 13286 5964 13288
rect 6020 13286 6044 13288
rect 6100 13286 6124 13288
rect 5786 13234 5798 13286
rect 5860 13234 5862 13286
rect 6042 13234 6044 13286
rect 6106 13234 6118 13286
rect 5780 13232 5804 13234
rect 5860 13232 5884 13234
rect 5940 13232 5964 13234
rect 6020 13232 6044 13234
rect 6100 13232 6124 13234
rect 6180 13232 6222 13288
rect 5682 13190 6222 13232
rect 6250 13062 6304 13068
rect 6974 13062 7026 13064
rect 6250 13060 7042 13062
rect 6302 13058 7042 13060
rect 6302 13008 6974 13058
rect 6250 13006 6974 13008
rect 7026 13006 7042 13058
rect 6250 13000 6304 13006
rect 6974 13000 7026 13006
rect 5934 12892 5986 12898
rect 6580 12852 6586 12904
rect 6638 12852 6644 12904
rect 5934 12834 5986 12840
rect 3979 12748 4673 12787
rect 4862 12778 4914 12784
rect 2818 12728 2824 12732
rect 2509 12712 2587 12714
rect 2522 12710 2574 12712
rect 2768 12688 2812 12728
rect 5015 12780 5067 12786
rect 4914 12738 5015 12767
rect 144 11382 212 12534
rect 274 12461 329 12650
rect 372 12614 378 12670
rect 434 12614 440 12670
rect 274 12455 332 12461
rect 274 12401 278 12455
rect 277 12280 332 12401
rect 378 12442 434 12614
rect 1324 12587 1960 12640
rect 1324 12585 1374 12587
rect 1430 12585 1454 12587
rect 1510 12585 1534 12587
rect 1590 12585 1614 12587
rect 1670 12585 1694 12587
rect 1750 12585 1774 12587
rect 1830 12585 1854 12587
rect 1910 12585 1960 12587
rect 1324 12533 1360 12585
rect 1604 12533 1614 12585
rect 1670 12533 1680 12585
rect 1924 12533 1960 12585
rect 1324 12531 1374 12533
rect 1430 12531 1454 12533
rect 1510 12531 1534 12533
rect 1590 12531 1614 12533
rect 1670 12531 1694 12533
rect 1750 12531 1774 12533
rect 1830 12531 1854 12533
rect 1910 12531 1960 12533
rect 1324 12500 1960 12531
rect 3564 12453 3605 12724
rect 4862 12720 4914 12726
rect 5015 12722 5067 12728
rect 5122 12724 5163 12804
rect 5282 12724 5323 12804
rect 5362 12724 5403 12804
rect 5442 12724 5483 12804
rect 5522 12724 5563 12804
rect 5938 12788 5976 12834
rect 6596 12788 6630 12852
rect 5938 12748 6632 12788
rect 6820 12778 6872 12784
rect 6974 12780 7026 12786
rect 6872 12738 6974 12768
rect 3704 12598 4244 12640
rect 3704 12542 3746 12598
rect 3802 12596 3826 12598
rect 3882 12596 3906 12598
rect 3962 12596 3986 12598
rect 4042 12596 4066 12598
rect 4122 12596 4146 12598
rect 3808 12544 3820 12596
rect 3882 12544 3884 12596
rect 4064 12544 4066 12596
rect 4128 12544 4140 12596
rect 3802 12542 3826 12544
rect 3882 12542 3906 12544
rect 3962 12542 3986 12544
rect 4042 12542 4066 12544
rect 4122 12542 4146 12544
rect 4202 12542 4244 12598
rect 4546 12595 4552 12647
rect 4604 12595 4610 12647
rect 3704 12500 4244 12542
rect 3564 12447 3617 12453
rect 274 11655 329 12280
rect 378 11826 433 12442
rect 3564 12395 3565 12447
rect 4559 12431 4598 12595
rect 3564 12389 3617 12395
rect 1348 12061 1880 12102
rect 1348 12005 1388 12061
rect 1444 12059 1468 12061
rect 1524 12059 1548 12061
rect 1604 12059 1628 12061
rect 1684 12059 1708 12061
rect 1764 12059 1788 12061
rect 1450 12007 1462 12059
rect 1524 12007 1526 12059
rect 1706 12007 1708 12059
rect 1770 12007 1782 12059
rect 1444 12005 1468 12007
rect 1524 12005 1548 12007
rect 1604 12005 1628 12007
rect 1684 12005 1708 12007
rect 1764 12005 1788 12007
rect 1844 12005 1880 12061
rect 560 11988 612 11994
rect 700 11986 756 11992
rect 612 11984 976 11986
rect 612 11936 702 11984
rect 560 11932 702 11936
rect 754 11932 976 11984
rect 1348 11962 1880 12005
rect 2759 11944 2827 11952
rect 560 11930 1268 11932
rect 700 11924 756 11930
rect 920 11924 1268 11930
rect 2759 11924 2769 11944
rect 920 11892 2769 11924
rect 2821 11892 2827 11944
rect 920 11880 2827 11892
rect 920 11876 1268 11880
rect 852 11834 904 11840
rect 372 11771 378 11826
rect 433 11771 439 11826
rect 1396 11835 2851 11844
rect 3268 11839 3320 11845
rect 1396 11830 3268 11835
rect 904 11800 3268 11830
rect 904 11786 1440 11800
rect 2851 11791 3268 11800
rect 852 11776 904 11782
rect 3268 11781 3320 11787
rect 1930 11754 1990 11765
rect 1004 11742 1056 11748
rect 1930 11743 1932 11754
rect 1056 11731 1242 11738
rect 1599 11731 1932 11743
rect 1056 11709 1932 11731
rect 1056 11697 1633 11709
rect 1930 11698 1932 11709
rect 1988 11743 1990 11754
rect 1988 11709 1991 11743
rect 1988 11698 1990 11709
rect 1056 11694 1242 11697
rect 1004 11684 1056 11690
rect 1930 11687 1990 11698
rect 3564 11679 3605 12389
rect 5023 12188 5029 12240
rect 5081 12188 5087 12240
rect 4744 12158 4796 12164
rect 5036 12152 5075 12188
rect 4796 12113 5075 12152
rect 3724 12060 4264 12102
rect 4744 12100 4796 12106
rect 3724 12004 3766 12060
rect 3822 12058 3846 12060
rect 3902 12058 3926 12060
rect 3982 12058 4006 12060
rect 4062 12058 4086 12060
rect 4142 12058 4166 12060
rect 3828 12006 3840 12058
rect 3902 12006 3904 12058
rect 4084 12006 4086 12058
rect 4148 12006 4160 12058
rect 3822 12004 3846 12006
rect 3902 12004 3926 12006
rect 3982 12004 4006 12006
rect 4062 12004 4086 12006
rect 4142 12004 4166 12006
rect 4222 12004 4264 12060
rect 3724 11962 4264 12004
rect 4291 11833 4346 11839
rect 5016 11833 5068 11836
rect 4291 11831 5084 11833
rect 4291 11779 4292 11831
rect 4344 11830 5084 11831
rect 4344 11779 5016 11830
rect 4291 11778 5016 11779
rect 5068 11778 5084 11830
rect 4291 11772 4346 11778
rect 5016 11772 5068 11778
rect 5122 11679 5164 12724
rect 5202 12453 5244 12724
rect 5197 12447 5249 12453
rect 5197 12389 5249 12395
rect 3561 11673 3613 11679
rect 1154 11655 1209 11661
rect 274 11653 1209 11655
rect 274 11601 1155 11653
rect 1207 11601 1209 11653
rect 274 11600 1209 11601
rect 1154 11594 1209 11600
rect 1754 11656 1814 11662
rect 2267 11656 2325 11665
rect 1754 11653 2325 11656
rect 2838 11653 2898 11658
rect 1754 11652 2898 11653
rect 1754 11600 1758 11652
rect 1810 11650 2908 11652
rect 1810 11600 2270 11650
rect 1754 11598 2270 11600
rect 2322 11648 2908 11650
rect 2322 11598 2842 11648
rect 1754 11596 2842 11598
rect 2894 11596 2908 11648
rect 1754 11590 1814 11596
rect 2267 11595 2908 11596
rect 2267 11583 2325 11595
rect 2838 11592 2908 11595
rect 3262 11594 3268 11646
rect 3320 11594 3326 11646
rect 3976 11664 4028 11670
rect 3561 11615 3613 11621
rect 3975 11615 3976 11658
rect 2838 11586 2898 11592
rect 2768 11552 2816 11556
rect 378 11541 433 11547
rect 1248 11542 1300 11548
rect 433 11538 619 11541
rect 433 11494 1248 11538
rect 433 11486 619 11494
rect 2020 11542 2072 11548
rect 2522 11544 2574 11546
rect 1300 11494 2020 11538
rect 378 11480 433 11486
rect 1248 11484 1300 11490
rect 2020 11484 2072 11490
rect 2509 11542 2587 11544
rect 2509 11486 2520 11542
rect 2576 11486 2587 11542
rect 2760 11500 2766 11552
rect 2818 11548 2824 11552
rect 3270 11548 3314 11594
rect 3564 11576 3605 11615
rect 4622 11623 4628 11675
rect 4680 11623 4686 11675
rect 5117 11673 5169 11679
rect 3976 11606 4028 11612
rect 2818 11504 3314 11548
rect 3979 11559 4018 11606
rect 4637 11559 4671 11623
rect 5117 11615 5169 11621
rect 5122 11576 5164 11615
rect 5202 11576 5244 12389
rect 5282 11576 5324 12724
rect 5362 11576 5404 12724
rect 5442 11576 5484 12724
rect 5522 11576 5564 12724
rect 6820 12720 6872 12726
rect 6974 12722 7026 12728
rect 5662 12598 6202 12640
rect 5662 12542 5704 12598
rect 5760 12596 5784 12598
rect 5840 12596 5864 12598
rect 5920 12596 5944 12598
rect 6000 12596 6024 12598
rect 6080 12596 6104 12598
rect 5766 12544 5778 12596
rect 5840 12544 5842 12596
rect 6022 12544 6024 12596
rect 6086 12544 6098 12596
rect 5760 12542 5784 12544
rect 5840 12542 5864 12544
rect 5920 12542 5944 12544
rect 6000 12542 6024 12544
rect 6080 12542 6104 12544
rect 6160 12542 6202 12598
rect 6504 12596 6510 12648
rect 6562 12596 6568 12648
rect 5662 12500 6202 12542
rect 6518 12432 6556 12596
rect 7101 12308 7107 12360
rect 7159 12308 7165 12360
rect 6868 12158 6920 12164
rect 7119 12152 7147 12308
rect 6920 12113 7147 12152
rect 5682 12060 6222 12102
rect 6868 12100 6920 12106
rect 5682 12004 5724 12060
rect 5780 12058 5804 12060
rect 5860 12058 5884 12060
rect 5940 12058 5964 12060
rect 6020 12058 6044 12060
rect 6100 12058 6124 12060
rect 5786 12006 5798 12058
rect 5860 12006 5862 12058
rect 6042 12006 6044 12058
rect 6106 12006 6118 12058
rect 5780 12004 5804 12006
rect 5860 12004 5884 12006
rect 5940 12004 5964 12006
rect 6020 12004 6044 12006
rect 6100 12004 6124 12006
rect 6180 12004 6222 12060
rect 5682 11962 6222 12004
rect 6250 11834 6304 11840
rect 6974 11834 7026 11836
rect 6250 11832 7042 11834
rect 6302 11830 7042 11832
rect 6302 11780 6974 11830
rect 6250 11778 6974 11780
rect 7026 11778 7042 11830
rect 6250 11772 6304 11778
rect 6974 11772 7026 11778
rect 5934 11664 5986 11670
rect 6580 11624 6586 11676
rect 6638 11624 6644 11676
rect 5934 11606 5986 11612
rect 3979 11520 4673 11559
rect 4862 11550 4914 11556
rect 2818 11500 2824 11504
rect 2509 11484 2587 11486
rect 2522 11482 2574 11484
rect 2768 11460 2812 11500
rect 5015 11552 5067 11558
rect 4914 11510 5015 11539
rect 144 10146 212 11314
rect 274 11233 329 11422
rect 372 11386 378 11442
rect 434 11386 440 11442
rect 274 11227 332 11233
rect 274 11173 278 11227
rect 277 11052 332 11173
rect 378 11214 434 11386
rect 1324 11359 1960 11412
rect 1324 11357 1374 11359
rect 1430 11357 1454 11359
rect 1510 11357 1534 11359
rect 1590 11357 1614 11359
rect 1670 11357 1694 11359
rect 1750 11357 1774 11359
rect 1830 11357 1854 11359
rect 1910 11357 1960 11359
rect 1324 11305 1360 11357
rect 1604 11305 1614 11357
rect 1670 11305 1680 11357
rect 1924 11305 1960 11357
rect 1324 11303 1374 11305
rect 1430 11303 1454 11305
rect 1510 11303 1534 11305
rect 1590 11303 1614 11305
rect 1670 11303 1694 11305
rect 1750 11303 1774 11305
rect 1830 11303 1854 11305
rect 1910 11303 1960 11305
rect 1324 11272 1960 11303
rect 3564 11225 3605 11496
rect 4862 11492 4914 11498
rect 5015 11494 5067 11500
rect 5202 11496 5243 11576
rect 5282 11496 5323 11576
rect 5362 11496 5403 11576
rect 5442 11496 5483 11576
rect 5522 11496 5563 11576
rect 5938 11560 5976 11606
rect 6596 11560 6630 11624
rect 5938 11520 6632 11560
rect 6820 11550 6872 11556
rect 6974 11552 7026 11558
rect 6872 11510 6974 11540
rect 3704 11370 4244 11412
rect 3704 11314 3746 11370
rect 3802 11368 3826 11370
rect 3882 11368 3906 11370
rect 3962 11368 3986 11370
rect 4042 11368 4066 11370
rect 4122 11368 4146 11370
rect 3808 11316 3820 11368
rect 3882 11316 3884 11368
rect 4064 11316 4066 11368
rect 4128 11316 4140 11368
rect 3802 11314 3826 11316
rect 3882 11314 3906 11316
rect 3962 11314 3986 11316
rect 4042 11314 4066 11316
rect 4122 11314 4146 11316
rect 4202 11314 4244 11370
rect 4546 11367 4552 11419
rect 4604 11367 4610 11419
rect 3704 11272 4244 11314
rect 3564 11219 3617 11225
rect 274 10427 329 11052
rect 378 10598 433 11214
rect 3564 11167 3565 11219
rect 4559 11203 4598 11367
rect 5122 11225 5164 11496
rect 5117 11219 5169 11225
rect 3564 11161 3617 11167
rect 5117 11161 5169 11167
rect 1348 10833 1880 10874
rect 1348 10777 1388 10833
rect 1444 10831 1468 10833
rect 1524 10831 1548 10833
rect 1604 10831 1628 10833
rect 1684 10831 1708 10833
rect 1764 10831 1788 10833
rect 1450 10779 1462 10831
rect 1524 10779 1526 10831
rect 1706 10779 1708 10831
rect 1770 10779 1782 10831
rect 1444 10777 1468 10779
rect 1524 10777 1548 10779
rect 1604 10777 1628 10779
rect 1684 10777 1708 10779
rect 1764 10777 1788 10779
rect 1844 10777 1880 10833
rect 560 10760 612 10766
rect 700 10758 756 10764
rect 612 10756 976 10758
rect 612 10708 702 10756
rect 560 10704 702 10708
rect 754 10704 976 10756
rect 1348 10734 1880 10777
rect 2759 10716 2827 10724
rect 560 10702 1268 10704
rect 700 10696 756 10702
rect 920 10696 1268 10702
rect 2759 10696 2769 10716
rect 920 10664 2769 10696
rect 2821 10664 2827 10716
rect 920 10652 2827 10664
rect 920 10648 1268 10652
rect 852 10606 904 10612
rect 372 10543 378 10598
rect 433 10543 439 10598
rect 1396 10607 2851 10616
rect 3268 10611 3320 10617
rect 1396 10602 3268 10607
rect 904 10572 3268 10602
rect 904 10558 1440 10572
rect 2851 10563 3268 10572
rect 852 10548 904 10554
rect 3268 10553 3320 10559
rect 1930 10526 1990 10537
rect 1004 10514 1056 10520
rect 1930 10515 1932 10526
rect 1056 10503 1242 10510
rect 1599 10503 1932 10515
rect 1056 10481 1932 10503
rect 1056 10469 1633 10481
rect 1930 10470 1932 10481
rect 1988 10515 1990 10526
rect 1988 10481 1991 10515
rect 1988 10470 1990 10481
rect 1056 10466 1242 10469
rect 1004 10456 1056 10462
rect 1930 10459 1990 10470
rect 3564 10451 3605 11161
rect 5029 10997 5035 11049
rect 5087 10997 5093 11049
rect 4744 10930 4796 10936
rect 5047 10924 5075 10997
rect 4796 10885 5075 10924
rect 3724 10832 4264 10874
rect 4744 10872 4796 10878
rect 3724 10776 3766 10832
rect 3822 10830 3846 10832
rect 3902 10830 3926 10832
rect 3982 10830 4006 10832
rect 4062 10830 4086 10832
rect 4142 10830 4166 10832
rect 3828 10778 3840 10830
rect 3902 10778 3904 10830
rect 4084 10778 4086 10830
rect 4148 10778 4160 10830
rect 3822 10776 3846 10778
rect 3902 10776 3926 10778
rect 3982 10776 4006 10778
rect 4062 10776 4086 10778
rect 4142 10776 4166 10778
rect 4222 10776 4264 10832
rect 3724 10734 4264 10776
rect 4291 10605 4346 10611
rect 5016 10605 5068 10608
rect 4291 10603 5084 10605
rect 4291 10551 4292 10603
rect 4344 10602 5084 10603
rect 4344 10551 5016 10602
rect 4291 10550 5016 10551
rect 5068 10550 5084 10602
rect 4291 10544 4346 10550
rect 5016 10544 5068 10550
rect 3561 10445 3613 10451
rect 1154 10427 1209 10433
rect 274 10425 1209 10427
rect 274 10373 1155 10425
rect 1207 10373 1209 10425
rect 274 10372 1209 10373
rect 1154 10366 1209 10372
rect 1754 10428 1814 10434
rect 2267 10428 2325 10437
rect 1754 10425 2325 10428
rect 2838 10425 2898 10430
rect 1754 10424 2898 10425
rect 1754 10372 1758 10424
rect 1810 10422 2908 10424
rect 1810 10372 2270 10422
rect 1754 10370 2270 10372
rect 2322 10420 2908 10422
rect 2322 10370 2842 10420
rect 1754 10368 2842 10370
rect 2894 10368 2908 10420
rect 1754 10362 1814 10368
rect 2267 10367 2908 10368
rect 2267 10355 2325 10367
rect 2838 10364 2908 10367
rect 3262 10366 3268 10418
rect 3320 10366 3326 10418
rect 3976 10436 4028 10442
rect 3561 10387 3613 10393
rect 3975 10387 3976 10430
rect 2838 10358 2898 10364
rect 2768 10324 2816 10328
rect 378 10313 433 10319
rect 1248 10314 1300 10320
rect 433 10310 619 10313
rect 433 10266 1248 10310
rect 433 10258 619 10266
rect 2020 10314 2072 10320
rect 2522 10316 2574 10318
rect 1300 10266 2020 10310
rect 378 10252 433 10258
rect 1248 10256 1300 10262
rect 2020 10256 2072 10262
rect 2509 10314 2587 10316
rect 2509 10258 2520 10314
rect 2576 10258 2587 10314
rect 2760 10272 2766 10324
rect 2818 10320 2824 10324
rect 3270 10320 3314 10366
rect 3564 10348 3605 10387
rect 4622 10395 4628 10447
rect 4680 10395 4686 10447
rect 3976 10378 4028 10384
rect 2818 10276 3314 10320
rect 3979 10331 4018 10378
rect 4637 10331 4671 10395
rect 5122 10348 5164 11161
rect 5202 10348 5244 11496
rect 5282 10348 5324 11496
rect 5362 10451 5404 11496
rect 5356 10445 5408 10451
rect 5356 10387 5408 10393
rect 5362 10348 5404 10387
rect 5442 10348 5484 11496
rect 5522 10348 5564 11496
rect 6820 11492 6872 11498
rect 6974 11494 7026 11500
rect 5662 11370 6202 11412
rect 5662 11314 5704 11370
rect 5760 11368 5784 11370
rect 5840 11368 5864 11370
rect 5920 11368 5944 11370
rect 6000 11368 6024 11370
rect 6080 11368 6104 11370
rect 5766 11316 5778 11368
rect 5840 11316 5842 11368
rect 6022 11316 6024 11368
rect 6086 11316 6098 11368
rect 5760 11314 5784 11316
rect 5840 11314 5864 11316
rect 5920 11314 5944 11316
rect 6000 11314 6024 11316
rect 6080 11314 6104 11316
rect 6160 11314 6202 11370
rect 6504 11368 6510 11420
rect 6562 11368 6568 11420
rect 5662 11272 6202 11314
rect 6518 11204 6556 11368
rect 6974 11022 7026 11028
rect 7298 11011 7337 14887
rect 7026 10981 7337 11011
rect 6974 10964 7026 10970
rect 6835 10930 6887 10936
rect 6887 10885 7150 10924
rect 5682 10832 6222 10874
rect 6835 10872 6887 10878
rect 5682 10776 5724 10832
rect 5780 10830 5804 10832
rect 5860 10830 5884 10832
rect 5940 10830 5964 10832
rect 6020 10830 6044 10832
rect 6100 10830 6124 10832
rect 5786 10778 5798 10830
rect 5860 10778 5862 10830
rect 6042 10778 6044 10830
rect 6106 10778 6118 10830
rect 5780 10776 5804 10778
rect 5860 10776 5884 10778
rect 5940 10776 5964 10778
rect 6020 10776 6044 10778
rect 6100 10776 6124 10778
rect 6180 10776 6222 10832
rect 5682 10734 6222 10776
rect 7111 10802 7150 10885
rect 7111 10763 7360 10802
rect 6250 10606 6304 10612
rect 6974 10606 7026 10608
rect 6250 10604 7042 10606
rect 6302 10602 7042 10604
rect 6302 10552 6974 10602
rect 6250 10550 6974 10552
rect 7026 10550 7042 10602
rect 6250 10544 6304 10550
rect 6974 10544 7026 10550
rect 5934 10436 5986 10442
rect 6580 10396 6586 10448
rect 6638 10396 6644 10448
rect 5934 10378 5986 10384
rect 3979 10292 4673 10331
rect 4862 10322 4914 10328
rect 2818 10272 2824 10276
rect 2509 10256 2587 10258
rect 2522 10254 2574 10256
rect 2768 10232 2812 10272
rect 5015 10324 5067 10330
rect 4914 10282 5015 10311
rect 144 8926 212 10078
rect 274 10037 329 10194
rect 372 10158 378 10214
rect 434 10158 440 10214
rect 274 9999 332 10037
rect 274 9945 278 9999
rect 277 9824 332 9945
rect 378 9986 434 10158
rect 1324 10131 1960 10184
rect 1324 10129 1374 10131
rect 1430 10129 1454 10131
rect 1510 10129 1534 10131
rect 1590 10129 1614 10131
rect 1670 10129 1694 10131
rect 1750 10129 1774 10131
rect 1830 10129 1854 10131
rect 1910 10129 1960 10131
rect 1324 10077 1360 10129
rect 1604 10077 1614 10129
rect 1670 10077 1680 10129
rect 1924 10077 1960 10129
rect 1324 10075 1374 10077
rect 1430 10075 1454 10077
rect 1510 10075 1534 10077
rect 1590 10075 1614 10077
rect 1670 10075 1694 10077
rect 1750 10075 1774 10077
rect 1830 10075 1854 10077
rect 1910 10075 1960 10077
rect 1324 10044 1960 10075
rect 3564 9997 3605 10268
rect 4862 10264 4914 10270
rect 5015 10266 5067 10272
rect 5122 10268 5163 10348
rect 5202 10268 5243 10348
rect 5282 10268 5323 10348
rect 5442 10268 5483 10348
rect 5522 10268 5563 10348
rect 5938 10332 5976 10378
rect 6596 10332 6630 10396
rect 5938 10292 6632 10332
rect 6820 10322 6872 10328
rect 6974 10324 7026 10330
rect 6872 10282 6974 10312
rect 3704 10142 4244 10184
rect 3704 10086 3746 10142
rect 3802 10140 3826 10142
rect 3882 10140 3906 10142
rect 3962 10140 3986 10142
rect 4042 10140 4066 10142
rect 4122 10140 4146 10142
rect 3808 10088 3820 10140
rect 3882 10088 3884 10140
rect 4064 10088 4066 10140
rect 4128 10088 4140 10140
rect 3802 10086 3826 10088
rect 3882 10086 3906 10088
rect 3962 10086 3986 10088
rect 4042 10086 4066 10088
rect 4122 10086 4146 10088
rect 4202 10086 4244 10142
rect 4546 10139 4552 10191
rect 4604 10139 4610 10191
rect 3704 10044 4244 10086
rect 3564 9991 3617 9997
rect 274 9199 329 9824
rect 378 9370 433 9986
rect 3564 9939 3565 9991
rect 4559 9975 4598 10139
rect 3564 9933 3617 9939
rect 1348 9605 1880 9646
rect 1348 9549 1388 9605
rect 1444 9603 1468 9605
rect 1524 9603 1548 9605
rect 1604 9603 1628 9605
rect 1684 9603 1708 9605
rect 1764 9603 1788 9605
rect 1450 9551 1462 9603
rect 1524 9551 1526 9603
rect 1706 9551 1708 9603
rect 1770 9551 1782 9603
rect 1444 9549 1468 9551
rect 1524 9549 1548 9551
rect 1604 9549 1628 9551
rect 1684 9549 1708 9551
rect 1764 9549 1788 9551
rect 1844 9549 1880 9605
rect 560 9532 612 9538
rect 700 9530 756 9536
rect 612 9528 976 9530
rect 612 9480 702 9528
rect 560 9476 702 9480
rect 754 9476 976 9528
rect 1348 9506 1880 9549
rect 2759 9488 2827 9496
rect 560 9474 1268 9476
rect 700 9468 756 9474
rect 920 9468 1268 9474
rect 2759 9468 2769 9488
rect 920 9436 2769 9468
rect 2821 9436 2827 9488
rect 920 9424 2827 9436
rect 920 9420 1268 9424
rect 852 9378 904 9384
rect 372 9315 378 9370
rect 433 9315 439 9370
rect 1396 9379 2851 9388
rect 3268 9383 3320 9389
rect 1396 9374 3268 9379
rect 904 9344 3268 9374
rect 904 9330 1440 9344
rect 2851 9335 3268 9344
rect 852 9320 904 9326
rect 3268 9325 3320 9331
rect 1930 9298 1990 9309
rect 1004 9286 1056 9292
rect 1930 9287 1932 9298
rect 1056 9275 1242 9282
rect 1599 9275 1932 9287
rect 1056 9253 1932 9275
rect 1056 9241 1633 9253
rect 1930 9242 1932 9253
rect 1988 9287 1990 9298
rect 1988 9253 1991 9287
rect 1988 9242 1990 9253
rect 1056 9238 1242 9241
rect 1004 9228 1056 9234
rect 1930 9231 1990 9242
rect 3564 9223 3605 9933
rect 5023 9732 5029 9784
rect 5081 9732 5087 9784
rect 4744 9702 4796 9708
rect 5036 9696 5075 9732
rect 4796 9657 5075 9696
rect 3724 9604 4264 9646
rect 4744 9644 4796 9650
rect 3724 9548 3766 9604
rect 3822 9602 3846 9604
rect 3902 9602 3926 9604
rect 3982 9602 4006 9604
rect 4062 9602 4086 9604
rect 4142 9602 4166 9604
rect 3828 9550 3840 9602
rect 3902 9550 3904 9602
rect 4084 9550 4086 9602
rect 4148 9550 4160 9602
rect 3822 9548 3846 9550
rect 3902 9548 3926 9550
rect 3982 9548 4006 9550
rect 4062 9548 4086 9550
rect 4142 9548 4166 9550
rect 4222 9548 4264 9604
rect 3724 9506 4264 9548
rect 4291 9377 4346 9383
rect 5016 9377 5068 9380
rect 4291 9375 5084 9377
rect 4291 9323 4292 9375
rect 4344 9374 5084 9375
rect 4344 9323 5016 9374
rect 4291 9322 5016 9323
rect 5068 9322 5084 9374
rect 4291 9316 4346 9322
rect 5016 9316 5068 9322
rect 5122 9223 5164 10268
rect 3561 9217 3613 9223
rect 1154 9199 1209 9205
rect 274 9197 1209 9199
rect 274 9145 1155 9197
rect 1207 9145 1209 9197
rect 274 9144 1209 9145
rect 1154 9138 1209 9144
rect 1754 9200 1814 9206
rect 2267 9200 2325 9209
rect 1754 9197 2325 9200
rect 2838 9197 2898 9202
rect 1754 9196 2898 9197
rect 1754 9144 1758 9196
rect 1810 9194 2908 9196
rect 1810 9144 2270 9194
rect 1754 9142 2270 9144
rect 2322 9192 2908 9194
rect 2322 9142 2842 9192
rect 1754 9140 2842 9142
rect 2894 9140 2908 9192
rect 1754 9134 1814 9140
rect 2267 9139 2908 9140
rect 2267 9127 2325 9139
rect 2838 9136 2908 9139
rect 3262 9138 3268 9190
rect 3320 9138 3326 9190
rect 3976 9208 4028 9214
rect 3561 9159 3613 9165
rect 3975 9159 3976 9202
rect 2838 9130 2898 9136
rect 2768 9096 2816 9100
rect 378 9085 433 9091
rect 1248 9086 1300 9092
rect 433 9082 619 9085
rect 433 9038 1248 9082
rect 433 9030 619 9038
rect 2020 9086 2072 9092
rect 2522 9088 2574 9090
rect 1300 9038 2020 9082
rect 378 9024 433 9030
rect 1248 9028 1300 9034
rect 2020 9028 2072 9034
rect 2509 9086 2587 9088
rect 2509 9030 2520 9086
rect 2576 9030 2587 9086
rect 2760 9044 2766 9096
rect 2818 9092 2824 9096
rect 3270 9092 3314 9138
rect 3564 9120 3605 9159
rect 4622 9167 4628 9219
rect 4680 9167 4686 9219
rect 5117 9217 5169 9223
rect 3976 9150 4028 9156
rect 2818 9048 3314 9092
rect 3979 9103 4018 9150
rect 4637 9103 4671 9167
rect 5117 9159 5169 9165
rect 5122 9120 5164 9159
rect 5202 9120 5244 10268
rect 5282 9120 5324 10268
rect 5362 9997 5404 10268
rect 5354 9991 5406 9997
rect 5354 9933 5406 9939
rect 5362 9120 5404 9933
rect 5442 9120 5484 10268
rect 5522 9120 5564 10268
rect 6820 10264 6872 10270
rect 6974 10266 7026 10272
rect 5662 10142 6202 10184
rect 5662 10086 5704 10142
rect 5760 10140 5784 10142
rect 5840 10140 5864 10142
rect 5920 10140 5944 10142
rect 6000 10140 6024 10142
rect 6080 10140 6104 10142
rect 5766 10088 5778 10140
rect 5840 10088 5842 10140
rect 6022 10088 6024 10140
rect 6086 10088 6098 10140
rect 5760 10086 5784 10088
rect 5840 10086 5864 10088
rect 5920 10086 5944 10088
rect 6000 10086 6024 10088
rect 6080 10086 6104 10088
rect 6160 10086 6202 10142
rect 6504 10140 6510 10192
rect 6562 10140 6568 10192
rect 5662 10044 6202 10086
rect 6518 9976 6556 10140
rect 7085 10010 7137 10016
rect 7137 9970 7322 9998
rect 7085 9952 7137 9958
rect 6868 9702 6920 9708
rect 6920 9657 7147 9696
rect 5682 9604 6222 9646
rect 6868 9644 6920 9650
rect 5682 9548 5724 9604
rect 5780 9602 5804 9604
rect 5860 9602 5884 9604
rect 5940 9602 5964 9604
rect 6020 9602 6044 9604
rect 6100 9602 6124 9604
rect 5786 9550 5798 9602
rect 5860 9550 5862 9602
rect 6042 9550 6044 9602
rect 6106 9550 6118 9602
rect 5780 9548 5804 9550
rect 5860 9548 5884 9550
rect 5940 9548 5964 9550
rect 6020 9548 6044 9550
rect 6100 9548 6124 9550
rect 6180 9548 6222 9604
rect 5682 9506 6222 9548
rect 6250 9378 6304 9384
rect 6974 9378 7026 9380
rect 6250 9376 7042 9378
rect 6302 9374 7042 9376
rect 6302 9324 6974 9374
rect 6250 9322 6974 9324
rect 7026 9322 7042 9374
rect 6250 9316 6304 9322
rect 6974 9316 7026 9322
rect 5934 9208 5986 9214
rect 6580 9168 6586 9220
rect 6638 9168 6644 9220
rect 5934 9150 5986 9156
rect 3979 9064 4673 9103
rect 4862 9094 4914 9100
rect 2818 9044 2824 9048
rect 2509 9028 2587 9030
rect 2522 9026 2574 9028
rect 2768 9004 2812 9044
rect 5015 9096 5067 9102
rect 4914 9054 5015 9083
rect 144 7690 212 8858
rect 274 8777 329 8966
rect 372 8930 378 8986
rect 434 8930 440 8986
rect 274 8771 332 8777
rect 274 8717 278 8771
rect 277 8596 332 8717
rect 378 8758 434 8930
rect 1324 8903 1960 8956
rect 1324 8901 1374 8903
rect 1430 8901 1454 8903
rect 1510 8901 1534 8903
rect 1590 8901 1614 8903
rect 1670 8901 1694 8903
rect 1750 8901 1774 8903
rect 1830 8901 1854 8903
rect 1910 8901 1960 8903
rect 1324 8849 1360 8901
rect 1604 8849 1614 8901
rect 1670 8849 1680 8901
rect 1924 8849 1960 8901
rect 1324 8847 1374 8849
rect 1430 8847 1454 8849
rect 1510 8847 1534 8849
rect 1590 8847 1614 8849
rect 1670 8847 1694 8849
rect 1750 8847 1774 8849
rect 1830 8847 1854 8849
rect 1910 8847 1960 8849
rect 1324 8816 1960 8847
rect 3564 8769 3605 9040
rect 4862 9036 4914 9042
rect 5015 9038 5067 9044
rect 5202 9040 5243 9120
rect 5282 9040 5323 9120
rect 5362 9040 5403 9120
rect 5442 9040 5483 9120
rect 5522 9040 5563 9120
rect 5938 9104 5976 9150
rect 6596 9104 6630 9168
rect 5938 9064 6632 9104
rect 6820 9094 6872 9100
rect 6974 9096 7026 9102
rect 6872 9054 6974 9084
rect 3704 8914 4244 8956
rect 3704 8858 3746 8914
rect 3802 8912 3826 8914
rect 3882 8912 3906 8914
rect 3962 8912 3986 8914
rect 4042 8912 4066 8914
rect 4122 8912 4146 8914
rect 3808 8860 3820 8912
rect 3882 8860 3884 8912
rect 4064 8860 4066 8912
rect 4128 8860 4140 8912
rect 3802 8858 3826 8860
rect 3882 8858 3906 8860
rect 3962 8858 3986 8860
rect 4042 8858 4066 8860
rect 4122 8858 4146 8860
rect 4202 8858 4244 8914
rect 4546 8911 4552 8963
rect 4604 8911 4610 8963
rect 3704 8816 4244 8858
rect 3564 8763 3617 8769
rect 274 7971 329 8596
rect 378 8142 433 8758
rect 3564 8711 3565 8763
rect 4559 8747 4598 8911
rect 5122 8769 5164 9040
rect 5117 8763 5169 8769
rect 3564 8705 3617 8711
rect 5117 8705 5169 8711
rect 1348 8377 1880 8418
rect 1348 8321 1388 8377
rect 1444 8375 1468 8377
rect 1524 8375 1548 8377
rect 1604 8375 1628 8377
rect 1684 8375 1708 8377
rect 1764 8375 1788 8377
rect 1450 8323 1462 8375
rect 1524 8323 1526 8375
rect 1706 8323 1708 8375
rect 1770 8323 1782 8375
rect 1444 8321 1468 8323
rect 1524 8321 1548 8323
rect 1604 8321 1628 8323
rect 1684 8321 1708 8323
rect 1764 8321 1788 8323
rect 1844 8321 1880 8377
rect 560 8304 612 8310
rect 700 8302 756 8308
rect 612 8300 976 8302
rect 612 8252 702 8300
rect 560 8248 702 8252
rect 754 8248 976 8300
rect 1348 8278 1880 8321
rect 2759 8260 2827 8268
rect 560 8246 1268 8248
rect 700 8240 756 8246
rect 920 8240 1268 8246
rect 2759 8240 2769 8260
rect 920 8208 2769 8240
rect 2821 8208 2827 8260
rect 920 8196 2827 8208
rect 920 8192 1268 8196
rect 852 8150 904 8156
rect 372 8087 378 8142
rect 433 8087 439 8142
rect 1396 8151 2851 8160
rect 3268 8155 3320 8161
rect 1396 8146 3268 8151
rect 904 8116 3268 8146
rect 904 8102 1440 8116
rect 2851 8107 3268 8116
rect 852 8092 904 8098
rect 3268 8097 3320 8103
rect 1930 8070 1990 8081
rect 1004 8058 1056 8064
rect 1930 8059 1932 8070
rect 1056 8047 1242 8054
rect 1599 8047 1932 8059
rect 1056 8025 1932 8047
rect 1056 8013 1633 8025
rect 1930 8014 1932 8025
rect 1988 8059 1990 8070
rect 1988 8025 1991 8059
rect 1988 8014 1990 8025
rect 1056 8010 1242 8013
rect 1004 8000 1056 8006
rect 1930 8003 1990 8014
rect 3564 7995 3605 8705
rect 5029 8541 5035 8593
rect 5087 8541 5093 8593
rect 4744 8474 4796 8480
rect 5047 8468 5075 8541
rect 4796 8429 5075 8468
rect 3724 8376 4264 8418
rect 4744 8416 4796 8422
rect 3724 8320 3766 8376
rect 3822 8374 3846 8376
rect 3902 8374 3926 8376
rect 3982 8374 4006 8376
rect 4062 8374 4086 8376
rect 4142 8374 4166 8376
rect 3828 8322 3840 8374
rect 3902 8322 3904 8374
rect 4084 8322 4086 8374
rect 4148 8322 4160 8374
rect 3822 8320 3846 8322
rect 3902 8320 3926 8322
rect 3982 8320 4006 8322
rect 4062 8320 4086 8322
rect 4142 8320 4166 8322
rect 4222 8320 4264 8376
rect 3724 8278 4264 8320
rect 4291 8149 4346 8155
rect 5016 8149 5068 8152
rect 4291 8147 5084 8149
rect 4291 8095 4292 8147
rect 4344 8146 5084 8147
rect 4344 8095 5016 8146
rect 4291 8094 5016 8095
rect 5068 8094 5084 8146
rect 4291 8088 4346 8094
rect 5016 8088 5068 8094
rect 3561 7989 3613 7995
rect 1154 7971 1209 7977
rect 274 7969 1209 7971
rect 274 7917 1155 7969
rect 1207 7917 1209 7969
rect 274 7916 1209 7917
rect 1154 7910 1209 7916
rect 1754 7972 1814 7978
rect 2267 7972 2325 7981
rect 1754 7969 2325 7972
rect 2838 7969 2898 7974
rect 1754 7968 2898 7969
rect 1754 7916 1758 7968
rect 1810 7966 2908 7968
rect 1810 7916 2270 7966
rect 1754 7914 2270 7916
rect 2322 7964 2908 7966
rect 2322 7914 2842 7964
rect 1754 7912 2842 7914
rect 2894 7912 2908 7964
rect 1754 7906 1814 7912
rect 2267 7911 2908 7912
rect 2267 7899 2325 7911
rect 2838 7908 2908 7911
rect 3262 7910 3268 7962
rect 3320 7910 3326 7962
rect 3976 7980 4028 7986
rect 3561 7931 3613 7937
rect 3975 7931 3976 7974
rect 2838 7902 2898 7908
rect 2768 7868 2816 7872
rect 378 7857 433 7863
rect 1248 7858 1300 7864
rect 433 7854 619 7857
rect 433 7810 1248 7854
rect 433 7802 619 7810
rect 2020 7858 2072 7864
rect 2522 7860 2574 7862
rect 1300 7810 2020 7854
rect 378 7796 433 7802
rect 1248 7800 1300 7806
rect 2020 7800 2072 7806
rect 2509 7858 2587 7860
rect 2509 7802 2520 7858
rect 2576 7802 2587 7858
rect 2760 7816 2766 7868
rect 2818 7864 2824 7868
rect 3270 7864 3314 7910
rect 3564 7892 3605 7931
rect 4622 7939 4628 7991
rect 4680 7939 4686 7991
rect 3976 7922 4028 7928
rect 2818 7820 3314 7864
rect 3979 7875 4018 7922
rect 4637 7875 4671 7939
rect 5122 7892 5164 8705
rect 5202 7995 5244 9040
rect 5197 7989 5249 7995
rect 5197 7931 5249 7937
rect 5202 7892 5244 7931
rect 5282 7892 5324 9040
rect 5362 7892 5404 9040
rect 5442 7892 5484 9040
rect 5522 7892 5564 9040
rect 6820 9036 6872 9042
rect 6974 9038 7026 9044
rect 5662 8914 6202 8956
rect 5662 8858 5704 8914
rect 5760 8912 5784 8914
rect 5840 8912 5864 8914
rect 5920 8912 5944 8914
rect 6000 8912 6024 8914
rect 6080 8912 6104 8914
rect 5766 8860 5778 8912
rect 5840 8860 5842 8912
rect 6022 8860 6024 8912
rect 6086 8860 6098 8912
rect 5760 8858 5784 8860
rect 5840 8858 5864 8860
rect 5920 8858 5944 8860
rect 6000 8858 6024 8860
rect 6080 8858 6104 8860
rect 6160 8858 6202 8914
rect 6504 8912 6510 8964
rect 6562 8912 6568 8964
rect 5662 8816 6202 8858
rect 6518 8748 6556 8912
rect 6523 8678 6553 8748
rect 6506 8626 6512 8678
rect 6564 8626 6570 8678
rect 6843 8474 6895 8480
rect 6895 8429 7241 8468
rect 5682 8376 6222 8418
rect 6843 8416 6895 8422
rect 5682 8320 5724 8376
rect 5780 8374 5804 8376
rect 5860 8374 5884 8376
rect 5940 8374 5964 8376
rect 6020 8374 6044 8376
rect 6100 8374 6124 8376
rect 5786 8322 5798 8374
rect 5860 8322 5862 8374
rect 6042 8322 6044 8374
rect 6106 8322 6118 8374
rect 5780 8320 5804 8322
rect 5860 8320 5884 8322
rect 5940 8320 5964 8322
rect 6020 8320 6044 8322
rect 6100 8320 6124 8322
rect 6180 8320 6222 8376
rect 5682 8278 6222 8320
rect 6250 8150 6304 8156
rect 6974 8150 7026 8152
rect 6250 8148 7042 8150
rect 6302 8146 7042 8148
rect 6302 8096 6974 8146
rect 6250 8094 6974 8096
rect 7026 8094 7042 8146
rect 6250 8088 6304 8094
rect 6974 8088 7026 8094
rect 5934 7980 5986 7986
rect 6580 7940 6586 7992
rect 6638 7940 6644 7992
rect 5934 7922 5986 7928
rect 3979 7836 4673 7875
rect 4862 7866 4914 7872
rect 2818 7816 2824 7820
rect 2509 7800 2587 7802
rect 2522 7798 2574 7800
rect 2768 7776 2812 7816
rect 5015 7868 5067 7874
rect 4914 7826 5015 7855
rect 144 6470 212 7622
rect 274 7549 329 7738
rect 372 7702 378 7758
rect 434 7702 440 7758
rect 274 7543 332 7549
rect 274 7489 278 7543
rect 277 7368 332 7489
rect 378 7530 434 7702
rect 1324 7675 1960 7728
rect 1324 7673 1374 7675
rect 1430 7673 1454 7675
rect 1510 7673 1534 7675
rect 1590 7673 1614 7675
rect 1670 7673 1694 7675
rect 1750 7673 1774 7675
rect 1830 7673 1854 7675
rect 1910 7673 1960 7675
rect 1324 7621 1360 7673
rect 1604 7621 1614 7673
rect 1670 7621 1680 7673
rect 1924 7621 1960 7673
rect 1324 7619 1374 7621
rect 1430 7619 1454 7621
rect 1510 7619 1534 7621
rect 1590 7619 1614 7621
rect 1670 7619 1694 7621
rect 1750 7619 1774 7621
rect 1830 7619 1854 7621
rect 1910 7619 1960 7621
rect 1324 7588 1960 7619
rect 3564 7541 3605 7812
rect 4862 7808 4914 7814
rect 5015 7810 5067 7816
rect 5122 7812 5163 7892
rect 5282 7812 5323 7892
rect 5362 7812 5403 7892
rect 5442 7812 5483 7892
rect 5522 7812 5563 7892
rect 5938 7876 5976 7922
rect 6596 7876 6630 7940
rect 5938 7836 6632 7876
rect 6820 7866 6872 7872
rect 6974 7868 7026 7874
rect 6872 7826 6974 7856
rect 3704 7686 4244 7728
rect 3704 7630 3746 7686
rect 3802 7684 3826 7686
rect 3882 7684 3906 7686
rect 3962 7684 3986 7686
rect 4042 7684 4066 7686
rect 4122 7684 4146 7686
rect 3808 7632 3820 7684
rect 3882 7632 3884 7684
rect 4064 7632 4066 7684
rect 4128 7632 4140 7684
rect 3802 7630 3826 7632
rect 3882 7630 3906 7632
rect 3962 7630 3986 7632
rect 4042 7630 4066 7632
rect 4122 7630 4146 7632
rect 4202 7630 4244 7686
rect 4546 7683 4552 7735
rect 4604 7683 4610 7735
rect 3704 7588 4244 7630
rect 3564 7535 3617 7541
rect 274 6743 329 7368
rect 378 6914 433 7530
rect 3564 7483 3565 7535
rect 4559 7519 4598 7683
rect 3564 7477 3617 7483
rect 1348 7149 1880 7190
rect 1348 7093 1388 7149
rect 1444 7147 1468 7149
rect 1524 7147 1548 7149
rect 1604 7147 1628 7149
rect 1684 7147 1708 7149
rect 1764 7147 1788 7149
rect 1450 7095 1462 7147
rect 1524 7095 1526 7147
rect 1706 7095 1708 7147
rect 1770 7095 1782 7147
rect 1444 7093 1468 7095
rect 1524 7093 1548 7095
rect 1604 7093 1628 7095
rect 1684 7093 1708 7095
rect 1764 7093 1788 7095
rect 1844 7093 1880 7149
rect 560 7076 612 7082
rect 700 7074 756 7080
rect 612 7072 976 7074
rect 612 7024 702 7072
rect 560 7020 702 7024
rect 754 7020 976 7072
rect 1348 7050 1880 7093
rect 2759 7032 2827 7040
rect 560 7018 1268 7020
rect 700 7012 756 7018
rect 920 7012 1268 7018
rect 2759 7012 2769 7032
rect 920 6980 2769 7012
rect 2821 6980 2827 7032
rect 920 6968 2827 6980
rect 920 6964 1268 6968
rect 852 6922 904 6928
rect 372 6859 378 6914
rect 433 6859 439 6914
rect 1396 6923 2851 6932
rect 3268 6927 3320 6933
rect 1396 6918 3268 6923
rect 904 6888 3268 6918
rect 904 6874 1440 6888
rect 2851 6879 3268 6888
rect 852 6864 904 6870
rect 3268 6869 3320 6875
rect 1930 6842 1990 6853
rect 1004 6830 1056 6836
rect 1930 6831 1932 6842
rect 1056 6819 1242 6826
rect 1599 6819 1932 6831
rect 1056 6797 1932 6819
rect 1056 6785 1633 6797
rect 1930 6786 1932 6797
rect 1988 6831 1990 6842
rect 1988 6797 1991 6831
rect 1988 6786 1990 6797
rect 1056 6782 1242 6785
rect 1004 6772 1056 6778
rect 1930 6775 1990 6786
rect 3564 6767 3605 7477
rect 5023 7276 5029 7328
rect 5081 7276 5087 7328
rect 4744 7246 4796 7252
rect 5036 7240 5075 7276
rect 4796 7201 5075 7240
rect 3724 7148 4264 7190
rect 4744 7188 4796 7194
rect 3724 7092 3766 7148
rect 3822 7146 3846 7148
rect 3902 7146 3926 7148
rect 3982 7146 4006 7148
rect 4062 7146 4086 7148
rect 4142 7146 4166 7148
rect 3828 7094 3840 7146
rect 3902 7094 3904 7146
rect 4084 7094 4086 7146
rect 4148 7094 4160 7146
rect 3822 7092 3846 7094
rect 3902 7092 3926 7094
rect 3982 7092 4006 7094
rect 4062 7092 4086 7094
rect 4142 7092 4166 7094
rect 4222 7092 4264 7148
rect 3724 7050 4264 7092
rect 4291 6921 4346 6927
rect 5016 6921 5068 6924
rect 4291 6919 5084 6921
rect 4291 6867 4292 6919
rect 4344 6918 5084 6919
rect 4344 6867 5016 6918
rect 4291 6866 5016 6867
rect 5068 6866 5084 6918
rect 4291 6860 4346 6866
rect 5016 6860 5068 6866
rect 5122 6767 5164 7812
rect 5202 7541 5244 7812
rect 5197 7535 5249 7541
rect 5197 7477 5249 7483
rect 3561 6761 3613 6767
rect 1154 6743 1209 6749
rect 274 6741 1209 6743
rect 274 6689 1155 6741
rect 1207 6689 1209 6741
rect 274 6688 1209 6689
rect 1154 6682 1209 6688
rect 1754 6744 1814 6750
rect 2267 6744 2325 6753
rect 1754 6741 2325 6744
rect 2838 6741 2898 6746
rect 1754 6740 2898 6741
rect 1754 6688 1758 6740
rect 1810 6738 2908 6740
rect 1810 6688 2270 6738
rect 1754 6686 2270 6688
rect 2322 6736 2908 6738
rect 2322 6686 2842 6736
rect 1754 6684 2842 6686
rect 2894 6684 2908 6736
rect 1754 6678 1814 6684
rect 2267 6683 2908 6684
rect 2267 6671 2325 6683
rect 2838 6680 2908 6683
rect 3262 6682 3268 6734
rect 3320 6682 3326 6734
rect 3976 6752 4028 6758
rect 3561 6703 3613 6709
rect 3975 6703 3976 6746
rect 2838 6674 2898 6680
rect 2768 6640 2816 6644
rect 378 6629 433 6635
rect 1248 6630 1300 6636
rect 433 6626 619 6629
rect 433 6582 1248 6626
rect 433 6574 619 6582
rect 2020 6630 2072 6636
rect 2522 6632 2574 6634
rect 1300 6582 2020 6626
rect 378 6568 433 6574
rect 1248 6572 1300 6578
rect 2020 6572 2072 6578
rect 2509 6630 2587 6632
rect 2509 6574 2520 6630
rect 2576 6574 2587 6630
rect 2760 6588 2766 6640
rect 2818 6636 2824 6640
rect 3270 6636 3314 6682
rect 3564 6664 3605 6703
rect 4622 6711 4628 6763
rect 4680 6711 4686 6763
rect 5117 6761 5169 6767
rect 3976 6694 4028 6700
rect 2818 6592 3314 6636
rect 3979 6647 4018 6694
rect 4637 6647 4671 6711
rect 5117 6703 5169 6709
rect 5122 6664 5164 6703
rect 5202 6664 5244 7477
rect 5282 6664 5324 7812
rect 5362 6664 5404 7812
rect 5442 6664 5484 7812
rect 5522 6664 5564 7812
rect 6820 7808 6872 7814
rect 6974 7810 7026 7816
rect 5662 7686 6202 7728
rect 5662 7630 5704 7686
rect 5760 7684 5784 7686
rect 5840 7684 5864 7686
rect 5920 7684 5944 7686
rect 6000 7684 6024 7686
rect 6080 7684 6104 7686
rect 5766 7632 5778 7684
rect 5840 7632 5842 7684
rect 6022 7632 6024 7684
rect 6086 7632 6098 7684
rect 5760 7630 5784 7632
rect 5840 7630 5864 7632
rect 5920 7630 5944 7632
rect 6000 7630 6024 7632
rect 6080 7630 6104 7632
rect 6160 7630 6202 7686
rect 6504 7684 6510 7736
rect 6562 7684 6568 7736
rect 5662 7588 6202 7630
rect 6518 7520 6556 7684
rect 7101 7396 7107 7448
rect 7159 7396 7165 7448
rect 6868 7246 6920 7252
rect 7119 7240 7147 7396
rect 6920 7201 7147 7240
rect 5682 7148 6222 7190
rect 6868 7188 6920 7194
rect 5682 7092 5724 7148
rect 5780 7146 5804 7148
rect 5860 7146 5884 7148
rect 5940 7146 5964 7148
rect 6020 7146 6044 7148
rect 6100 7146 6124 7148
rect 5786 7094 5798 7146
rect 5860 7094 5862 7146
rect 6042 7094 6044 7146
rect 6106 7094 6118 7146
rect 5780 7092 5804 7094
rect 5860 7092 5884 7094
rect 5940 7092 5964 7094
rect 6020 7092 6044 7094
rect 6100 7092 6124 7094
rect 6180 7092 6222 7148
rect 5682 7050 6222 7092
rect 6250 6922 6304 6928
rect 6974 6922 7026 6924
rect 6250 6920 7042 6922
rect 6302 6918 7042 6920
rect 6302 6868 6974 6918
rect 6250 6866 6974 6868
rect 7026 6866 7042 6918
rect 6250 6860 6304 6866
rect 6974 6860 7026 6866
rect 5934 6752 5986 6758
rect 6580 6712 6586 6764
rect 6638 6712 6644 6764
rect 5934 6694 5986 6700
rect 3979 6608 4673 6647
rect 4862 6638 4914 6644
rect 2818 6588 2824 6592
rect 2509 6572 2587 6574
rect 2522 6570 2574 6572
rect 2768 6548 2812 6588
rect 5015 6640 5067 6646
rect 4914 6598 5015 6627
rect 144 5234 212 6402
rect 274 6321 329 6510
rect 372 6474 378 6530
rect 434 6474 440 6530
rect 274 6315 332 6321
rect 274 6261 278 6315
rect 277 6140 332 6261
rect 378 6302 434 6474
rect 1324 6447 1960 6500
rect 1324 6445 1374 6447
rect 1430 6445 1454 6447
rect 1510 6445 1534 6447
rect 1590 6445 1614 6447
rect 1670 6445 1694 6447
rect 1750 6445 1774 6447
rect 1830 6445 1854 6447
rect 1910 6445 1960 6447
rect 1324 6393 1360 6445
rect 1604 6393 1614 6445
rect 1670 6393 1680 6445
rect 1924 6393 1960 6445
rect 1324 6391 1374 6393
rect 1430 6391 1454 6393
rect 1510 6391 1534 6393
rect 1590 6391 1614 6393
rect 1670 6391 1694 6393
rect 1750 6391 1774 6393
rect 1830 6391 1854 6393
rect 1910 6391 1960 6393
rect 1324 6360 1960 6391
rect 3564 6313 3605 6584
rect 4862 6580 4914 6586
rect 5015 6582 5067 6588
rect 5202 6584 5243 6664
rect 5282 6584 5323 6664
rect 5362 6584 5403 6664
rect 5442 6584 5483 6664
rect 5522 6584 5563 6664
rect 5938 6648 5976 6694
rect 6596 6648 6630 6712
rect 5938 6608 6632 6648
rect 6820 6638 6872 6644
rect 6974 6640 7026 6646
rect 6872 6598 6974 6628
rect 3704 6458 4244 6500
rect 3704 6402 3746 6458
rect 3802 6456 3826 6458
rect 3882 6456 3906 6458
rect 3962 6456 3986 6458
rect 4042 6456 4066 6458
rect 4122 6456 4146 6458
rect 3808 6404 3820 6456
rect 3882 6404 3884 6456
rect 4064 6404 4066 6456
rect 4128 6404 4140 6456
rect 3802 6402 3826 6404
rect 3882 6402 3906 6404
rect 3962 6402 3986 6404
rect 4042 6402 4066 6404
rect 4122 6402 4146 6404
rect 4202 6402 4244 6458
rect 4546 6455 4552 6507
rect 4604 6455 4610 6507
rect 3704 6360 4244 6402
rect 3564 6307 3617 6313
rect 274 5515 329 6140
rect 378 5686 433 6302
rect 3564 6255 3565 6307
rect 4559 6291 4598 6455
rect 5122 6313 5164 6584
rect 5117 6307 5169 6313
rect 3564 6249 3617 6255
rect 5117 6249 5169 6255
rect 1348 5921 1880 5962
rect 1348 5865 1388 5921
rect 1444 5919 1468 5921
rect 1524 5919 1548 5921
rect 1604 5919 1628 5921
rect 1684 5919 1708 5921
rect 1764 5919 1788 5921
rect 1450 5867 1462 5919
rect 1524 5867 1526 5919
rect 1706 5867 1708 5919
rect 1770 5867 1782 5919
rect 1444 5865 1468 5867
rect 1524 5865 1548 5867
rect 1604 5865 1628 5867
rect 1684 5865 1708 5867
rect 1764 5865 1788 5867
rect 1844 5865 1880 5921
rect 560 5848 612 5854
rect 700 5846 756 5852
rect 612 5844 976 5846
rect 612 5796 702 5844
rect 560 5792 702 5796
rect 754 5792 976 5844
rect 1348 5822 1880 5865
rect 2759 5804 2827 5812
rect 560 5790 1268 5792
rect 700 5784 756 5790
rect 920 5784 1268 5790
rect 2759 5784 2769 5804
rect 920 5752 2769 5784
rect 2821 5752 2827 5804
rect 920 5740 2827 5752
rect 920 5736 1268 5740
rect 852 5694 904 5700
rect 372 5631 378 5686
rect 433 5631 439 5686
rect 1396 5695 2851 5704
rect 3268 5699 3320 5705
rect 1396 5690 3268 5695
rect 904 5660 3268 5690
rect 904 5646 1440 5660
rect 2851 5651 3268 5660
rect 852 5636 904 5642
rect 3268 5641 3320 5647
rect 1930 5614 1990 5625
rect 1004 5602 1056 5608
rect 1930 5603 1932 5614
rect 1056 5591 1242 5598
rect 1599 5591 1932 5603
rect 1056 5569 1932 5591
rect 1056 5557 1633 5569
rect 1930 5558 1932 5569
rect 1988 5603 1990 5614
rect 1988 5569 1991 5603
rect 1988 5558 1990 5569
rect 1056 5554 1242 5557
rect 1004 5544 1056 5550
rect 1930 5547 1990 5558
rect 3564 5539 3605 6249
rect 5029 6085 5035 6137
rect 5087 6085 5093 6137
rect 4744 6018 4796 6024
rect 5047 6012 5075 6085
rect 4796 5973 5075 6012
rect 3724 5920 4264 5962
rect 4744 5960 4796 5966
rect 3724 5864 3766 5920
rect 3822 5918 3846 5920
rect 3902 5918 3926 5920
rect 3982 5918 4006 5920
rect 4062 5918 4086 5920
rect 4142 5918 4166 5920
rect 3828 5866 3840 5918
rect 3902 5866 3904 5918
rect 4084 5866 4086 5918
rect 4148 5866 4160 5918
rect 3822 5864 3846 5866
rect 3902 5864 3926 5866
rect 3982 5864 4006 5866
rect 4062 5864 4086 5866
rect 4142 5864 4166 5866
rect 4222 5864 4264 5920
rect 3724 5822 4264 5864
rect 4291 5693 4346 5699
rect 5016 5693 5068 5696
rect 4291 5691 5084 5693
rect 4291 5639 4292 5691
rect 4344 5690 5084 5691
rect 4344 5639 5016 5690
rect 4291 5638 5016 5639
rect 5068 5638 5084 5690
rect 4291 5632 4346 5638
rect 5016 5632 5068 5638
rect 3561 5533 3613 5539
rect 1154 5515 1209 5521
rect 274 5513 1209 5515
rect 274 5461 1155 5513
rect 1207 5461 1209 5513
rect 274 5460 1209 5461
rect 1154 5454 1209 5460
rect 1754 5516 1814 5522
rect 2267 5516 2325 5525
rect 1754 5513 2325 5516
rect 2838 5513 2898 5518
rect 1754 5512 2898 5513
rect 1754 5460 1758 5512
rect 1810 5510 2908 5512
rect 1810 5460 2270 5510
rect 1754 5458 2270 5460
rect 2322 5508 2908 5510
rect 2322 5458 2842 5508
rect 1754 5456 2842 5458
rect 2894 5456 2908 5508
rect 1754 5450 1814 5456
rect 2267 5455 2908 5456
rect 2267 5443 2325 5455
rect 2838 5452 2908 5455
rect 3262 5454 3268 5506
rect 3320 5454 3326 5506
rect 3976 5524 4028 5530
rect 3561 5475 3613 5481
rect 3975 5475 3976 5518
rect 2838 5446 2898 5452
rect 2768 5412 2816 5416
rect 378 5401 433 5407
rect 1248 5402 1300 5408
rect 433 5398 619 5401
rect 433 5354 1248 5398
rect 433 5346 619 5354
rect 2020 5402 2072 5408
rect 2522 5404 2574 5406
rect 1300 5354 2020 5398
rect 378 5340 433 5346
rect 1248 5344 1300 5350
rect 2020 5344 2072 5350
rect 2509 5402 2587 5404
rect 2509 5346 2520 5402
rect 2576 5346 2587 5402
rect 2760 5360 2766 5412
rect 2818 5408 2824 5412
rect 3270 5408 3314 5454
rect 3564 5436 3605 5475
rect 4622 5483 4628 5535
rect 4680 5483 4686 5535
rect 3976 5466 4028 5472
rect 2818 5364 3314 5408
rect 3979 5419 4018 5466
rect 4637 5419 4671 5483
rect 5122 5436 5164 6249
rect 5202 5436 5244 6584
rect 5282 5539 5324 6584
rect 5279 5533 5331 5539
rect 5279 5475 5331 5481
rect 5282 5436 5324 5475
rect 5362 5436 5404 6584
rect 5442 5436 5484 6584
rect 5522 5436 5564 6584
rect 6820 6580 6872 6586
rect 6974 6582 7026 6588
rect 5662 6458 6202 6500
rect 5662 6402 5704 6458
rect 5760 6456 5784 6458
rect 5840 6456 5864 6458
rect 5920 6456 5944 6458
rect 6000 6456 6024 6458
rect 6080 6456 6104 6458
rect 5766 6404 5778 6456
rect 5840 6404 5842 6456
rect 6022 6404 6024 6456
rect 6086 6404 6098 6456
rect 5760 6402 5784 6404
rect 5840 6402 5864 6404
rect 5920 6402 5944 6404
rect 6000 6402 6024 6404
rect 6080 6402 6104 6404
rect 6160 6402 6202 6458
rect 6504 6456 6510 6508
rect 6562 6456 6568 6508
rect 5662 6360 6202 6402
rect 6518 6292 6556 6456
rect 6974 6138 7026 6144
rect 7202 6127 7241 8429
rect 7026 6097 7241 6127
rect 6974 6080 7026 6086
rect 5682 5920 6222 5962
rect 5682 5864 5724 5920
rect 5780 5918 5804 5920
rect 5860 5918 5884 5920
rect 5940 5918 5964 5920
rect 6020 5918 6044 5920
rect 6100 5918 6124 5920
rect 5786 5866 5798 5918
rect 5860 5866 5862 5918
rect 6042 5866 6044 5918
rect 6106 5866 6118 5918
rect 5780 5864 5804 5866
rect 5860 5864 5884 5866
rect 5940 5864 5964 5866
rect 6020 5864 6044 5866
rect 6100 5864 6124 5866
rect 6180 5864 6222 5920
rect 5682 5822 6222 5864
rect 6250 5694 6304 5700
rect 6974 5694 7026 5696
rect 6250 5692 7042 5694
rect 6302 5690 7042 5692
rect 6302 5640 6974 5690
rect 6250 5638 6974 5640
rect 7026 5638 7042 5690
rect 6250 5632 6304 5638
rect 6974 5632 7026 5638
rect 5934 5524 5986 5530
rect 6580 5484 6586 5536
rect 6638 5484 6644 5536
rect 5934 5466 5986 5472
rect 3979 5380 4673 5419
rect 4862 5410 4914 5416
rect 2818 5360 2824 5364
rect 2509 5344 2587 5346
rect 2522 5342 2574 5344
rect 2768 5320 2812 5360
rect 5015 5412 5067 5418
rect 4914 5370 5015 5399
rect 144 4014 212 5166
rect 274 5093 329 5282
rect 372 5246 378 5302
rect 434 5246 440 5302
rect 274 5087 332 5093
rect 274 5033 278 5087
rect 277 4912 332 5033
rect 378 5074 434 5246
rect 1324 5219 1960 5272
rect 1324 5217 1374 5219
rect 1430 5217 1454 5219
rect 1510 5217 1534 5219
rect 1590 5217 1614 5219
rect 1670 5217 1694 5219
rect 1750 5217 1774 5219
rect 1830 5217 1854 5219
rect 1910 5217 1960 5219
rect 1324 5165 1360 5217
rect 1604 5165 1614 5217
rect 1670 5165 1680 5217
rect 1924 5165 1960 5217
rect 1324 5163 1374 5165
rect 1430 5163 1454 5165
rect 1510 5163 1534 5165
rect 1590 5163 1614 5165
rect 1670 5163 1694 5165
rect 1750 5163 1774 5165
rect 1830 5163 1854 5165
rect 1910 5163 1960 5165
rect 1324 5132 1960 5163
rect 3564 5085 3605 5356
rect 4862 5352 4914 5358
rect 5015 5354 5067 5360
rect 5122 5356 5163 5436
rect 5202 5356 5243 5436
rect 5362 5356 5403 5436
rect 5442 5356 5483 5436
rect 5522 5356 5563 5436
rect 5938 5420 5976 5466
rect 6596 5420 6630 5484
rect 5938 5380 6632 5420
rect 6820 5410 6872 5416
rect 6974 5412 7026 5418
rect 6872 5370 6974 5400
rect 3704 5230 4244 5272
rect 3704 5174 3746 5230
rect 3802 5228 3826 5230
rect 3882 5228 3906 5230
rect 3962 5228 3986 5230
rect 4042 5228 4066 5230
rect 4122 5228 4146 5230
rect 3808 5176 3820 5228
rect 3882 5176 3884 5228
rect 4064 5176 4066 5228
rect 4128 5176 4140 5228
rect 3802 5174 3826 5176
rect 3882 5174 3906 5176
rect 3962 5174 3986 5176
rect 4042 5174 4066 5176
rect 4122 5174 4146 5176
rect 4202 5174 4244 5230
rect 4546 5227 4552 5279
rect 4604 5227 4610 5279
rect 3704 5132 4244 5174
rect 3564 5079 3617 5085
rect 274 4287 329 4912
rect 378 4458 433 5074
rect 3564 5027 3565 5079
rect 4559 5063 4598 5227
rect 3564 5021 3617 5027
rect 1348 4693 1880 4734
rect 1348 4637 1388 4693
rect 1444 4691 1468 4693
rect 1524 4691 1548 4693
rect 1604 4691 1628 4693
rect 1684 4691 1708 4693
rect 1764 4691 1788 4693
rect 1450 4639 1462 4691
rect 1524 4639 1526 4691
rect 1706 4639 1708 4691
rect 1770 4639 1782 4691
rect 1444 4637 1468 4639
rect 1524 4637 1548 4639
rect 1604 4637 1628 4639
rect 1684 4637 1708 4639
rect 1764 4637 1788 4639
rect 1844 4637 1880 4693
rect 560 4620 612 4626
rect 700 4618 756 4624
rect 612 4616 976 4618
rect 612 4568 702 4616
rect 560 4564 702 4568
rect 754 4564 976 4616
rect 1348 4594 1880 4637
rect 2759 4576 2827 4584
rect 560 4562 1268 4564
rect 700 4556 756 4562
rect 920 4556 1268 4562
rect 2759 4556 2769 4576
rect 920 4524 2769 4556
rect 2821 4524 2827 4576
rect 920 4512 2827 4524
rect 920 4508 1268 4512
rect 852 4466 904 4472
rect 372 4403 378 4458
rect 433 4403 439 4458
rect 1396 4467 2851 4476
rect 3268 4471 3320 4477
rect 1396 4462 3268 4467
rect 904 4432 3268 4462
rect 904 4418 1440 4432
rect 2851 4423 3268 4432
rect 852 4408 904 4414
rect 3268 4413 3320 4419
rect 1930 4386 1990 4397
rect 1004 4374 1056 4380
rect 1930 4375 1932 4386
rect 1056 4363 1242 4370
rect 1599 4363 1932 4375
rect 1056 4341 1932 4363
rect 1056 4329 1633 4341
rect 1930 4330 1932 4341
rect 1988 4375 1990 4386
rect 1988 4341 1991 4375
rect 1988 4330 1990 4341
rect 1056 4326 1242 4329
rect 1004 4316 1056 4322
rect 1930 4319 1990 4330
rect 3564 4311 3605 5021
rect 5023 4820 5029 4872
rect 5081 4820 5087 4872
rect 4744 4790 4796 4796
rect 5036 4784 5075 4820
rect 4796 4745 5075 4784
rect 3724 4692 4264 4734
rect 4744 4732 4796 4738
rect 3724 4636 3766 4692
rect 3822 4690 3846 4692
rect 3902 4690 3926 4692
rect 3982 4690 4006 4692
rect 4062 4690 4086 4692
rect 4142 4690 4166 4692
rect 3828 4638 3840 4690
rect 3902 4638 3904 4690
rect 4084 4638 4086 4690
rect 4148 4638 4160 4690
rect 3822 4636 3846 4638
rect 3902 4636 3926 4638
rect 3982 4636 4006 4638
rect 4062 4636 4086 4638
rect 4142 4636 4166 4638
rect 4222 4636 4264 4692
rect 3724 4594 4264 4636
rect 4291 4465 4346 4471
rect 5016 4465 5068 4468
rect 4291 4463 5084 4465
rect 4291 4411 4292 4463
rect 4344 4462 5084 4463
rect 4344 4411 5016 4462
rect 4291 4410 5016 4411
rect 5068 4410 5084 4462
rect 4291 4404 4346 4410
rect 5016 4404 5068 4410
rect 5122 4311 5164 5356
rect 3561 4305 3613 4311
rect 1154 4287 1209 4293
rect 274 4285 1209 4287
rect 274 4233 1155 4285
rect 1207 4233 1209 4285
rect 274 4232 1209 4233
rect 1154 4226 1209 4232
rect 1754 4288 1814 4294
rect 2267 4288 2325 4297
rect 1754 4285 2325 4288
rect 2838 4285 2898 4290
rect 1754 4284 2898 4285
rect 1754 4232 1758 4284
rect 1810 4282 2908 4284
rect 1810 4232 2270 4282
rect 1754 4230 2270 4232
rect 2322 4280 2908 4282
rect 2322 4230 2842 4280
rect 1754 4228 2842 4230
rect 2894 4228 2908 4280
rect 1754 4222 1814 4228
rect 2267 4227 2908 4228
rect 2267 4215 2325 4227
rect 2838 4224 2908 4227
rect 3262 4226 3268 4278
rect 3320 4226 3326 4278
rect 3976 4296 4028 4302
rect 3561 4247 3613 4253
rect 3975 4247 3976 4290
rect 2838 4218 2898 4224
rect 2768 4184 2816 4188
rect 378 4173 433 4179
rect 1248 4174 1300 4180
rect 433 4170 619 4173
rect 433 4126 1248 4170
rect 433 4118 619 4126
rect 2020 4174 2072 4180
rect 2522 4176 2574 4178
rect 1300 4126 2020 4170
rect 378 4112 433 4118
rect 1248 4116 1300 4122
rect 2020 4116 2072 4122
rect 2509 4174 2587 4176
rect 2509 4118 2520 4174
rect 2576 4118 2587 4174
rect 2760 4132 2766 4184
rect 2818 4180 2824 4184
rect 3270 4180 3314 4226
rect 3564 4208 3605 4247
rect 4622 4255 4628 4307
rect 4680 4255 4686 4307
rect 5117 4305 5169 4311
rect 3976 4238 4028 4244
rect 2818 4136 3314 4180
rect 3979 4191 4018 4238
rect 4637 4191 4671 4255
rect 5117 4247 5169 4253
rect 5122 4208 5164 4247
rect 5202 4208 5244 5356
rect 5282 5085 5324 5356
rect 5279 5079 5331 5085
rect 5279 5021 5331 5027
rect 5282 4208 5324 5021
rect 5362 4208 5404 5356
rect 5442 4208 5484 5356
rect 5522 4208 5564 5356
rect 6820 5352 6872 5358
rect 6974 5354 7026 5360
rect 5662 5230 6202 5272
rect 5662 5174 5704 5230
rect 5760 5228 5784 5230
rect 5840 5228 5864 5230
rect 5920 5228 5944 5230
rect 6000 5228 6024 5230
rect 6080 5228 6104 5230
rect 5766 5176 5778 5228
rect 5840 5176 5842 5228
rect 6022 5176 6024 5228
rect 6086 5176 6098 5228
rect 5760 5174 5784 5176
rect 5840 5174 5864 5176
rect 5920 5174 5944 5176
rect 6000 5174 6024 5176
rect 6080 5174 6104 5176
rect 6160 5174 6202 5230
rect 6504 5228 6510 5280
rect 6562 5228 6568 5280
rect 5662 5132 6202 5174
rect 6518 5102 6556 5228
rect 7283 5102 7322 9970
rect 6517 5063 7322 5102
rect 6868 4790 6920 4796
rect 6920 4745 7147 4784
rect 5682 4692 6222 4734
rect 6868 4732 6920 4738
rect 5682 4636 5724 4692
rect 5780 4690 5804 4692
rect 5860 4690 5884 4692
rect 5940 4690 5964 4692
rect 6020 4690 6044 4692
rect 6100 4690 6124 4692
rect 5786 4638 5798 4690
rect 5860 4638 5862 4690
rect 6042 4638 6044 4690
rect 6106 4638 6118 4690
rect 5780 4636 5804 4638
rect 5860 4636 5884 4638
rect 5940 4636 5964 4638
rect 6020 4636 6044 4638
rect 6100 4636 6124 4638
rect 6180 4636 6222 4692
rect 5682 4594 6222 4636
rect 7188 4620 7194 4672
rect 7246 4620 7252 4672
rect 6250 4466 6304 4472
rect 6974 4466 7026 4468
rect 6250 4464 7042 4466
rect 6302 4462 7042 4464
rect 6302 4412 6974 4462
rect 6250 4410 6974 4412
rect 7026 4410 7042 4462
rect 6250 4404 6304 4410
rect 6974 4404 7026 4410
rect 5934 4296 5986 4302
rect 6580 4256 6586 4308
rect 6638 4256 6644 4308
rect 5934 4238 5986 4244
rect 3979 4152 4673 4191
rect 4862 4182 4914 4188
rect 2818 4132 2824 4136
rect 2509 4116 2587 4118
rect 2522 4114 2574 4116
rect 2768 4092 2812 4132
rect 5015 4184 5067 4190
rect 4914 4142 5015 4171
rect 144 2778 212 3946
rect 274 3865 329 4054
rect 372 4018 378 4074
rect 434 4018 440 4074
rect 274 3859 332 3865
rect 274 3805 278 3859
rect 277 3684 332 3805
rect 378 3846 434 4018
rect 1324 3991 1960 4044
rect 1324 3989 1374 3991
rect 1430 3989 1454 3991
rect 1510 3989 1534 3991
rect 1590 3989 1614 3991
rect 1670 3989 1694 3991
rect 1750 3989 1774 3991
rect 1830 3989 1854 3991
rect 1910 3989 1960 3991
rect 1324 3937 1360 3989
rect 1604 3937 1614 3989
rect 1670 3937 1680 3989
rect 1924 3937 1960 3989
rect 1324 3935 1374 3937
rect 1430 3935 1454 3937
rect 1510 3935 1534 3937
rect 1590 3935 1614 3937
rect 1670 3935 1694 3937
rect 1750 3935 1774 3937
rect 1830 3935 1854 3937
rect 1910 3935 1960 3937
rect 1324 3904 1960 3935
rect 3564 3857 3605 4128
rect 4862 4124 4914 4130
rect 5015 4126 5067 4132
rect 5202 4128 5243 4208
rect 5282 4128 5323 4208
rect 5362 4128 5403 4208
rect 5442 4128 5483 4208
rect 5522 4128 5563 4208
rect 5938 4192 5976 4238
rect 6596 4192 6630 4256
rect 5938 4152 6632 4192
rect 6820 4182 6872 4188
rect 6974 4184 7026 4190
rect 6872 4142 6974 4172
rect 3704 4002 4244 4044
rect 3704 3946 3746 4002
rect 3802 4000 3826 4002
rect 3882 4000 3906 4002
rect 3962 4000 3986 4002
rect 4042 4000 4066 4002
rect 4122 4000 4146 4002
rect 3808 3948 3820 4000
rect 3882 3948 3884 4000
rect 4064 3948 4066 4000
rect 4128 3948 4140 4000
rect 3802 3946 3826 3948
rect 3882 3946 3906 3948
rect 3962 3946 3986 3948
rect 4042 3946 4066 3948
rect 4122 3946 4146 3948
rect 4202 3946 4244 4002
rect 4546 3999 4552 4051
rect 4604 3999 4610 4051
rect 3704 3904 4244 3946
rect 3564 3851 3617 3857
rect 274 3059 329 3684
rect 378 3230 433 3846
rect 3564 3799 3565 3851
rect 4559 3835 4598 3999
rect 5122 3857 5164 4128
rect 5117 3851 5169 3857
rect 3564 3793 3617 3799
rect 5117 3793 5169 3799
rect 1348 3465 1880 3506
rect 1348 3409 1388 3465
rect 1444 3463 1468 3465
rect 1524 3463 1548 3465
rect 1604 3463 1628 3465
rect 1684 3463 1708 3465
rect 1764 3463 1788 3465
rect 1450 3411 1462 3463
rect 1524 3411 1526 3463
rect 1706 3411 1708 3463
rect 1770 3411 1782 3463
rect 1444 3409 1468 3411
rect 1524 3409 1548 3411
rect 1604 3409 1628 3411
rect 1684 3409 1708 3411
rect 1764 3409 1788 3411
rect 1844 3409 1880 3465
rect 560 3392 612 3398
rect 700 3390 756 3396
rect 612 3388 976 3390
rect 612 3340 702 3388
rect 560 3336 702 3340
rect 754 3336 976 3388
rect 1348 3366 1880 3409
rect 2759 3348 2827 3356
rect 560 3334 1268 3336
rect 700 3328 756 3334
rect 920 3328 1268 3334
rect 2759 3328 2769 3348
rect 920 3296 2769 3328
rect 2821 3296 2827 3348
rect 920 3284 2827 3296
rect 920 3280 1268 3284
rect 852 3238 904 3244
rect 372 3175 378 3230
rect 433 3175 439 3230
rect 1396 3239 2851 3248
rect 3268 3243 3320 3249
rect 1396 3234 3268 3239
rect 904 3204 3268 3234
rect 904 3190 1440 3204
rect 2851 3195 3268 3204
rect 852 3180 904 3186
rect 3268 3185 3320 3191
rect 1930 3158 1990 3169
rect 1004 3146 1056 3152
rect 1930 3147 1932 3158
rect 1056 3135 1242 3142
rect 1599 3135 1932 3147
rect 1056 3113 1932 3135
rect 1056 3101 1633 3113
rect 1930 3102 1932 3113
rect 1988 3147 1990 3158
rect 1988 3113 1991 3147
rect 1988 3102 1990 3113
rect 1056 3098 1242 3101
rect 1004 3088 1056 3094
rect 1930 3091 1990 3102
rect 3564 3083 3605 3793
rect 5029 3629 5035 3681
rect 5087 3629 5093 3681
rect 4744 3562 4796 3568
rect 5047 3556 5075 3629
rect 4796 3517 5075 3556
rect 3724 3464 4264 3506
rect 4744 3504 4796 3510
rect 3724 3408 3766 3464
rect 3822 3462 3846 3464
rect 3902 3462 3926 3464
rect 3982 3462 4006 3464
rect 4062 3462 4086 3464
rect 4142 3462 4166 3464
rect 3828 3410 3840 3462
rect 3902 3410 3904 3462
rect 4084 3410 4086 3462
rect 4148 3410 4160 3462
rect 3822 3408 3846 3410
rect 3902 3408 3926 3410
rect 3982 3408 4006 3410
rect 4062 3408 4086 3410
rect 4142 3408 4166 3410
rect 4222 3408 4264 3464
rect 3724 3366 4264 3408
rect 4291 3237 4346 3243
rect 5016 3237 5068 3240
rect 4291 3235 5084 3237
rect 4291 3183 4292 3235
rect 4344 3234 5084 3235
rect 4344 3183 5016 3234
rect 4291 3182 5016 3183
rect 5068 3182 5084 3234
rect 4291 3176 4346 3182
rect 5016 3176 5068 3182
rect 3561 3077 3613 3083
rect 1154 3059 1209 3065
rect 274 3057 1209 3059
rect 274 3005 1155 3057
rect 1207 3005 1209 3057
rect 274 3004 1209 3005
rect 1154 2998 1209 3004
rect 1754 3060 1814 3066
rect 2267 3060 2325 3069
rect 1754 3057 2325 3060
rect 2838 3057 2898 3062
rect 1754 3056 2898 3057
rect 1754 3004 1758 3056
rect 1810 3054 2908 3056
rect 1810 3004 2270 3054
rect 1754 3002 2270 3004
rect 2322 3052 2908 3054
rect 2322 3002 2842 3052
rect 1754 3000 2842 3002
rect 2894 3000 2908 3052
rect 1754 2994 1814 3000
rect 2267 2999 2908 3000
rect 2267 2987 2325 2999
rect 2838 2996 2908 2999
rect 3262 2998 3268 3050
rect 3320 2998 3326 3050
rect 3976 3068 4028 3074
rect 3561 3019 3613 3025
rect 3975 3019 3976 3062
rect 2838 2990 2898 2996
rect 2768 2956 2816 2960
rect 378 2945 433 2951
rect 1248 2946 1300 2952
rect 433 2942 619 2945
rect 433 2898 1248 2942
rect 433 2890 619 2898
rect 2020 2946 2072 2952
rect 2522 2948 2574 2950
rect 1300 2898 2020 2942
rect 378 2884 433 2890
rect 1248 2888 1300 2894
rect 2020 2888 2072 2894
rect 2509 2946 2587 2948
rect 2509 2890 2520 2946
rect 2576 2890 2587 2946
rect 2760 2904 2766 2956
rect 2818 2952 2824 2956
rect 3270 2952 3314 2998
rect 3564 2980 3605 3019
rect 4622 3027 4628 3079
rect 4680 3027 4686 3079
rect 3976 3010 4028 3016
rect 2818 2908 3314 2952
rect 3979 2963 4018 3010
rect 4637 2963 4671 3027
rect 5122 2980 5164 3793
rect 5202 3083 5244 4128
rect 5197 3077 5249 3083
rect 5197 3019 5249 3025
rect 5202 2980 5244 3019
rect 5282 2980 5324 4128
rect 5362 2980 5404 4128
rect 5442 2980 5484 4128
rect 5522 2980 5564 4128
rect 6820 4124 6872 4130
rect 6974 4126 7026 4132
rect 5662 4002 6202 4044
rect 5662 3946 5704 4002
rect 5760 4000 5784 4002
rect 5840 4000 5864 4002
rect 5920 4000 5944 4002
rect 6000 4000 6024 4002
rect 6080 4000 6104 4002
rect 5766 3948 5778 4000
rect 5840 3948 5842 4000
rect 6022 3948 6024 4000
rect 6086 3948 6098 4000
rect 5760 3946 5784 3948
rect 5840 3946 5864 3948
rect 5920 3946 5944 3948
rect 6000 3946 6024 3948
rect 6080 3946 6104 3948
rect 6160 3946 6202 4002
rect 6504 4000 6510 4052
rect 6562 4000 6568 4052
rect 5662 3904 6202 3946
rect 6518 3836 6556 4000
rect 6523 3766 6553 3836
rect 6506 3714 6512 3766
rect 6564 3714 6570 3766
rect 6843 3562 6895 3568
rect 7196 3556 7235 4620
rect 6895 3517 7235 3556
rect 5682 3464 6222 3506
rect 6843 3504 6895 3510
rect 5682 3408 5724 3464
rect 5780 3462 5804 3464
rect 5860 3462 5884 3464
rect 5940 3462 5964 3464
rect 6020 3462 6044 3464
rect 6100 3462 6124 3464
rect 5786 3410 5798 3462
rect 5860 3410 5862 3462
rect 6042 3410 6044 3462
rect 6106 3410 6118 3462
rect 5780 3408 5804 3410
rect 5860 3408 5884 3410
rect 5940 3408 5964 3410
rect 6020 3408 6044 3410
rect 6100 3408 6124 3410
rect 6180 3408 6222 3464
rect 5682 3366 6222 3408
rect 6250 3238 6304 3244
rect 6974 3238 7026 3240
rect 6250 3236 7042 3238
rect 6302 3234 7042 3236
rect 6302 3184 6974 3234
rect 6250 3182 6974 3184
rect 7026 3182 7042 3234
rect 6250 3176 6304 3182
rect 6974 3176 7026 3182
rect 5934 3068 5986 3074
rect 6580 3028 6586 3080
rect 6638 3028 6644 3080
rect 5934 3010 5986 3016
rect 3979 2924 4673 2963
rect 4862 2954 4914 2960
rect 2818 2904 2824 2908
rect 2509 2888 2587 2890
rect 2522 2886 2574 2888
rect 2768 2864 2812 2904
rect 5015 2956 5067 2962
rect 4914 2914 5015 2943
rect 144 1558 212 2710
rect 274 2637 329 2826
rect 372 2790 378 2846
rect 434 2790 440 2846
rect 274 2631 332 2637
rect 274 2577 278 2631
rect 277 2456 332 2577
rect 378 2618 434 2790
rect 1324 2763 1960 2816
rect 1324 2761 1374 2763
rect 1430 2761 1454 2763
rect 1510 2761 1534 2763
rect 1590 2761 1614 2763
rect 1670 2761 1694 2763
rect 1750 2761 1774 2763
rect 1830 2761 1854 2763
rect 1910 2761 1960 2763
rect 1324 2709 1360 2761
rect 1604 2709 1614 2761
rect 1670 2709 1680 2761
rect 1924 2709 1960 2761
rect 1324 2707 1374 2709
rect 1430 2707 1454 2709
rect 1510 2707 1534 2709
rect 1590 2707 1614 2709
rect 1670 2707 1694 2709
rect 1750 2707 1774 2709
rect 1830 2707 1854 2709
rect 1910 2707 1960 2709
rect 1324 2676 1960 2707
rect 3564 2629 3605 2900
rect 4862 2896 4914 2902
rect 5015 2898 5067 2904
rect 5122 2900 5163 2980
rect 5282 2900 5323 2980
rect 5362 2900 5403 2980
rect 5442 2900 5483 2980
rect 5522 2900 5563 2980
rect 5938 2964 5976 3010
rect 6596 2964 6630 3028
rect 5938 2924 6632 2964
rect 6820 2954 6872 2960
rect 6974 2956 7026 2962
rect 6872 2914 6974 2944
rect 3704 2774 4244 2816
rect 3704 2718 3746 2774
rect 3802 2772 3826 2774
rect 3882 2772 3906 2774
rect 3962 2772 3986 2774
rect 4042 2772 4066 2774
rect 4122 2772 4146 2774
rect 3808 2720 3820 2772
rect 3882 2720 3884 2772
rect 4064 2720 4066 2772
rect 4128 2720 4140 2772
rect 3802 2718 3826 2720
rect 3882 2718 3906 2720
rect 3962 2718 3986 2720
rect 4042 2718 4066 2720
rect 4122 2718 4146 2720
rect 4202 2718 4244 2774
rect 4546 2771 4552 2823
rect 4604 2771 4610 2823
rect 3704 2676 4244 2718
rect 3564 2623 3617 2629
rect 274 1831 329 2456
rect 378 2002 433 2618
rect 3564 2571 3565 2623
rect 4559 2607 4598 2771
rect 3564 2565 3617 2571
rect 1348 2237 1880 2278
rect 1348 2181 1388 2237
rect 1444 2235 1468 2237
rect 1524 2235 1548 2237
rect 1604 2235 1628 2237
rect 1684 2235 1708 2237
rect 1764 2235 1788 2237
rect 1450 2183 1462 2235
rect 1524 2183 1526 2235
rect 1706 2183 1708 2235
rect 1770 2183 1782 2235
rect 1444 2181 1468 2183
rect 1524 2181 1548 2183
rect 1604 2181 1628 2183
rect 1684 2181 1708 2183
rect 1764 2181 1788 2183
rect 1844 2181 1880 2237
rect 560 2164 612 2170
rect 700 2162 756 2168
rect 612 2160 976 2162
rect 612 2112 702 2160
rect 560 2108 702 2112
rect 754 2108 976 2160
rect 1348 2138 1880 2181
rect 2759 2120 2827 2128
rect 560 2106 1268 2108
rect 700 2100 756 2106
rect 920 2100 1268 2106
rect 2759 2100 2769 2120
rect 920 2068 2769 2100
rect 2821 2068 2827 2120
rect 920 2056 2827 2068
rect 920 2052 1268 2056
rect 852 2010 904 2016
rect 372 1947 378 2002
rect 433 1947 439 2002
rect 1396 2011 2851 2020
rect 3268 2015 3320 2021
rect 1396 2006 3268 2011
rect 904 1976 3268 2006
rect 904 1962 1440 1976
rect 2851 1967 3268 1976
rect 852 1952 904 1958
rect 3268 1957 3320 1963
rect 1930 1930 1990 1941
rect 1004 1918 1056 1924
rect 1930 1919 1932 1930
rect 1056 1907 1242 1914
rect 1599 1907 1932 1919
rect 1056 1885 1932 1907
rect 1056 1873 1633 1885
rect 1930 1874 1932 1885
rect 1988 1919 1990 1930
rect 1988 1885 1991 1919
rect 1988 1874 1990 1885
rect 1056 1870 1242 1873
rect 1004 1860 1056 1866
rect 1930 1863 1990 1874
rect 3564 1855 3605 2565
rect 5023 2364 5029 2416
rect 5081 2364 5087 2416
rect 4744 2334 4796 2340
rect 5036 2328 5075 2364
rect 4796 2289 5075 2328
rect 3724 2236 4264 2278
rect 4744 2276 4796 2282
rect 3724 2180 3766 2236
rect 3822 2234 3846 2236
rect 3902 2234 3926 2236
rect 3982 2234 4006 2236
rect 4062 2234 4086 2236
rect 4142 2234 4166 2236
rect 3828 2182 3840 2234
rect 3902 2182 3904 2234
rect 4084 2182 4086 2234
rect 4148 2182 4160 2234
rect 3822 2180 3846 2182
rect 3902 2180 3926 2182
rect 3982 2180 4006 2182
rect 4062 2180 4086 2182
rect 4142 2180 4166 2182
rect 4222 2180 4264 2236
rect 3724 2138 4264 2180
rect 4291 2009 4346 2015
rect 5016 2009 5068 2012
rect 4291 2007 5084 2009
rect 4291 1955 4292 2007
rect 4344 2006 5084 2007
rect 4344 1955 5016 2006
rect 4291 1954 5016 1955
rect 5068 1954 5084 2006
rect 4291 1948 4346 1954
rect 5016 1948 5068 1954
rect 5122 1855 5164 2900
rect 5202 2629 5244 2900
rect 5197 2623 5249 2629
rect 5197 2565 5249 2571
rect 3561 1849 3613 1855
rect 1154 1831 1209 1837
rect 274 1829 1209 1831
rect 274 1777 1155 1829
rect 1207 1777 1209 1829
rect 274 1776 1209 1777
rect 1154 1770 1209 1776
rect 1754 1832 1814 1838
rect 2267 1832 2325 1841
rect 1754 1829 2325 1832
rect 2838 1829 2898 1834
rect 1754 1828 2898 1829
rect 1754 1776 1758 1828
rect 1810 1826 2908 1828
rect 1810 1776 2270 1826
rect 1754 1774 2270 1776
rect 2322 1824 2908 1826
rect 2322 1774 2842 1824
rect 1754 1772 2842 1774
rect 2894 1772 2908 1824
rect 1754 1766 1814 1772
rect 2267 1771 2908 1772
rect 2267 1759 2325 1771
rect 2838 1768 2908 1771
rect 3262 1770 3268 1822
rect 3320 1770 3326 1822
rect 3976 1840 4028 1846
rect 3561 1791 3613 1797
rect 3975 1791 3976 1834
rect 2838 1762 2898 1768
rect 2768 1728 2816 1732
rect 378 1717 433 1723
rect 1248 1718 1300 1724
rect 433 1714 619 1717
rect 433 1670 1248 1714
rect 433 1662 619 1670
rect 2020 1718 2072 1724
rect 2522 1720 2574 1722
rect 1300 1670 2020 1714
rect 378 1656 433 1662
rect 1248 1660 1300 1666
rect 2020 1660 2072 1666
rect 2509 1718 2587 1720
rect 2509 1662 2520 1718
rect 2576 1662 2587 1718
rect 2760 1676 2766 1728
rect 2818 1724 2824 1728
rect 3270 1724 3314 1770
rect 3564 1752 3605 1791
rect 4622 1799 4628 1851
rect 4680 1799 4686 1851
rect 5117 1849 5169 1855
rect 3976 1782 4028 1788
rect 2818 1680 3314 1724
rect 3979 1735 4018 1782
rect 4637 1735 4671 1799
rect 5117 1791 5169 1797
rect 5122 1752 5164 1791
rect 5202 1752 5244 2565
rect 5282 1752 5324 2900
rect 5362 1752 5404 2900
rect 5442 1752 5484 2900
rect 5522 1752 5564 2900
rect 6820 2896 6872 2902
rect 6974 2898 7026 2904
rect 5662 2774 6202 2816
rect 5662 2718 5704 2774
rect 5760 2772 5784 2774
rect 5840 2772 5864 2774
rect 5920 2772 5944 2774
rect 6000 2772 6024 2774
rect 6080 2772 6104 2774
rect 5766 2720 5778 2772
rect 5840 2720 5842 2772
rect 6022 2720 6024 2772
rect 6086 2720 6098 2772
rect 5760 2718 5784 2720
rect 5840 2718 5864 2720
rect 5920 2718 5944 2720
rect 6000 2718 6024 2720
rect 6080 2718 6104 2720
rect 6160 2718 6202 2774
rect 6504 2772 6510 2824
rect 6562 2772 6568 2824
rect 5662 2676 6202 2718
rect 6518 2608 6556 2772
rect 7101 2484 7107 2536
rect 7159 2484 7165 2536
rect 6868 2334 6920 2340
rect 7119 2328 7147 2484
rect 6920 2289 7147 2328
rect 5682 2236 6222 2278
rect 6868 2276 6920 2282
rect 5682 2180 5724 2236
rect 5780 2234 5804 2236
rect 5860 2234 5884 2236
rect 5940 2234 5964 2236
rect 6020 2234 6044 2236
rect 6100 2234 6124 2236
rect 5786 2182 5798 2234
rect 5860 2182 5862 2234
rect 6042 2182 6044 2234
rect 6106 2182 6118 2234
rect 5780 2180 5804 2182
rect 5860 2180 5884 2182
rect 5940 2180 5964 2182
rect 6020 2180 6044 2182
rect 6100 2180 6124 2182
rect 6180 2180 6222 2236
rect 5682 2138 6222 2180
rect 6250 2010 6304 2016
rect 6974 2010 7026 2012
rect 6250 2008 7042 2010
rect 6302 2006 7042 2008
rect 6302 1956 6974 2006
rect 6250 1954 6974 1956
rect 7026 1954 7042 2006
rect 6250 1948 6304 1954
rect 6974 1948 7026 1954
rect 5934 1840 5986 1846
rect 6580 1800 6586 1852
rect 6638 1800 6644 1852
rect 5934 1782 5986 1788
rect 3979 1696 4673 1735
rect 4862 1726 4914 1732
rect 2818 1676 2824 1680
rect 2509 1660 2587 1662
rect 2522 1658 2574 1660
rect 2768 1636 2812 1676
rect 5015 1728 5067 1734
rect 4914 1686 5015 1715
rect 144 322 212 1490
rect 274 1409 329 1598
rect 372 1562 378 1618
rect 434 1562 440 1618
rect 274 1403 332 1409
rect 274 1349 278 1403
rect 277 1228 332 1349
rect 378 1390 434 1562
rect 1324 1535 1960 1588
rect 1324 1533 1374 1535
rect 1430 1533 1454 1535
rect 1510 1533 1534 1535
rect 1590 1533 1614 1535
rect 1670 1533 1694 1535
rect 1750 1533 1774 1535
rect 1830 1533 1854 1535
rect 1910 1533 1960 1535
rect 1324 1481 1360 1533
rect 1604 1481 1614 1533
rect 1670 1481 1680 1533
rect 1924 1481 1960 1533
rect 1324 1479 1374 1481
rect 1430 1479 1454 1481
rect 1510 1479 1534 1481
rect 1590 1479 1614 1481
rect 1670 1479 1694 1481
rect 1750 1479 1774 1481
rect 1830 1479 1854 1481
rect 1910 1479 1960 1481
rect 1324 1448 1960 1479
rect 3564 1401 3605 1672
rect 4862 1668 4914 1674
rect 5015 1670 5067 1676
rect 5202 1672 5243 1752
rect 5282 1672 5323 1752
rect 5362 1672 5403 1752
rect 5442 1672 5483 1752
rect 5522 1672 5563 1752
rect 5938 1736 5976 1782
rect 6596 1736 6630 1800
rect 5938 1696 6632 1736
rect 6820 1726 6872 1732
rect 6974 1728 7026 1734
rect 6872 1686 6974 1716
rect 3704 1546 4244 1588
rect 3704 1490 3746 1546
rect 3802 1544 3826 1546
rect 3882 1544 3906 1546
rect 3962 1544 3986 1546
rect 4042 1544 4066 1546
rect 4122 1544 4146 1546
rect 3808 1492 3820 1544
rect 3882 1492 3884 1544
rect 4064 1492 4066 1544
rect 4128 1492 4140 1544
rect 3802 1490 3826 1492
rect 3882 1490 3906 1492
rect 3962 1490 3986 1492
rect 4042 1490 4066 1492
rect 4122 1490 4146 1492
rect 4202 1490 4244 1546
rect 4546 1543 4552 1595
rect 4604 1543 4610 1595
rect 3704 1448 4244 1490
rect 3564 1395 3617 1401
rect 274 603 329 1228
rect 378 774 433 1390
rect 3564 1343 3565 1395
rect 4559 1379 4598 1543
rect 5122 1401 5164 1672
rect 5117 1395 5169 1401
rect 3564 1337 3617 1343
rect 5117 1337 5169 1343
rect 1348 1009 1880 1050
rect 1348 953 1388 1009
rect 1444 1007 1468 1009
rect 1524 1007 1548 1009
rect 1604 1007 1628 1009
rect 1684 1007 1708 1009
rect 1764 1007 1788 1009
rect 1450 955 1462 1007
rect 1524 955 1526 1007
rect 1706 955 1708 1007
rect 1770 955 1782 1007
rect 1444 953 1468 955
rect 1524 953 1548 955
rect 1604 953 1628 955
rect 1684 953 1708 955
rect 1764 953 1788 955
rect 1844 953 1880 1009
rect 560 936 612 942
rect 700 934 756 940
rect 612 932 976 934
rect 612 884 702 932
rect 560 880 702 884
rect 754 880 976 932
rect 1348 910 1880 953
rect 2759 892 2827 900
rect 560 878 1268 880
rect 700 872 756 878
rect 920 872 1268 878
rect 2759 872 2769 892
rect 920 840 2769 872
rect 2821 840 2827 892
rect 920 828 2827 840
rect 920 824 1268 828
rect 852 782 904 788
rect 372 719 378 774
rect 433 719 439 774
rect 1396 783 2851 792
rect 3268 787 3320 793
rect 1396 778 3268 783
rect 904 748 3268 778
rect 904 734 1440 748
rect 2851 739 3268 748
rect 852 724 904 730
rect 3268 729 3320 735
rect 1930 702 1990 713
rect 1004 690 1056 696
rect 1930 691 1932 702
rect 1056 679 1242 686
rect 1599 679 1932 691
rect 1056 657 1932 679
rect 1056 645 1633 657
rect 1930 646 1932 657
rect 1988 691 1990 702
rect 1988 657 1991 691
rect 1988 646 1990 657
rect 1056 642 1242 645
rect 1004 632 1056 638
rect 1930 635 1990 646
rect 3564 627 3605 1337
rect 5029 1173 5035 1225
rect 5087 1173 5093 1225
rect 4744 1106 4796 1112
rect 5047 1100 5075 1173
rect 5122 1142 5164 1337
rect 5202 1142 5244 1672
rect 5282 1142 5324 1672
rect 5362 1142 5404 1672
rect 5442 1142 5484 1672
rect 5522 1142 5564 1672
rect 6820 1668 6872 1674
rect 6974 1670 7026 1676
rect 5662 1546 6202 1588
rect 5662 1490 5704 1546
rect 5760 1544 5784 1546
rect 5840 1544 5864 1546
rect 5920 1544 5944 1546
rect 6000 1544 6024 1546
rect 6080 1544 6104 1546
rect 5766 1492 5778 1544
rect 5840 1492 5842 1544
rect 6022 1492 6024 1544
rect 6086 1492 6098 1544
rect 5760 1490 5784 1492
rect 5840 1490 5864 1492
rect 5920 1490 5944 1492
rect 6000 1490 6024 1492
rect 6080 1490 6104 1492
rect 6160 1490 6202 1546
rect 6504 1544 6510 1596
rect 6562 1544 6568 1596
rect 5662 1448 6202 1490
rect 6518 1380 6556 1544
rect 4796 1061 5075 1100
rect 3724 1008 4264 1050
rect 4744 1048 4796 1054
rect 3724 952 3766 1008
rect 3822 1006 3846 1008
rect 3902 1006 3926 1008
rect 3982 1006 4006 1008
rect 4062 1006 4086 1008
rect 4142 1006 4166 1008
rect 3828 954 3840 1006
rect 3902 954 3904 1006
rect 4084 954 4086 1006
rect 4148 954 4160 1006
rect 3822 952 3846 954
rect 3902 952 3926 954
rect 3982 952 4006 954
rect 4062 952 4086 954
rect 4142 952 4166 954
rect 4222 952 4264 1008
rect 3724 910 4264 952
rect 4291 781 4346 787
rect 5016 781 5068 784
rect 4291 779 5084 781
rect 4291 727 4292 779
rect 4344 778 5084 779
rect 4344 727 5016 778
rect 4291 726 5016 727
rect 5068 726 5084 778
rect 4291 720 4346 726
rect 5016 720 5068 726
rect 3561 621 3613 627
rect 1154 603 1209 609
rect 274 601 1209 603
rect 274 549 1155 601
rect 1207 549 1209 601
rect 274 548 1209 549
rect 1154 542 1209 548
rect 1754 604 1814 610
rect 2267 604 2325 613
rect 1754 601 2325 604
rect 2838 601 2898 606
rect 1754 600 2898 601
rect 1754 548 1758 600
rect 1810 598 2908 600
rect 1810 548 2270 598
rect 1754 546 2270 548
rect 2322 596 2908 598
rect 2322 546 2842 596
rect 1754 544 2842 546
rect 2894 544 2908 596
rect 1754 538 1814 544
rect 2267 543 2908 544
rect 2267 531 2325 543
rect 2838 540 2908 543
rect 3262 542 3268 594
rect 3320 542 3326 594
rect 3976 612 4028 618
rect 3561 563 3613 569
rect 3975 563 3976 606
rect 2838 534 2898 540
rect 2768 500 2816 504
rect 378 489 433 495
rect 1248 490 1300 496
rect 433 486 619 489
rect 433 442 1248 486
rect 433 434 619 442
rect 2020 490 2072 496
rect 2522 492 2574 494
rect 1300 442 2020 486
rect 378 428 433 434
rect 1248 432 1300 438
rect 2020 432 2072 438
rect 2509 490 2587 492
rect 2509 434 2520 490
rect 2576 434 2587 490
rect 2760 448 2766 500
rect 2818 496 2824 500
rect 3270 496 3314 542
rect 3564 524 3605 563
rect 4622 571 4628 623
rect 4680 571 4686 623
rect 3976 554 4028 560
rect 2818 452 3314 496
rect 3979 507 4018 554
rect 4637 507 4671 571
rect 3979 468 4673 507
rect 4862 498 4914 504
rect 2818 448 2824 452
rect 2509 432 2587 434
rect 2522 430 2574 432
rect 2768 408 2812 448
rect 5015 500 5067 506
rect 4914 458 5015 487
rect 144 245 212 254
rect 274 225 329 370
rect 372 334 378 390
rect 434 334 440 390
rect 274 175 332 225
rect 274 121 278 175
rect 277 0 332 121
rect 378 162 434 334
rect 1324 307 1960 360
rect 1324 305 1374 307
rect 1430 305 1454 307
rect 1510 305 1534 307
rect 1590 305 1614 307
rect 1670 305 1694 307
rect 1750 305 1774 307
rect 1830 305 1854 307
rect 1910 305 1960 307
rect 1324 253 1360 305
rect 1604 253 1614 305
rect 1670 253 1680 305
rect 1924 253 1960 305
rect 1324 251 1374 253
rect 1430 251 1454 253
rect 1510 251 1534 253
rect 1590 251 1614 253
rect 1670 251 1694 253
rect 1750 251 1774 253
rect 1830 251 1854 253
rect 1910 251 1960 253
rect 1324 220 1960 251
rect 3564 173 3605 444
rect 4862 440 4914 446
rect 5015 442 5067 448
rect 3704 318 4244 360
rect 3704 262 3746 318
rect 3802 316 3826 318
rect 3882 316 3906 318
rect 3962 316 3986 318
rect 4042 316 4066 318
rect 4122 316 4146 318
rect 3808 264 3820 316
rect 3882 264 3884 316
rect 4064 264 4066 316
rect 4128 264 4140 316
rect 3802 262 3826 264
rect 3882 262 3906 264
rect 3962 262 3986 264
rect 4042 262 4066 264
rect 4122 262 4146 264
rect 4202 262 4244 318
rect 4546 315 4552 367
rect 4604 315 4610 367
rect 3704 220 4244 262
rect 3564 167 3617 173
rect 378 0 433 162
rect 3564 115 3565 167
rect 4559 151 4598 315
rect 3564 109 3617 115
rect 3564 0 3605 109
<< via2 >>
rect 42 19358 110 19426
rect 1388 19427 1444 19429
rect 1468 19427 1524 19429
rect 1548 19427 1604 19429
rect 1628 19427 1684 19429
rect 1708 19427 1764 19429
rect 1788 19427 1844 19429
rect 1388 19375 1398 19427
rect 1398 19375 1444 19427
rect 1468 19375 1514 19427
rect 1514 19375 1524 19427
rect 1548 19375 1578 19427
rect 1578 19375 1590 19427
rect 1590 19375 1604 19427
rect 1628 19375 1642 19427
rect 1642 19375 1654 19427
rect 1654 19375 1684 19427
rect 1708 19375 1718 19427
rect 1718 19375 1764 19427
rect 1788 19375 1834 19427
rect 1834 19375 1844 19427
rect 1388 19373 1444 19375
rect 1468 19373 1524 19375
rect 1548 19373 1604 19375
rect 1628 19373 1684 19375
rect 1708 19373 1764 19375
rect 1788 19373 1844 19375
rect 1932 19121 1988 19122
rect 1932 19069 1935 19121
rect 1935 19069 1987 19121
rect 1987 19069 1988 19121
rect 1932 19066 1988 19069
rect 3766 19426 3822 19428
rect 3846 19426 3902 19428
rect 3926 19426 3982 19428
rect 4006 19426 4062 19428
rect 4086 19426 4142 19428
rect 4166 19426 4222 19428
rect 3766 19374 3776 19426
rect 3776 19374 3822 19426
rect 3846 19374 3892 19426
rect 3892 19374 3902 19426
rect 3926 19374 3956 19426
rect 3956 19374 3968 19426
rect 3968 19374 3982 19426
rect 4006 19374 4020 19426
rect 4020 19374 4032 19426
rect 4032 19374 4062 19426
rect 4086 19374 4096 19426
rect 4096 19374 4142 19426
rect 4166 19374 4212 19426
rect 4212 19374 4222 19426
rect 3766 19372 3822 19374
rect 3846 19372 3902 19374
rect 3926 19372 3982 19374
rect 4006 19372 4062 19374
rect 4086 19372 4142 19374
rect 4166 19372 4222 19374
rect 2520 18908 2576 18910
rect 2520 18856 2522 18908
rect 2522 18856 2574 18908
rect 2574 18856 2576 18908
rect 2520 18854 2576 18856
rect 5724 19426 5780 19428
rect 5804 19426 5860 19428
rect 5884 19426 5940 19428
rect 5964 19426 6020 19428
rect 6044 19426 6100 19428
rect 6124 19426 6180 19428
rect 5724 19374 5734 19426
rect 5734 19374 5780 19426
rect 5804 19374 5850 19426
rect 5850 19374 5860 19426
rect 5884 19374 5914 19426
rect 5914 19374 5926 19426
rect 5926 19374 5940 19426
rect 5964 19374 5978 19426
rect 5978 19374 5990 19426
rect 5990 19374 6020 19426
rect 6044 19374 6054 19426
rect 6054 19374 6100 19426
rect 6124 19374 6170 19426
rect 6170 19374 6180 19426
rect 5724 19372 5780 19374
rect 5804 19372 5860 19374
rect 5884 19372 5940 19374
rect 5964 19372 6020 19374
rect 6044 19372 6100 19374
rect 6124 19372 6180 19374
rect 42 18152 110 18220
rect 42 16902 110 16970
rect 42 15696 110 15764
rect 42 14446 110 14514
rect 42 13240 110 13308
rect 42 11990 110 12058
rect 42 10784 110 10852
rect 42 9534 110 9602
rect 42 8328 110 8396
rect 42 7078 110 7146
rect 42 5872 110 5940
rect 42 4622 110 4690
rect 42 3416 110 3484
rect 42 2166 110 2234
rect 42 960 110 1028
rect 144 18682 212 18750
rect 1374 18725 1430 18727
rect 1454 18725 1510 18727
rect 1534 18725 1590 18727
rect 1614 18725 1670 18727
rect 1694 18725 1750 18727
rect 1774 18725 1830 18727
rect 1854 18725 1910 18727
rect 1374 18673 1412 18725
rect 1412 18673 1424 18725
rect 1424 18673 1430 18725
rect 1454 18673 1476 18725
rect 1476 18673 1488 18725
rect 1488 18673 1510 18725
rect 1534 18673 1540 18725
rect 1540 18673 1552 18725
rect 1552 18673 1590 18725
rect 1614 18673 1616 18725
rect 1616 18673 1668 18725
rect 1668 18673 1670 18725
rect 1694 18673 1732 18725
rect 1732 18673 1744 18725
rect 1744 18673 1750 18725
rect 1774 18673 1796 18725
rect 1796 18673 1808 18725
rect 1808 18673 1830 18725
rect 1854 18673 1860 18725
rect 1860 18673 1872 18725
rect 1872 18673 1910 18725
rect 1374 18671 1430 18673
rect 1454 18671 1510 18673
rect 1534 18671 1590 18673
rect 1614 18671 1670 18673
rect 1694 18671 1750 18673
rect 1774 18671 1830 18673
rect 1854 18671 1910 18673
rect 3746 18736 3802 18738
rect 3826 18736 3882 18738
rect 3906 18736 3962 18738
rect 3986 18736 4042 18738
rect 4066 18736 4122 18738
rect 4146 18736 4202 18738
rect 3746 18684 3756 18736
rect 3756 18684 3802 18736
rect 3826 18684 3872 18736
rect 3872 18684 3882 18736
rect 3906 18684 3936 18736
rect 3936 18684 3948 18736
rect 3948 18684 3962 18736
rect 3986 18684 4000 18736
rect 4000 18684 4012 18736
rect 4012 18684 4042 18736
rect 4066 18684 4076 18736
rect 4076 18684 4122 18736
rect 4146 18684 4192 18736
rect 4192 18684 4202 18736
rect 3746 18682 3802 18684
rect 3826 18682 3882 18684
rect 3906 18682 3962 18684
rect 3986 18682 4042 18684
rect 4066 18682 4122 18684
rect 4146 18682 4202 18684
rect 1388 18199 1444 18201
rect 1468 18199 1524 18201
rect 1548 18199 1604 18201
rect 1628 18199 1684 18201
rect 1708 18199 1764 18201
rect 1788 18199 1844 18201
rect 1388 18147 1398 18199
rect 1398 18147 1444 18199
rect 1468 18147 1514 18199
rect 1514 18147 1524 18199
rect 1548 18147 1578 18199
rect 1578 18147 1590 18199
rect 1590 18147 1604 18199
rect 1628 18147 1642 18199
rect 1642 18147 1654 18199
rect 1654 18147 1684 18199
rect 1708 18147 1718 18199
rect 1718 18147 1764 18199
rect 1788 18147 1834 18199
rect 1834 18147 1844 18199
rect 1388 18145 1444 18147
rect 1468 18145 1524 18147
rect 1548 18145 1604 18147
rect 1628 18145 1684 18147
rect 1708 18145 1764 18147
rect 1788 18145 1844 18147
rect 1932 17893 1988 17894
rect 1932 17841 1935 17893
rect 1935 17841 1987 17893
rect 1987 17841 1988 17893
rect 1932 17838 1988 17841
rect 3766 18198 3822 18200
rect 3846 18198 3902 18200
rect 3926 18198 3982 18200
rect 4006 18198 4062 18200
rect 4086 18198 4142 18200
rect 4166 18198 4222 18200
rect 3766 18146 3776 18198
rect 3776 18146 3822 18198
rect 3846 18146 3892 18198
rect 3892 18146 3902 18198
rect 3926 18146 3956 18198
rect 3956 18146 3968 18198
rect 3968 18146 3982 18198
rect 4006 18146 4020 18198
rect 4020 18146 4032 18198
rect 4032 18146 4062 18198
rect 4086 18146 4096 18198
rect 4096 18146 4142 18198
rect 4166 18146 4212 18198
rect 4212 18146 4222 18198
rect 3766 18144 3822 18146
rect 3846 18144 3902 18146
rect 3926 18144 3982 18146
rect 4006 18144 4062 18146
rect 4086 18144 4142 18146
rect 4166 18144 4222 18146
rect 2520 17680 2576 17682
rect 2520 17628 2522 17680
rect 2522 17628 2574 17680
rect 2574 17628 2576 17680
rect 2520 17626 2576 17628
rect 5704 18736 5760 18738
rect 5784 18736 5840 18738
rect 5864 18736 5920 18738
rect 5944 18736 6000 18738
rect 6024 18736 6080 18738
rect 6104 18736 6160 18738
rect 5704 18684 5714 18736
rect 5714 18684 5760 18736
rect 5784 18684 5830 18736
rect 5830 18684 5840 18736
rect 5864 18684 5894 18736
rect 5894 18684 5906 18736
rect 5906 18684 5920 18736
rect 5944 18684 5958 18736
rect 5958 18684 5970 18736
rect 5970 18684 6000 18736
rect 6024 18684 6034 18736
rect 6034 18684 6080 18736
rect 6104 18684 6150 18736
rect 6150 18684 6160 18736
rect 5704 18682 5760 18684
rect 5784 18682 5840 18684
rect 5864 18682 5920 18684
rect 5944 18682 6000 18684
rect 6024 18682 6080 18684
rect 6104 18682 6160 18684
rect 5724 18198 5780 18200
rect 5804 18198 5860 18200
rect 5884 18198 5940 18200
rect 5964 18198 6020 18200
rect 6044 18198 6100 18200
rect 6124 18198 6180 18200
rect 5724 18146 5734 18198
rect 5734 18146 5780 18198
rect 5804 18146 5850 18198
rect 5850 18146 5860 18198
rect 5884 18146 5914 18198
rect 5914 18146 5926 18198
rect 5926 18146 5940 18198
rect 5964 18146 5978 18198
rect 5978 18146 5990 18198
rect 5990 18146 6020 18198
rect 6044 18146 6054 18198
rect 6054 18146 6100 18198
rect 6124 18146 6170 18198
rect 6170 18146 6180 18198
rect 5724 18144 5780 18146
rect 5804 18144 5860 18146
rect 5884 18144 5940 18146
rect 5964 18144 6020 18146
rect 6044 18144 6100 18146
rect 6124 18144 6180 18146
rect 144 17446 212 17514
rect 1374 17497 1430 17499
rect 1454 17497 1510 17499
rect 1534 17497 1590 17499
rect 1614 17497 1670 17499
rect 1694 17497 1750 17499
rect 1774 17497 1830 17499
rect 1854 17497 1910 17499
rect 1374 17445 1412 17497
rect 1412 17445 1424 17497
rect 1424 17445 1430 17497
rect 1454 17445 1476 17497
rect 1476 17445 1488 17497
rect 1488 17445 1510 17497
rect 1534 17445 1540 17497
rect 1540 17445 1552 17497
rect 1552 17445 1590 17497
rect 1614 17445 1616 17497
rect 1616 17445 1668 17497
rect 1668 17445 1670 17497
rect 1694 17445 1732 17497
rect 1732 17445 1744 17497
rect 1744 17445 1750 17497
rect 1774 17445 1796 17497
rect 1796 17445 1808 17497
rect 1808 17445 1830 17497
rect 1854 17445 1860 17497
rect 1860 17445 1872 17497
rect 1872 17445 1910 17497
rect 1374 17443 1430 17445
rect 1454 17443 1510 17445
rect 1534 17443 1590 17445
rect 1614 17443 1670 17445
rect 1694 17443 1750 17445
rect 1774 17443 1830 17445
rect 1854 17443 1910 17445
rect 3746 17508 3802 17510
rect 3826 17508 3882 17510
rect 3906 17508 3962 17510
rect 3986 17508 4042 17510
rect 4066 17508 4122 17510
rect 4146 17508 4202 17510
rect 3746 17456 3756 17508
rect 3756 17456 3802 17508
rect 3826 17456 3872 17508
rect 3872 17456 3882 17508
rect 3906 17456 3936 17508
rect 3936 17456 3948 17508
rect 3948 17456 3962 17508
rect 3986 17456 4000 17508
rect 4000 17456 4012 17508
rect 4012 17456 4042 17508
rect 4066 17456 4076 17508
rect 4076 17456 4122 17508
rect 4146 17456 4192 17508
rect 4192 17456 4202 17508
rect 3746 17454 3802 17456
rect 3826 17454 3882 17456
rect 3906 17454 3962 17456
rect 3986 17454 4042 17456
rect 4066 17454 4122 17456
rect 4146 17454 4202 17456
rect 1388 16971 1444 16973
rect 1468 16971 1524 16973
rect 1548 16971 1604 16973
rect 1628 16971 1684 16973
rect 1708 16971 1764 16973
rect 1788 16971 1844 16973
rect 1388 16919 1398 16971
rect 1398 16919 1444 16971
rect 1468 16919 1514 16971
rect 1514 16919 1524 16971
rect 1548 16919 1578 16971
rect 1578 16919 1590 16971
rect 1590 16919 1604 16971
rect 1628 16919 1642 16971
rect 1642 16919 1654 16971
rect 1654 16919 1684 16971
rect 1708 16919 1718 16971
rect 1718 16919 1764 16971
rect 1788 16919 1834 16971
rect 1834 16919 1844 16971
rect 1388 16917 1444 16919
rect 1468 16917 1524 16919
rect 1548 16917 1604 16919
rect 1628 16917 1684 16919
rect 1708 16917 1764 16919
rect 1788 16917 1844 16919
rect 1932 16665 1988 16666
rect 1932 16613 1935 16665
rect 1935 16613 1987 16665
rect 1987 16613 1988 16665
rect 1932 16610 1988 16613
rect 3766 16970 3822 16972
rect 3846 16970 3902 16972
rect 3926 16970 3982 16972
rect 4006 16970 4062 16972
rect 4086 16970 4142 16972
rect 4166 16970 4222 16972
rect 3766 16918 3776 16970
rect 3776 16918 3822 16970
rect 3846 16918 3892 16970
rect 3892 16918 3902 16970
rect 3926 16918 3956 16970
rect 3956 16918 3968 16970
rect 3968 16918 3982 16970
rect 4006 16918 4020 16970
rect 4020 16918 4032 16970
rect 4032 16918 4062 16970
rect 4086 16918 4096 16970
rect 4096 16918 4142 16970
rect 4166 16918 4212 16970
rect 4212 16918 4222 16970
rect 3766 16916 3822 16918
rect 3846 16916 3902 16918
rect 3926 16916 3982 16918
rect 4006 16916 4062 16918
rect 4086 16916 4142 16918
rect 4166 16916 4222 16918
rect 2520 16452 2576 16454
rect 2520 16400 2522 16452
rect 2522 16400 2574 16452
rect 2574 16400 2576 16452
rect 2520 16398 2576 16400
rect 5704 17508 5760 17510
rect 5784 17508 5840 17510
rect 5864 17508 5920 17510
rect 5944 17508 6000 17510
rect 6024 17508 6080 17510
rect 6104 17508 6160 17510
rect 5704 17456 5714 17508
rect 5714 17456 5760 17508
rect 5784 17456 5830 17508
rect 5830 17456 5840 17508
rect 5864 17456 5894 17508
rect 5894 17456 5906 17508
rect 5906 17456 5920 17508
rect 5944 17456 5958 17508
rect 5958 17456 5970 17508
rect 5970 17456 6000 17508
rect 6024 17456 6034 17508
rect 6034 17456 6080 17508
rect 6104 17456 6150 17508
rect 6150 17456 6160 17508
rect 5704 17454 5760 17456
rect 5784 17454 5840 17456
rect 5864 17454 5920 17456
rect 5944 17454 6000 17456
rect 6024 17454 6080 17456
rect 6104 17454 6160 17456
rect 5724 16970 5780 16972
rect 5804 16970 5860 16972
rect 5884 16970 5940 16972
rect 5964 16970 6020 16972
rect 6044 16970 6100 16972
rect 6124 16970 6180 16972
rect 5724 16918 5734 16970
rect 5734 16918 5780 16970
rect 5804 16918 5850 16970
rect 5850 16918 5860 16970
rect 5884 16918 5914 16970
rect 5914 16918 5926 16970
rect 5926 16918 5940 16970
rect 5964 16918 5978 16970
rect 5978 16918 5990 16970
rect 5990 16918 6020 16970
rect 6044 16918 6054 16970
rect 6054 16918 6100 16970
rect 6124 16918 6170 16970
rect 6170 16918 6180 16970
rect 5724 16916 5780 16918
rect 5804 16916 5860 16918
rect 5884 16916 5940 16918
rect 5964 16916 6020 16918
rect 6044 16916 6100 16918
rect 6124 16916 6180 16918
rect 144 16226 212 16294
rect 1374 16269 1430 16271
rect 1454 16269 1510 16271
rect 1534 16269 1590 16271
rect 1614 16269 1670 16271
rect 1694 16269 1750 16271
rect 1774 16269 1830 16271
rect 1854 16269 1910 16271
rect 1374 16217 1412 16269
rect 1412 16217 1424 16269
rect 1424 16217 1430 16269
rect 1454 16217 1476 16269
rect 1476 16217 1488 16269
rect 1488 16217 1510 16269
rect 1534 16217 1540 16269
rect 1540 16217 1552 16269
rect 1552 16217 1590 16269
rect 1614 16217 1616 16269
rect 1616 16217 1668 16269
rect 1668 16217 1670 16269
rect 1694 16217 1732 16269
rect 1732 16217 1744 16269
rect 1744 16217 1750 16269
rect 1774 16217 1796 16269
rect 1796 16217 1808 16269
rect 1808 16217 1830 16269
rect 1854 16217 1860 16269
rect 1860 16217 1872 16269
rect 1872 16217 1910 16269
rect 1374 16215 1430 16217
rect 1454 16215 1510 16217
rect 1534 16215 1590 16217
rect 1614 16215 1670 16217
rect 1694 16215 1750 16217
rect 1774 16215 1830 16217
rect 1854 16215 1910 16217
rect 3746 16280 3802 16282
rect 3826 16280 3882 16282
rect 3906 16280 3962 16282
rect 3986 16280 4042 16282
rect 4066 16280 4122 16282
rect 4146 16280 4202 16282
rect 3746 16228 3756 16280
rect 3756 16228 3802 16280
rect 3826 16228 3872 16280
rect 3872 16228 3882 16280
rect 3906 16228 3936 16280
rect 3936 16228 3948 16280
rect 3948 16228 3962 16280
rect 3986 16228 4000 16280
rect 4000 16228 4012 16280
rect 4012 16228 4042 16280
rect 4066 16228 4076 16280
rect 4076 16228 4122 16280
rect 4146 16228 4192 16280
rect 4192 16228 4202 16280
rect 3746 16226 3802 16228
rect 3826 16226 3882 16228
rect 3906 16226 3962 16228
rect 3986 16226 4042 16228
rect 4066 16226 4122 16228
rect 4146 16226 4202 16228
rect 1388 15743 1444 15745
rect 1468 15743 1524 15745
rect 1548 15743 1604 15745
rect 1628 15743 1684 15745
rect 1708 15743 1764 15745
rect 1788 15743 1844 15745
rect 1388 15691 1398 15743
rect 1398 15691 1444 15743
rect 1468 15691 1514 15743
rect 1514 15691 1524 15743
rect 1548 15691 1578 15743
rect 1578 15691 1590 15743
rect 1590 15691 1604 15743
rect 1628 15691 1642 15743
rect 1642 15691 1654 15743
rect 1654 15691 1684 15743
rect 1708 15691 1718 15743
rect 1718 15691 1764 15743
rect 1788 15691 1834 15743
rect 1834 15691 1844 15743
rect 1388 15689 1444 15691
rect 1468 15689 1524 15691
rect 1548 15689 1604 15691
rect 1628 15689 1684 15691
rect 1708 15689 1764 15691
rect 1788 15689 1844 15691
rect 1932 15437 1988 15438
rect 1932 15385 1935 15437
rect 1935 15385 1987 15437
rect 1987 15385 1988 15437
rect 1932 15382 1988 15385
rect 3766 15742 3822 15744
rect 3846 15742 3902 15744
rect 3926 15742 3982 15744
rect 4006 15742 4062 15744
rect 4086 15742 4142 15744
rect 4166 15742 4222 15744
rect 3766 15690 3776 15742
rect 3776 15690 3822 15742
rect 3846 15690 3892 15742
rect 3892 15690 3902 15742
rect 3926 15690 3956 15742
rect 3956 15690 3968 15742
rect 3968 15690 3982 15742
rect 4006 15690 4020 15742
rect 4020 15690 4032 15742
rect 4032 15690 4062 15742
rect 4086 15690 4096 15742
rect 4096 15690 4142 15742
rect 4166 15690 4212 15742
rect 4212 15690 4222 15742
rect 3766 15688 3822 15690
rect 3846 15688 3902 15690
rect 3926 15688 3982 15690
rect 4006 15688 4062 15690
rect 4086 15688 4142 15690
rect 4166 15688 4222 15690
rect 2520 15224 2576 15226
rect 2520 15172 2522 15224
rect 2522 15172 2574 15224
rect 2574 15172 2576 15224
rect 2520 15170 2576 15172
rect 5704 16280 5760 16282
rect 5784 16280 5840 16282
rect 5864 16280 5920 16282
rect 5944 16280 6000 16282
rect 6024 16280 6080 16282
rect 6104 16280 6160 16282
rect 5704 16228 5714 16280
rect 5714 16228 5760 16280
rect 5784 16228 5830 16280
rect 5830 16228 5840 16280
rect 5864 16228 5894 16280
rect 5894 16228 5906 16280
rect 5906 16228 5920 16280
rect 5944 16228 5958 16280
rect 5958 16228 5970 16280
rect 5970 16228 6000 16280
rect 6024 16228 6034 16280
rect 6034 16228 6080 16280
rect 6104 16228 6150 16280
rect 6150 16228 6160 16280
rect 5704 16226 5760 16228
rect 5784 16226 5840 16228
rect 5864 16226 5920 16228
rect 5944 16226 6000 16228
rect 6024 16226 6080 16228
rect 6104 16226 6160 16228
rect 5724 15742 5780 15744
rect 5804 15742 5860 15744
rect 5884 15742 5940 15744
rect 5964 15742 6020 15744
rect 6044 15742 6100 15744
rect 6124 15742 6180 15744
rect 5724 15690 5734 15742
rect 5734 15690 5780 15742
rect 5804 15690 5850 15742
rect 5850 15690 5860 15742
rect 5884 15690 5914 15742
rect 5914 15690 5926 15742
rect 5926 15690 5940 15742
rect 5964 15690 5978 15742
rect 5978 15690 5990 15742
rect 5990 15690 6020 15742
rect 6044 15690 6054 15742
rect 6054 15690 6100 15742
rect 6124 15690 6170 15742
rect 6170 15690 6180 15742
rect 5724 15688 5780 15690
rect 5804 15688 5860 15690
rect 5884 15688 5940 15690
rect 5964 15688 6020 15690
rect 6044 15688 6100 15690
rect 6124 15688 6180 15690
rect 144 14990 212 15058
rect 1374 15041 1430 15043
rect 1454 15041 1510 15043
rect 1534 15041 1590 15043
rect 1614 15041 1670 15043
rect 1694 15041 1750 15043
rect 1774 15041 1830 15043
rect 1854 15041 1910 15043
rect 1374 14989 1412 15041
rect 1412 14989 1424 15041
rect 1424 14989 1430 15041
rect 1454 14989 1476 15041
rect 1476 14989 1488 15041
rect 1488 14989 1510 15041
rect 1534 14989 1540 15041
rect 1540 14989 1552 15041
rect 1552 14989 1590 15041
rect 1614 14989 1616 15041
rect 1616 14989 1668 15041
rect 1668 14989 1670 15041
rect 1694 14989 1732 15041
rect 1732 14989 1744 15041
rect 1744 14989 1750 15041
rect 1774 14989 1796 15041
rect 1796 14989 1808 15041
rect 1808 14989 1830 15041
rect 1854 14989 1860 15041
rect 1860 14989 1872 15041
rect 1872 14989 1910 15041
rect 1374 14987 1430 14989
rect 1454 14987 1510 14989
rect 1534 14987 1590 14989
rect 1614 14987 1670 14989
rect 1694 14987 1750 14989
rect 1774 14987 1830 14989
rect 1854 14987 1910 14989
rect 3746 15052 3802 15054
rect 3826 15052 3882 15054
rect 3906 15052 3962 15054
rect 3986 15052 4042 15054
rect 4066 15052 4122 15054
rect 4146 15052 4202 15054
rect 3746 15000 3756 15052
rect 3756 15000 3802 15052
rect 3826 15000 3872 15052
rect 3872 15000 3882 15052
rect 3906 15000 3936 15052
rect 3936 15000 3948 15052
rect 3948 15000 3962 15052
rect 3986 15000 4000 15052
rect 4000 15000 4012 15052
rect 4012 15000 4042 15052
rect 4066 15000 4076 15052
rect 4076 15000 4122 15052
rect 4146 15000 4192 15052
rect 4192 15000 4202 15052
rect 3746 14998 3802 15000
rect 3826 14998 3882 15000
rect 3906 14998 3962 15000
rect 3986 14998 4042 15000
rect 4066 14998 4122 15000
rect 4146 14998 4202 15000
rect 1388 14515 1444 14517
rect 1468 14515 1524 14517
rect 1548 14515 1604 14517
rect 1628 14515 1684 14517
rect 1708 14515 1764 14517
rect 1788 14515 1844 14517
rect 1388 14463 1398 14515
rect 1398 14463 1444 14515
rect 1468 14463 1514 14515
rect 1514 14463 1524 14515
rect 1548 14463 1578 14515
rect 1578 14463 1590 14515
rect 1590 14463 1604 14515
rect 1628 14463 1642 14515
rect 1642 14463 1654 14515
rect 1654 14463 1684 14515
rect 1708 14463 1718 14515
rect 1718 14463 1764 14515
rect 1788 14463 1834 14515
rect 1834 14463 1844 14515
rect 1388 14461 1444 14463
rect 1468 14461 1524 14463
rect 1548 14461 1604 14463
rect 1628 14461 1684 14463
rect 1708 14461 1764 14463
rect 1788 14461 1844 14463
rect 1932 14209 1988 14210
rect 1932 14157 1935 14209
rect 1935 14157 1987 14209
rect 1987 14157 1988 14209
rect 1932 14154 1988 14157
rect 3766 14514 3822 14516
rect 3846 14514 3902 14516
rect 3926 14514 3982 14516
rect 4006 14514 4062 14516
rect 4086 14514 4142 14516
rect 4166 14514 4222 14516
rect 3766 14462 3776 14514
rect 3776 14462 3822 14514
rect 3846 14462 3892 14514
rect 3892 14462 3902 14514
rect 3926 14462 3956 14514
rect 3956 14462 3968 14514
rect 3968 14462 3982 14514
rect 4006 14462 4020 14514
rect 4020 14462 4032 14514
rect 4032 14462 4062 14514
rect 4086 14462 4096 14514
rect 4096 14462 4142 14514
rect 4166 14462 4212 14514
rect 4212 14462 4222 14514
rect 3766 14460 3822 14462
rect 3846 14460 3902 14462
rect 3926 14460 3982 14462
rect 4006 14460 4062 14462
rect 4086 14460 4142 14462
rect 4166 14460 4222 14462
rect 2520 13996 2576 13998
rect 2520 13944 2522 13996
rect 2522 13944 2574 13996
rect 2574 13944 2576 13996
rect 2520 13942 2576 13944
rect 5704 15052 5760 15054
rect 5784 15052 5840 15054
rect 5864 15052 5920 15054
rect 5944 15052 6000 15054
rect 6024 15052 6080 15054
rect 6104 15052 6160 15054
rect 5704 15000 5714 15052
rect 5714 15000 5760 15052
rect 5784 15000 5830 15052
rect 5830 15000 5840 15052
rect 5864 15000 5894 15052
rect 5894 15000 5906 15052
rect 5906 15000 5920 15052
rect 5944 15000 5958 15052
rect 5958 15000 5970 15052
rect 5970 15000 6000 15052
rect 6024 15000 6034 15052
rect 6034 15000 6080 15052
rect 6104 15000 6150 15052
rect 6150 15000 6160 15052
rect 5704 14998 5760 15000
rect 5784 14998 5840 15000
rect 5864 14998 5920 15000
rect 5944 14998 6000 15000
rect 6024 14998 6080 15000
rect 6104 14998 6160 15000
rect 5724 14514 5780 14516
rect 5804 14514 5860 14516
rect 5884 14514 5940 14516
rect 5964 14514 6020 14516
rect 6044 14514 6100 14516
rect 6124 14514 6180 14516
rect 5724 14462 5734 14514
rect 5734 14462 5780 14514
rect 5804 14462 5850 14514
rect 5850 14462 5860 14514
rect 5884 14462 5914 14514
rect 5914 14462 5926 14514
rect 5926 14462 5940 14514
rect 5964 14462 5978 14514
rect 5978 14462 5990 14514
rect 5990 14462 6020 14514
rect 6044 14462 6054 14514
rect 6054 14462 6100 14514
rect 6124 14462 6170 14514
rect 6170 14462 6180 14514
rect 5724 14460 5780 14462
rect 5804 14460 5860 14462
rect 5884 14460 5940 14462
rect 5964 14460 6020 14462
rect 6044 14460 6100 14462
rect 6124 14460 6180 14462
rect 144 13770 212 13838
rect 1374 13813 1430 13815
rect 1454 13813 1510 13815
rect 1534 13813 1590 13815
rect 1614 13813 1670 13815
rect 1694 13813 1750 13815
rect 1774 13813 1830 13815
rect 1854 13813 1910 13815
rect 1374 13761 1412 13813
rect 1412 13761 1424 13813
rect 1424 13761 1430 13813
rect 1454 13761 1476 13813
rect 1476 13761 1488 13813
rect 1488 13761 1510 13813
rect 1534 13761 1540 13813
rect 1540 13761 1552 13813
rect 1552 13761 1590 13813
rect 1614 13761 1616 13813
rect 1616 13761 1668 13813
rect 1668 13761 1670 13813
rect 1694 13761 1732 13813
rect 1732 13761 1744 13813
rect 1744 13761 1750 13813
rect 1774 13761 1796 13813
rect 1796 13761 1808 13813
rect 1808 13761 1830 13813
rect 1854 13761 1860 13813
rect 1860 13761 1872 13813
rect 1872 13761 1910 13813
rect 1374 13759 1430 13761
rect 1454 13759 1510 13761
rect 1534 13759 1590 13761
rect 1614 13759 1670 13761
rect 1694 13759 1750 13761
rect 1774 13759 1830 13761
rect 1854 13759 1910 13761
rect 3746 13824 3802 13826
rect 3826 13824 3882 13826
rect 3906 13824 3962 13826
rect 3986 13824 4042 13826
rect 4066 13824 4122 13826
rect 4146 13824 4202 13826
rect 3746 13772 3756 13824
rect 3756 13772 3802 13824
rect 3826 13772 3872 13824
rect 3872 13772 3882 13824
rect 3906 13772 3936 13824
rect 3936 13772 3948 13824
rect 3948 13772 3962 13824
rect 3986 13772 4000 13824
rect 4000 13772 4012 13824
rect 4012 13772 4042 13824
rect 4066 13772 4076 13824
rect 4076 13772 4122 13824
rect 4146 13772 4192 13824
rect 4192 13772 4202 13824
rect 3746 13770 3802 13772
rect 3826 13770 3882 13772
rect 3906 13770 3962 13772
rect 3986 13770 4042 13772
rect 4066 13770 4122 13772
rect 4146 13770 4202 13772
rect 1388 13287 1444 13289
rect 1468 13287 1524 13289
rect 1548 13287 1604 13289
rect 1628 13287 1684 13289
rect 1708 13287 1764 13289
rect 1788 13287 1844 13289
rect 1388 13235 1398 13287
rect 1398 13235 1444 13287
rect 1468 13235 1514 13287
rect 1514 13235 1524 13287
rect 1548 13235 1578 13287
rect 1578 13235 1590 13287
rect 1590 13235 1604 13287
rect 1628 13235 1642 13287
rect 1642 13235 1654 13287
rect 1654 13235 1684 13287
rect 1708 13235 1718 13287
rect 1718 13235 1764 13287
rect 1788 13235 1834 13287
rect 1834 13235 1844 13287
rect 1388 13233 1444 13235
rect 1468 13233 1524 13235
rect 1548 13233 1604 13235
rect 1628 13233 1684 13235
rect 1708 13233 1764 13235
rect 1788 13233 1844 13235
rect 1932 12981 1988 12982
rect 1932 12929 1935 12981
rect 1935 12929 1987 12981
rect 1987 12929 1988 12981
rect 1932 12926 1988 12929
rect 3766 13286 3822 13288
rect 3846 13286 3902 13288
rect 3926 13286 3982 13288
rect 4006 13286 4062 13288
rect 4086 13286 4142 13288
rect 4166 13286 4222 13288
rect 3766 13234 3776 13286
rect 3776 13234 3822 13286
rect 3846 13234 3892 13286
rect 3892 13234 3902 13286
rect 3926 13234 3956 13286
rect 3956 13234 3968 13286
rect 3968 13234 3982 13286
rect 4006 13234 4020 13286
rect 4020 13234 4032 13286
rect 4032 13234 4062 13286
rect 4086 13234 4096 13286
rect 4096 13234 4142 13286
rect 4166 13234 4212 13286
rect 4212 13234 4222 13286
rect 3766 13232 3822 13234
rect 3846 13232 3902 13234
rect 3926 13232 3982 13234
rect 4006 13232 4062 13234
rect 4086 13232 4142 13234
rect 4166 13232 4222 13234
rect 2520 12768 2576 12770
rect 2520 12716 2522 12768
rect 2522 12716 2574 12768
rect 2574 12716 2576 12768
rect 2520 12714 2576 12716
rect 5704 13824 5760 13826
rect 5784 13824 5840 13826
rect 5864 13824 5920 13826
rect 5944 13824 6000 13826
rect 6024 13824 6080 13826
rect 6104 13824 6160 13826
rect 5704 13772 5714 13824
rect 5714 13772 5760 13824
rect 5784 13772 5830 13824
rect 5830 13772 5840 13824
rect 5864 13772 5894 13824
rect 5894 13772 5906 13824
rect 5906 13772 5920 13824
rect 5944 13772 5958 13824
rect 5958 13772 5970 13824
rect 5970 13772 6000 13824
rect 6024 13772 6034 13824
rect 6034 13772 6080 13824
rect 6104 13772 6150 13824
rect 6150 13772 6160 13824
rect 5704 13770 5760 13772
rect 5784 13770 5840 13772
rect 5864 13770 5920 13772
rect 5944 13770 6000 13772
rect 6024 13770 6080 13772
rect 6104 13770 6160 13772
rect 5724 13286 5780 13288
rect 5804 13286 5860 13288
rect 5884 13286 5940 13288
rect 5964 13286 6020 13288
rect 6044 13286 6100 13288
rect 6124 13286 6180 13288
rect 5724 13234 5734 13286
rect 5734 13234 5780 13286
rect 5804 13234 5850 13286
rect 5850 13234 5860 13286
rect 5884 13234 5914 13286
rect 5914 13234 5926 13286
rect 5926 13234 5940 13286
rect 5964 13234 5978 13286
rect 5978 13234 5990 13286
rect 5990 13234 6020 13286
rect 6044 13234 6054 13286
rect 6054 13234 6100 13286
rect 6124 13234 6170 13286
rect 6170 13234 6180 13286
rect 5724 13232 5780 13234
rect 5804 13232 5860 13234
rect 5884 13232 5940 13234
rect 5964 13232 6020 13234
rect 6044 13232 6100 13234
rect 6124 13232 6180 13234
rect 144 12534 212 12602
rect 1374 12585 1430 12587
rect 1454 12585 1510 12587
rect 1534 12585 1590 12587
rect 1614 12585 1670 12587
rect 1694 12585 1750 12587
rect 1774 12585 1830 12587
rect 1854 12585 1910 12587
rect 1374 12533 1412 12585
rect 1412 12533 1424 12585
rect 1424 12533 1430 12585
rect 1454 12533 1476 12585
rect 1476 12533 1488 12585
rect 1488 12533 1510 12585
rect 1534 12533 1540 12585
rect 1540 12533 1552 12585
rect 1552 12533 1590 12585
rect 1614 12533 1616 12585
rect 1616 12533 1668 12585
rect 1668 12533 1670 12585
rect 1694 12533 1732 12585
rect 1732 12533 1744 12585
rect 1744 12533 1750 12585
rect 1774 12533 1796 12585
rect 1796 12533 1808 12585
rect 1808 12533 1830 12585
rect 1854 12533 1860 12585
rect 1860 12533 1872 12585
rect 1872 12533 1910 12585
rect 1374 12531 1430 12533
rect 1454 12531 1510 12533
rect 1534 12531 1590 12533
rect 1614 12531 1670 12533
rect 1694 12531 1750 12533
rect 1774 12531 1830 12533
rect 1854 12531 1910 12533
rect 3746 12596 3802 12598
rect 3826 12596 3882 12598
rect 3906 12596 3962 12598
rect 3986 12596 4042 12598
rect 4066 12596 4122 12598
rect 4146 12596 4202 12598
rect 3746 12544 3756 12596
rect 3756 12544 3802 12596
rect 3826 12544 3872 12596
rect 3872 12544 3882 12596
rect 3906 12544 3936 12596
rect 3936 12544 3948 12596
rect 3948 12544 3962 12596
rect 3986 12544 4000 12596
rect 4000 12544 4012 12596
rect 4012 12544 4042 12596
rect 4066 12544 4076 12596
rect 4076 12544 4122 12596
rect 4146 12544 4192 12596
rect 4192 12544 4202 12596
rect 3746 12542 3802 12544
rect 3826 12542 3882 12544
rect 3906 12542 3962 12544
rect 3986 12542 4042 12544
rect 4066 12542 4122 12544
rect 4146 12542 4202 12544
rect 1388 12059 1444 12061
rect 1468 12059 1524 12061
rect 1548 12059 1604 12061
rect 1628 12059 1684 12061
rect 1708 12059 1764 12061
rect 1788 12059 1844 12061
rect 1388 12007 1398 12059
rect 1398 12007 1444 12059
rect 1468 12007 1514 12059
rect 1514 12007 1524 12059
rect 1548 12007 1578 12059
rect 1578 12007 1590 12059
rect 1590 12007 1604 12059
rect 1628 12007 1642 12059
rect 1642 12007 1654 12059
rect 1654 12007 1684 12059
rect 1708 12007 1718 12059
rect 1718 12007 1764 12059
rect 1788 12007 1834 12059
rect 1834 12007 1844 12059
rect 1388 12005 1444 12007
rect 1468 12005 1524 12007
rect 1548 12005 1604 12007
rect 1628 12005 1684 12007
rect 1708 12005 1764 12007
rect 1788 12005 1844 12007
rect 1932 11753 1988 11754
rect 1932 11701 1935 11753
rect 1935 11701 1987 11753
rect 1987 11701 1988 11753
rect 1932 11698 1988 11701
rect 3766 12058 3822 12060
rect 3846 12058 3902 12060
rect 3926 12058 3982 12060
rect 4006 12058 4062 12060
rect 4086 12058 4142 12060
rect 4166 12058 4222 12060
rect 3766 12006 3776 12058
rect 3776 12006 3822 12058
rect 3846 12006 3892 12058
rect 3892 12006 3902 12058
rect 3926 12006 3956 12058
rect 3956 12006 3968 12058
rect 3968 12006 3982 12058
rect 4006 12006 4020 12058
rect 4020 12006 4032 12058
rect 4032 12006 4062 12058
rect 4086 12006 4096 12058
rect 4096 12006 4142 12058
rect 4166 12006 4212 12058
rect 4212 12006 4222 12058
rect 3766 12004 3822 12006
rect 3846 12004 3902 12006
rect 3926 12004 3982 12006
rect 4006 12004 4062 12006
rect 4086 12004 4142 12006
rect 4166 12004 4222 12006
rect 2520 11540 2576 11542
rect 2520 11488 2522 11540
rect 2522 11488 2574 11540
rect 2574 11488 2576 11540
rect 2520 11486 2576 11488
rect 5704 12596 5760 12598
rect 5784 12596 5840 12598
rect 5864 12596 5920 12598
rect 5944 12596 6000 12598
rect 6024 12596 6080 12598
rect 6104 12596 6160 12598
rect 5704 12544 5714 12596
rect 5714 12544 5760 12596
rect 5784 12544 5830 12596
rect 5830 12544 5840 12596
rect 5864 12544 5894 12596
rect 5894 12544 5906 12596
rect 5906 12544 5920 12596
rect 5944 12544 5958 12596
rect 5958 12544 5970 12596
rect 5970 12544 6000 12596
rect 6024 12544 6034 12596
rect 6034 12544 6080 12596
rect 6104 12544 6150 12596
rect 6150 12544 6160 12596
rect 5704 12542 5760 12544
rect 5784 12542 5840 12544
rect 5864 12542 5920 12544
rect 5944 12542 6000 12544
rect 6024 12542 6080 12544
rect 6104 12542 6160 12544
rect 5724 12058 5780 12060
rect 5804 12058 5860 12060
rect 5884 12058 5940 12060
rect 5964 12058 6020 12060
rect 6044 12058 6100 12060
rect 6124 12058 6180 12060
rect 5724 12006 5734 12058
rect 5734 12006 5780 12058
rect 5804 12006 5850 12058
rect 5850 12006 5860 12058
rect 5884 12006 5914 12058
rect 5914 12006 5926 12058
rect 5926 12006 5940 12058
rect 5964 12006 5978 12058
rect 5978 12006 5990 12058
rect 5990 12006 6020 12058
rect 6044 12006 6054 12058
rect 6054 12006 6100 12058
rect 6124 12006 6170 12058
rect 6170 12006 6180 12058
rect 5724 12004 5780 12006
rect 5804 12004 5860 12006
rect 5884 12004 5940 12006
rect 5964 12004 6020 12006
rect 6044 12004 6100 12006
rect 6124 12004 6180 12006
rect 144 11314 212 11382
rect 1374 11357 1430 11359
rect 1454 11357 1510 11359
rect 1534 11357 1590 11359
rect 1614 11357 1670 11359
rect 1694 11357 1750 11359
rect 1774 11357 1830 11359
rect 1854 11357 1910 11359
rect 1374 11305 1412 11357
rect 1412 11305 1424 11357
rect 1424 11305 1430 11357
rect 1454 11305 1476 11357
rect 1476 11305 1488 11357
rect 1488 11305 1510 11357
rect 1534 11305 1540 11357
rect 1540 11305 1552 11357
rect 1552 11305 1590 11357
rect 1614 11305 1616 11357
rect 1616 11305 1668 11357
rect 1668 11305 1670 11357
rect 1694 11305 1732 11357
rect 1732 11305 1744 11357
rect 1744 11305 1750 11357
rect 1774 11305 1796 11357
rect 1796 11305 1808 11357
rect 1808 11305 1830 11357
rect 1854 11305 1860 11357
rect 1860 11305 1872 11357
rect 1872 11305 1910 11357
rect 1374 11303 1430 11305
rect 1454 11303 1510 11305
rect 1534 11303 1590 11305
rect 1614 11303 1670 11305
rect 1694 11303 1750 11305
rect 1774 11303 1830 11305
rect 1854 11303 1910 11305
rect 3746 11368 3802 11370
rect 3826 11368 3882 11370
rect 3906 11368 3962 11370
rect 3986 11368 4042 11370
rect 4066 11368 4122 11370
rect 4146 11368 4202 11370
rect 3746 11316 3756 11368
rect 3756 11316 3802 11368
rect 3826 11316 3872 11368
rect 3872 11316 3882 11368
rect 3906 11316 3936 11368
rect 3936 11316 3948 11368
rect 3948 11316 3962 11368
rect 3986 11316 4000 11368
rect 4000 11316 4012 11368
rect 4012 11316 4042 11368
rect 4066 11316 4076 11368
rect 4076 11316 4122 11368
rect 4146 11316 4192 11368
rect 4192 11316 4202 11368
rect 3746 11314 3802 11316
rect 3826 11314 3882 11316
rect 3906 11314 3962 11316
rect 3986 11314 4042 11316
rect 4066 11314 4122 11316
rect 4146 11314 4202 11316
rect 1388 10831 1444 10833
rect 1468 10831 1524 10833
rect 1548 10831 1604 10833
rect 1628 10831 1684 10833
rect 1708 10831 1764 10833
rect 1788 10831 1844 10833
rect 1388 10779 1398 10831
rect 1398 10779 1444 10831
rect 1468 10779 1514 10831
rect 1514 10779 1524 10831
rect 1548 10779 1578 10831
rect 1578 10779 1590 10831
rect 1590 10779 1604 10831
rect 1628 10779 1642 10831
rect 1642 10779 1654 10831
rect 1654 10779 1684 10831
rect 1708 10779 1718 10831
rect 1718 10779 1764 10831
rect 1788 10779 1834 10831
rect 1834 10779 1844 10831
rect 1388 10777 1444 10779
rect 1468 10777 1524 10779
rect 1548 10777 1604 10779
rect 1628 10777 1684 10779
rect 1708 10777 1764 10779
rect 1788 10777 1844 10779
rect 1932 10525 1988 10526
rect 1932 10473 1935 10525
rect 1935 10473 1987 10525
rect 1987 10473 1988 10525
rect 1932 10470 1988 10473
rect 3766 10830 3822 10832
rect 3846 10830 3902 10832
rect 3926 10830 3982 10832
rect 4006 10830 4062 10832
rect 4086 10830 4142 10832
rect 4166 10830 4222 10832
rect 3766 10778 3776 10830
rect 3776 10778 3822 10830
rect 3846 10778 3892 10830
rect 3892 10778 3902 10830
rect 3926 10778 3956 10830
rect 3956 10778 3968 10830
rect 3968 10778 3982 10830
rect 4006 10778 4020 10830
rect 4020 10778 4032 10830
rect 4032 10778 4062 10830
rect 4086 10778 4096 10830
rect 4096 10778 4142 10830
rect 4166 10778 4212 10830
rect 4212 10778 4222 10830
rect 3766 10776 3822 10778
rect 3846 10776 3902 10778
rect 3926 10776 3982 10778
rect 4006 10776 4062 10778
rect 4086 10776 4142 10778
rect 4166 10776 4222 10778
rect 2520 10312 2576 10314
rect 2520 10260 2522 10312
rect 2522 10260 2574 10312
rect 2574 10260 2576 10312
rect 2520 10258 2576 10260
rect 5704 11368 5760 11370
rect 5784 11368 5840 11370
rect 5864 11368 5920 11370
rect 5944 11368 6000 11370
rect 6024 11368 6080 11370
rect 6104 11368 6160 11370
rect 5704 11316 5714 11368
rect 5714 11316 5760 11368
rect 5784 11316 5830 11368
rect 5830 11316 5840 11368
rect 5864 11316 5894 11368
rect 5894 11316 5906 11368
rect 5906 11316 5920 11368
rect 5944 11316 5958 11368
rect 5958 11316 5970 11368
rect 5970 11316 6000 11368
rect 6024 11316 6034 11368
rect 6034 11316 6080 11368
rect 6104 11316 6150 11368
rect 6150 11316 6160 11368
rect 5704 11314 5760 11316
rect 5784 11314 5840 11316
rect 5864 11314 5920 11316
rect 5944 11314 6000 11316
rect 6024 11314 6080 11316
rect 6104 11314 6160 11316
rect 5724 10830 5780 10832
rect 5804 10830 5860 10832
rect 5884 10830 5940 10832
rect 5964 10830 6020 10832
rect 6044 10830 6100 10832
rect 6124 10830 6180 10832
rect 5724 10778 5734 10830
rect 5734 10778 5780 10830
rect 5804 10778 5850 10830
rect 5850 10778 5860 10830
rect 5884 10778 5914 10830
rect 5914 10778 5926 10830
rect 5926 10778 5940 10830
rect 5964 10778 5978 10830
rect 5978 10778 5990 10830
rect 5990 10778 6020 10830
rect 6044 10778 6054 10830
rect 6054 10778 6100 10830
rect 6124 10778 6170 10830
rect 6170 10778 6180 10830
rect 5724 10776 5780 10778
rect 5804 10776 5860 10778
rect 5884 10776 5940 10778
rect 5964 10776 6020 10778
rect 6044 10776 6100 10778
rect 6124 10776 6180 10778
rect 144 10078 212 10146
rect 1374 10129 1430 10131
rect 1454 10129 1510 10131
rect 1534 10129 1590 10131
rect 1614 10129 1670 10131
rect 1694 10129 1750 10131
rect 1774 10129 1830 10131
rect 1854 10129 1910 10131
rect 1374 10077 1412 10129
rect 1412 10077 1424 10129
rect 1424 10077 1430 10129
rect 1454 10077 1476 10129
rect 1476 10077 1488 10129
rect 1488 10077 1510 10129
rect 1534 10077 1540 10129
rect 1540 10077 1552 10129
rect 1552 10077 1590 10129
rect 1614 10077 1616 10129
rect 1616 10077 1668 10129
rect 1668 10077 1670 10129
rect 1694 10077 1732 10129
rect 1732 10077 1744 10129
rect 1744 10077 1750 10129
rect 1774 10077 1796 10129
rect 1796 10077 1808 10129
rect 1808 10077 1830 10129
rect 1854 10077 1860 10129
rect 1860 10077 1872 10129
rect 1872 10077 1910 10129
rect 1374 10075 1430 10077
rect 1454 10075 1510 10077
rect 1534 10075 1590 10077
rect 1614 10075 1670 10077
rect 1694 10075 1750 10077
rect 1774 10075 1830 10077
rect 1854 10075 1910 10077
rect 3746 10140 3802 10142
rect 3826 10140 3882 10142
rect 3906 10140 3962 10142
rect 3986 10140 4042 10142
rect 4066 10140 4122 10142
rect 4146 10140 4202 10142
rect 3746 10088 3756 10140
rect 3756 10088 3802 10140
rect 3826 10088 3872 10140
rect 3872 10088 3882 10140
rect 3906 10088 3936 10140
rect 3936 10088 3948 10140
rect 3948 10088 3962 10140
rect 3986 10088 4000 10140
rect 4000 10088 4012 10140
rect 4012 10088 4042 10140
rect 4066 10088 4076 10140
rect 4076 10088 4122 10140
rect 4146 10088 4192 10140
rect 4192 10088 4202 10140
rect 3746 10086 3802 10088
rect 3826 10086 3882 10088
rect 3906 10086 3962 10088
rect 3986 10086 4042 10088
rect 4066 10086 4122 10088
rect 4146 10086 4202 10088
rect 1388 9603 1444 9605
rect 1468 9603 1524 9605
rect 1548 9603 1604 9605
rect 1628 9603 1684 9605
rect 1708 9603 1764 9605
rect 1788 9603 1844 9605
rect 1388 9551 1398 9603
rect 1398 9551 1444 9603
rect 1468 9551 1514 9603
rect 1514 9551 1524 9603
rect 1548 9551 1578 9603
rect 1578 9551 1590 9603
rect 1590 9551 1604 9603
rect 1628 9551 1642 9603
rect 1642 9551 1654 9603
rect 1654 9551 1684 9603
rect 1708 9551 1718 9603
rect 1718 9551 1764 9603
rect 1788 9551 1834 9603
rect 1834 9551 1844 9603
rect 1388 9549 1444 9551
rect 1468 9549 1524 9551
rect 1548 9549 1604 9551
rect 1628 9549 1684 9551
rect 1708 9549 1764 9551
rect 1788 9549 1844 9551
rect 1932 9297 1988 9298
rect 1932 9245 1935 9297
rect 1935 9245 1987 9297
rect 1987 9245 1988 9297
rect 1932 9242 1988 9245
rect 3766 9602 3822 9604
rect 3846 9602 3902 9604
rect 3926 9602 3982 9604
rect 4006 9602 4062 9604
rect 4086 9602 4142 9604
rect 4166 9602 4222 9604
rect 3766 9550 3776 9602
rect 3776 9550 3822 9602
rect 3846 9550 3892 9602
rect 3892 9550 3902 9602
rect 3926 9550 3956 9602
rect 3956 9550 3968 9602
rect 3968 9550 3982 9602
rect 4006 9550 4020 9602
rect 4020 9550 4032 9602
rect 4032 9550 4062 9602
rect 4086 9550 4096 9602
rect 4096 9550 4142 9602
rect 4166 9550 4212 9602
rect 4212 9550 4222 9602
rect 3766 9548 3822 9550
rect 3846 9548 3902 9550
rect 3926 9548 3982 9550
rect 4006 9548 4062 9550
rect 4086 9548 4142 9550
rect 4166 9548 4222 9550
rect 2520 9084 2576 9086
rect 2520 9032 2522 9084
rect 2522 9032 2574 9084
rect 2574 9032 2576 9084
rect 2520 9030 2576 9032
rect 5704 10140 5760 10142
rect 5784 10140 5840 10142
rect 5864 10140 5920 10142
rect 5944 10140 6000 10142
rect 6024 10140 6080 10142
rect 6104 10140 6160 10142
rect 5704 10088 5714 10140
rect 5714 10088 5760 10140
rect 5784 10088 5830 10140
rect 5830 10088 5840 10140
rect 5864 10088 5894 10140
rect 5894 10088 5906 10140
rect 5906 10088 5920 10140
rect 5944 10088 5958 10140
rect 5958 10088 5970 10140
rect 5970 10088 6000 10140
rect 6024 10088 6034 10140
rect 6034 10088 6080 10140
rect 6104 10088 6150 10140
rect 6150 10088 6160 10140
rect 5704 10086 5760 10088
rect 5784 10086 5840 10088
rect 5864 10086 5920 10088
rect 5944 10086 6000 10088
rect 6024 10086 6080 10088
rect 6104 10086 6160 10088
rect 5724 9602 5780 9604
rect 5804 9602 5860 9604
rect 5884 9602 5940 9604
rect 5964 9602 6020 9604
rect 6044 9602 6100 9604
rect 6124 9602 6180 9604
rect 5724 9550 5734 9602
rect 5734 9550 5780 9602
rect 5804 9550 5850 9602
rect 5850 9550 5860 9602
rect 5884 9550 5914 9602
rect 5914 9550 5926 9602
rect 5926 9550 5940 9602
rect 5964 9550 5978 9602
rect 5978 9550 5990 9602
rect 5990 9550 6020 9602
rect 6044 9550 6054 9602
rect 6054 9550 6100 9602
rect 6124 9550 6170 9602
rect 6170 9550 6180 9602
rect 5724 9548 5780 9550
rect 5804 9548 5860 9550
rect 5884 9548 5940 9550
rect 5964 9548 6020 9550
rect 6044 9548 6100 9550
rect 6124 9548 6180 9550
rect 144 8858 212 8926
rect 1374 8901 1430 8903
rect 1454 8901 1510 8903
rect 1534 8901 1590 8903
rect 1614 8901 1670 8903
rect 1694 8901 1750 8903
rect 1774 8901 1830 8903
rect 1854 8901 1910 8903
rect 1374 8849 1412 8901
rect 1412 8849 1424 8901
rect 1424 8849 1430 8901
rect 1454 8849 1476 8901
rect 1476 8849 1488 8901
rect 1488 8849 1510 8901
rect 1534 8849 1540 8901
rect 1540 8849 1552 8901
rect 1552 8849 1590 8901
rect 1614 8849 1616 8901
rect 1616 8849 1668 8901
rect 1668 8849 1670 8901
rect 1694 8849 1732 8901
rect 1732 8849 1744 8901
rect 1744 8849 1750 8901
rect 1774 8849 1796 8901
rect 1796 8849 1808 8901
rect 1808 8849 1830 8901
rect 1854 8849 1860 8901
rect 1860 8849 1872 8901
rect 1872 8849 1910 8901
rect 1374 8847 1430 8849
rect 1454 8847 1510 8849
rect 1534 8847 1590 8849
rect 1614 8847 1670 8849
rect 1694 8847 1750 8849
rect 1774 8847 1830 8849
rect 1854 8847 1910 8849
rect 3746 8912 3802 8914
rect 3826 8912 3882 8914
rect 3906 8912 3962 8914
rect 3986 8912 4042 8914
rect 4066 8912 4122 8914
rect 4146 8912 4202 8914
rect 3746 8860 3756 8912
rect 3756 8860 3802 8912
rect 3826 8860 3872 8912
rect 3872 8860 3882 8912
rect 3906 8860 3936 8912
rect 3936 8860 3948 8912
rect 3948 8860 3962 8912
rect 3986 8860 4000 8912
rect 4000 8860 4012 8912
rect 4012 8860 4042 8912
rect 4066 8860 4076 8912
rect 4076 8860 4122 8912
rect 4146 8860 4192 8912
rect 4192 8860 4202 8912
rect 3746 8858 3802 8860
rect 3826 8858 3882 8860
rect 3906 8858 3962 8860
rect 3986 8858 4042 8860
rect 4066 8858 4122 8860
rect 4146 8858 4202 8860
rect 1388 8375 1444 8377
rect 1468 8375 1524 8377
rect 1548 8375 1604 8377
rect 1628 8375 1684 8377
rect 1708 8375 1764 8377
rect 1788 8375 1844 8377
rect 1388 8323 1398 8375
rect 1398 8323 1444 8375
rect 1468 8323 1514 8375
rect 1514 8323 1524 8375
rect 1548 8323 1578 8375
rect 1578 8323 1590 8375
rect 1590 8323 1604 8375
rect 1628 8323 1642 8375
rect 1642 8323 1654 8375
rect 1654 8323 1684 8375
rect 1708 8323 1718 8375
rect 1718 8323 1764 8375
rect 1788 8323 1834 8375
rect 1834 8323 1844 8375
rect 1388 8321 1444 8323
rect 1468 8321 1524 8323
rect 1548 8321 1604 8323
rect 1628 8321 1684 8323
rect 1708 8321 1764 8323
rect 1788 8321 1844 8323
rect 1932 8069 1988 8070
rect 1932 8017 1935 8069
rect 1935 8017 1987 8069
rect 1987 8017 1988 8069
rect 1932 8014 1988 8017
rect 3766 8374 3822 8376
rect 3846 8374 3902 8376
rect 3926 8374 3982 8376
rect 4006 8374 4062 8376
rect 4086 8374 4142 8376
rect 4166 8374 4222 8376
rect 3766 8322 3776 8374
rect 3776 8322 3822 8374
rect 3846 8322 3892 8374
rect 3892 8322 3902 8374
rect 3926 8322 3956 8374
rect 3956 8322 3968 8374
rect 3968 8322 3982 8374
rect 4006 8322 4020 8374
rect 4020 8322 4032 8374
rect 4032 8322 4062 8374
rect 4086 8322 4096 8374
rect 4096 8322 4142 8374
rect 4166 8322 4212 8374
rect 4212 8322 4222 8374
rect 3766 8320 3822 8322
rect 3846 8320 3902 8322
rect 3926 8320 3982 8322
rect 4006 8320 4062 8322
rect 4086 8320 4142 8322
rect 4166 8320 4222 8322
rect 2520 7856 2576 7858
rect 2520 7804 2522 7856
rect 2522 7804 2574 7856
rect 2574 7804 2576 7856
rect 2520 7802 2576 7804
rect 5704 8912 5760 8914
rect 5784 8912 5840 8914
rect 5864 8912 5920 8914
rect 5944 8912 6000 8914
rect 6024 8912 6080 8914
rect 6104 8912 6160 8914
rect 5704 8860 5714 8912
rect 5714 8860 5760 8912
rect 5784 8860 5830 8912
rect 5830 8860 5840 8912
rect 5864 8860 5894 8912
rect 5894 8860 5906 8912
rect 5906 8860 5920 8912
rect 5944 8860 5958 8912
rect 5958 8860 5970 8912
rect 5970 8860 6000 8912
rect 6024 8860 6034 8912
rect 6034 8860 6080 8912
rect 6104 8860 6150 8912
rect 6150 8860 6160 8912
rect 5704 8858 5760 8860
rect 5784 8858 5840 8860
rect 5864 8858 5920 8860
rect 5944 8858 6000 8860
rect 6024 8858 6080 8860
rect 6104 8858 6160 8860
rect 5724 8374 5780 8376
rect 5804 8374 5860 8376
rect 5884 8374 5940 8376
rect 5964 8374 6020 8376
rect 6044 8374 6100 8376
rect 6124 8374 6180 8376
rect 5724 8322 5734 8374
rect 5734 8322 5780 8374
rect 5804 8322 5850 8374
rect 5850 8322 5860 8374
rect 5884 8322 5914 8374
rect 5914 8322 5926 8374
rect 5926 8322 5940 8374
rect 5964 8322 5978 8374
rect 5978 8322 5990 8374
rect 5990 8322 6020 8374
rect 6044 8322 6054 8374
rect 6054 8322 6100 8374
rect 6124 8322 6170 8374
rect 6170 8322 6180 8374
rect 5724 8320 5780 8322
rect 5804 8320 5860 8322
rect 5884 8320 5940 8322
rect 5964 8320 6020 8322
rect 6044 8320 6100 8322
rect 6124 8320 6180 8322
rect 144 7622 212 7690
rect 1374 7673 1430 7675
rect 1454 7673 1510 7675
rect 1534 7673 1590 7675
rect 1614 7673 1670 7675
rect 1694 7673 1750 7675
rect 1774 7673 1830 7675
rect 1854 7673 1910 7675
rect 1374 7621 1412 7673
rect 1412 7621 1424 7673
rect 1424 7621 1430 7673
rect 1454 7621 1476 7673
rect 1476 7621 1488 7673
rect 1488 7621 1510 7673
rect 1534 7621 1540 7673
rect 1540 7621 1552 7673
rect 1552 7621 1590 7673
rect 1614 7621 1616 7673
rect 1616 7621 1668 7673
rect 1668 7621 1670 7673
rect 1694 7621 1732 7673
rect 1732 7621 1744 7673
rect 1744 7621 1750 7673
rect 1774 7621 1796 7673
rect 1796 7621 1808 7673
rect 1808 7621 1830 7673
rect 1854 7621 1860 7673
rect 1860 7621 1872 7673
rect 1872 7621 1910 7673
rect 1374 7619 1430 7621
rect 1454 7619 1510 7621
rect 1534 7619 1590 7621
rect 1614 7619 1670 7621
rect 1694 7619 1750 7621
rect 1774 7619 1830 7621
rect 1854 7619 1910 7621
rect 3746 7684 3802 7686
rect 3826 7684 3882 7686
rect 3906 7684 3962 7686
rect 3986 7684 4042 7686
rect 4066 7684 4122 7686
rect 4146 7684 4202 7686
rect 3746 7632 3756 7684
rect 3756 7632 3802 7684
rect 3826 7632 3872 7684
rect 3872 7632 3882 7684
rect 3906 7632 3936 7684
rect 3936 7632 3948 7684
rect 3948 7632 3962 7684
rect 3986 7632 4000 7684
rect 4000 7632 4012 7684
rect 4012 7632 4042 7684
rect 4066 7632 4076 7684
rect 4076 7632 4122 7684
rect 4146 7632 4192 7684
rect 4192 7632 4202 7684
rect 3746 7630 3802 7632
rect 3826 7630 3882 7632
rect 3906 7630 3962 7632
rect 3986 7630 4042 7632
rect 4066 7630 4122 7632
rect 4146 7630 4202 7632
rect 1388 7147 1444 7149
rect 1468 7147 1524 7149
rect 1548 7147 1604 7149
rect 1628 7147 1684 7149
rect 1708 7147 1764 7149
rect 1788 7147 1844 7149
rect 1388 7095 1398 7147
rect 1398 7095 1444 7147
rect 1468 7095 1514 7147
rect 1514 7095 1524 7147
rect 1548 7095 1578 7147
rect 1578 7095 1590 7147
rect 1590 7095 1604 7147
rect 1628 7095 1642 7147
rect 1642 7095 1654 7147
rect 1654 7095 1684 7147
rect 1708 7095 1718 7147
rect 1718 7095 1764 7147
rect 1788 7095 1834 7147
rect 1834 7095 1844 7147
rect 1388 7093 1444 7095
rect 1468 7093 1524 7095
rect 1548 7093 1604 7095
rect 1628 7093 1684 7095
rect 1708 7093 1764 7095
rect 1788 7093 1844 7095
rect 1932 6841 1988 6842
rect 1932 6789 1935 6841
rect 1935 6789 1987 6841
rect 1987 6789 1988 6841
rect 1932 6786 1988 6789
rect 3766 7146 3822 7148
rect 3846 7146 3902 7148
rect 3926 7146 3982 7148
rect 4006 7146 4062 7148
rect 4086 7146 4142 7148
rect 4166 7146 4222 7148
rect 3766 7094 3776 7146
rect 3776 7094 3822 7146
rect 3846 7094 3892 7146
rect 3892 7094 3902 7146
rect 3926 7094 3956 7146
rect 3956 7094 3968 7146
rect 3968 7094 3982 7146
rect 4006 7094 4020 7146
rect 4020 7094 4032 7146
rect 4032 7094 4062 7146
rect 4086 7094 4096 7146
rect 4096 7094 4142 7146
rect 4166 7094 4212 7146
rect 4212 7094 4222 7146
rect 3766 7092 3822 7094
rect 3846 7092 3902 7094
rect 3926 7092 3982 7094
rect 4006 7092 4062 7094
rect 4086 7092 4142 7094
rect 4166 7092 4222 7094
rect 2520 6628 2576 6630
rect 2520 6576 2522 6628
rect 2522 6576 2574 6628
rect 2574 6576 2576 6628
rect 2520 6574 2576 6576
rect 5704 7684 5760 7686
rect 5784 7684 5840 7686
rect 5864 7684 5920 7686
rect 5944 7684 6000 7686
rect 6024 7684 6080 7686
rect 6104 7684 6160 7686
rect 5704 7632 5714 7684
rect 5714 7632 5760 7684
rect 5784 7632 5830 7684
rect 5830 7632 5840 7684
rect 5864 7632 5894 7684
rect 5894 7632 5906 7684
rect 5906 7632 5920 7684
rect 5944 7632 5958 7684
rect 5958 7632 5970 7684
rect 5970 7632 6000 7684
rect 6024 7632 6034 7684
rect 6034 7632 6080 7684
rect 6104 7632 6150 7684
rect 6150 7632 6160 7684
rect 5704 7630 5760 7632
rect 5784 7630 5840 7632
rect 5864 7630 5920 7632
rect 5944 7630 6000 7632
rect 6024 7630 6080 7632
rect 6104 7630 6160 7632
rect 5724 7146 5780 7148
rect 5804 7146 5860 7148
rect 5884 7146 5940 7148
rect 5964 7146 6020 7148
rect 6044 7146 6100 7148
rect 6124 7146 6180 7148
rect 5724 7094 5734 7146
rect 5734 7094 5780 7146
rect 5804 7094 5850 7146
rect 5850 7094 5860 7146
rect 5884 7094 5914 7146
rect 5914 7094 5926 7146
rect 5926 7094 5940 7146
rect 5964 7094 5978 7146
rect 5978 7094 5990 7146
rect 5990 7094 6020 7146
rect 6044 7094 6054 7146
rect 6054 7094 6100 7146
rect 6124 7094 6170 7146
rect 6170 7094 6180 7146
rect 5724 7092 5780 7094
rect 5804 7092 5860 7094
rect 5884 7092 5940 7094
rect 5964 7092 6020 7094
rect 6044 7092 6100 7094
rect 6124 7092 6180 7094
rect 144 6402 212 6470
rect 1374 6445 1430 6447
rect 1454 6445 1510 6447
rect 1534 6445 1590 6447
rect 1614 6445 1670 6447
rect 1694 6445 1750 6447
rect 1774 6445 1830 6447
rect 1854 6445 1910 6447
rect 1374 6393 1412 6445
rect 1412 6393 1424 6445
rect 1424 6393 1430 6445
rect 1454 6393 1476 6445
rect 1476 6393 1488 6445
rect 1488 6393 1510 6445
rect 1534 6393 1540 6445
rect 1540 6393 1552 6445
rect 1552 6393 1590 6445
rect 1614 6393 1616 6445
rect 1616 6393 1668 6445
rect 1668 6393 1670 6445
rect 1694 6393 1732 6445
rect 1732 6393 1744 6445
rect 1744 6393 1750 6445
rect 1774 6393 1796 6445
rect 1796 6393 1808 6445
rect 1808 6393 1830 6445
rect 1854 6393 1860 6445
rect 1860 6393 1872 6445
rect 1872 6393 1910 6445
rect 1374 6391 1430 6393
rect 1454 6391 1510 6393
rect 1534 6391 1590 6393
rect 1614 6391 1670 6393
rect 1694 6391 1750 6393
rect 1774 6391 1830 6393
rect 1854 6391 1910 6393
rect 3746 6456 3802 6458
rect 3826 6456 3882 6458
rect 3906 6456 3962 6458
rect 3986 6456 4042 6458
rect 4066 6456 4122 6458
rect 4146 6456 4202 6458
rect 3746 6404 3756 6456
rect 3756 6404 3802 6456
rect 3826 6404 3872 6456
rect 3872 6404 3882 6456
rect 3906 6404 3936 6456
rect 3936 6404 3948 6456
rect 3948 6404 3962 6456
rect 3986 6404 4000 6456
rect 4000 6404 4012 6456
rect 4012 6404 4042 6456
rect 4066 6404 4076 6456
rect 4076 6404 4122 6456
rect 4146 6404 4192 6456
rect 4192 6404 4202 6456
rect 3746 6402 3802 6404
rect 3826 6402 3882 6404
rect 3906 6402 3962 6404
rect 3986 6402 4042 6404
rect 4066 6402 4122 6404
rect 4146 6402 4202 6404
rect 1388 5919 1444 5921
rect 1468 5919 1524 5921
rect 1548 5919 1604 5921
rect 1628 5919 1684 5921
rect 1708 5919 1764 5921
rect 1788 5919 1844 5921
rect 1388 5867 1398 5919
rect 1398 5867 1444 5919
rect 1468 5867 1514 5919
rect 1514 5867 1524 5919
rect 1548 5867 1578 5919
rect 1578 5867 1590 5919
rect 1590 5867 1604 5919
rect 1628 5867 1642 5919
rect 1642 5867 1654 5919
rect 1654 5867 1684 5919
rect 1708 5867 1718 5919
rect 1718 5867 1764 5919
rect 1788 5867 1834 5919
rect 1834 5867 1844 5919
rect 1388 5865 1444 5867
rect 1468 5865 1524 5867
rect 1548 5865 1604 5867
rect 1628 5865 1684 5867
rect 1708 5865 1764 5867
rect 1788 5865 1844 5867
rect 1932 5613 1988 5614
rect 1932 5561 1935 5613
rect 1935 5561 1987 5613
rect 1987 5561 1988 5613
rect 1932 5558 1988 5561
rect 3766 5918 3822 5920
rect 3846 5918 3902 5920
rect 3926 5918 3982 5920
rect 4006 5918 4062 5920
rect 4086 5918 4142 5920
rect 4166 5918 4222 5920
rect 3766 5866 3776 5918
rect 3776 5866 3822 5918
rect 3846 5866 3892 5918
rect 3892 5866 3902 5918
rect 3926 5866 3956 5918
rect 3956 5866 3968 5918
rect 3968 5866 3982 5918
rect 4006 5866 4020 5918
rect 4020 5866 4032 5918
rect 4032 5866 4062 5918
rect 4086 5866 4096 5918
rect 4096 5866 4142 5918
rect 4166 5866 4212 5918
rect 4212 5866 4222 5918
rect 3766 5864 3822 5866
rect 3846 5864 3902 5866
rect 3926 5864 3982 5866
rect 4006 5864 4062 5866
rect 4086 5864 4142 5866
rect 4166 5864 4222 5866
rect 2520 5400 2576 5402
rect 2520 5348 2522 5400
rect 2522 5348 2574 5400
rect 2574 5348 2576 5400
rect 2520 5346 2576 5348
rect 5704 6456 5760 6458
rect 5784 6456 5840 6458
rect 5864 6456 5920 6458
rect 5944 6456 6000 6458
rect 6024 6456 6080 6458
rect 6104 6456 6160 6458
rect 5704 6404 5714 6456
rect 5714 6404 5760 6456
rect 5784 6404 5830 6456
rect 5830 6404 5840 6456
rect 5864 6404 5894 6456
rect 5894 6404 5906 6456
rect 5906 6404 5920 6456
rect 5944 6404 5958 6456
rect 5958 6404 5970 6456
rect 5970 6404 6000 6456
rect 6024 6404 6034 6456
rect 6034 6404 6080 6456
rect 6104 6404 6150 6456
rect 6150 6404 6160 6456
rect 5704 6402 5760 6404
rect 5784 6402 5840 6404
rect 5864 6402 5920 6404
rect 5944 6402 6000 6404
rect 6024 6402 6080 6404
rect 6104 6402 6160 6404
rect 5724 5918 5780 5920
rect 5804 5918 5860 5920
rect 5884 5918 5940 5920
rect 5964 5918 6020 5920
rect 6044 5918 6100 5920
rect 6124 5918 6180 5920
rect 5724 5866 5734 5918
rect 5734 5866 5780 5918
rect 5804 5866 5850 5918
rect 5850 5866 5860 5918
rect 5884 5866 5914 5918
rect 5914 5866 5926 5918
rect 5926 5866 5940 5918
rect 5964 5866 5978 5918
rect 5978 5866 5990 5918
rect 5990 5866 6020 5918
rect 6044 5866 6054 5918
rect 6054 5866 6100 5918
rect 6124 5866 6170 5918
rect 6170 5866 6180 5918
rect 5724 5864 5780 5866
rect 5804 5864 5860 5866
rect 5884 5864 5940 5866
rect 5964 5864 6020 5866
rect 6044 5864 6100 5866
rect 6124 5864 6180 5866
rect 144 5166 212 5234
rect 1374 5217 1430 5219
rect 1454 5217 1510 5219
rect 1534 5217 1590 5219
rect 1614 5217 1670 5219
rect 1694 5217 1750 5219
rect 1774 5217 1830 5219
rect 1854 5217 1910 5219
rect 1374 5165 1412 5217
rect 1412 5165 1424 5217
rect 1424 5165 1430 5217
rect 1454 5165 1476 5217
rect 1476 5165 1488 5217
rect 1488 5165 1510 5217
rect 1534 5165 1540 5217
rect 1540 5165 1552 5217
rect 1552 5165 1590 5217
rect 1614 5165 1616 5217
rect 1616 5165 1668 5217
rect 1668 5165 1670 5217
rect 1694 5165 1732 5217
rect 1732 5165 1744 5217
rect 1744 5165 1750 5217
rect 1774 5165 1796 5217
rect 1796 5165 1808 5217
rect 1808 5165 1830 5217
rect 1854 5165 1860 5217
rect 1860 5165 1872 5217
rect 1872 5165 1910 5217
rect 1374 5163 1430 5165
rect 1454 5163 1510 5165
rect 1534 5163 1590 5165
rect 1614 5163 1670 5165
rect 1694 5163 1750 5165
rect 1774 5163 1830 5165
rect 1854 5163 1910 5165
rect 3746 5228 3802 5230
rect 3826 5228 3882 5230
rect 3906 5228 3962 5230
rect 3986 5228 4042 5230
rect 4066 5228 4122 5230
rect 4146 5228 4202 5230
rect 3746 5176 3756 5228
rect 3756 5176 3802 5228
rect 3826 5176 3872 5228
rect 3872 5176 3882 5228
rect 3906 5176 3936 5228
rect 3936 5176 3948 5228
rect 3948 5176 3962 5228
rect 3986 5176 4000 5228
rect 4000 5176 4012 5228
rect 4012 5176 4042 5228
rect 4066 5176 4076 5228
rect 4076 5176 4122 5228
rect 4146 5176 4192 5228
rect 4192 5176 4202 5228
rect 3746 5174 3802 5176
rect 3826 5174 3882 5176
rect 3906 5174 3962 5176
rect 3986 5174 4042 5176
rect 4066 5174 4122 5176
rect 4146 5174 4202 5176
rect 1388 4691 1444 4693
rect 1468 4691 1524 4693
rect 1548 4691 1604 4693
rect 1628 4691 1684 4693
rect 1708 4691 1764 4693
rect 1788 4691 1844 4693
rect 1388 4639 1398 4691
rect 1398 4639 1444 4691
rect 1468 4639 1514 4691
rect 1514 4639 1524 4691
rect 1548 4639 1578 4691
rect 1578 4639 1590 4691
rect 1590 4639 1604 4691
rect 1628 4639 1642 4691
rect 1642 4639 1654 4691
rect 1654 4639 1684 4691
rect 1708 4639 1718 4691
rect 1718 4639 1764 4691
rect 1788 4639 1834 4691
rect 1834 4639 1844 4691
rect 1388 4637 1444 4639
rect 1468 4637 1524 4639
rect 1548 4637 1604 4639
rect 1628 4637 1684 4639
rect 1708 4637 1764 4639
rect 1788 4637 1844 4639
rect 1932 4385 1988 4386
rect 1932 4333 1935 4385
rect 1935 4333 1987 4385
rect 1987 4333 1988 4385
rect 1932 4330 1988 4333
rect 3766 4690 3822 4692
rect 3846 4690 3902 4692
rect 3926 4690 3982 4692
rect 4006 4690 4062 4692
rect 4086 4690 4142 4692
rect 4166 4690 4222 4692
rect 3766 4638 3776 4690
rect 3776 4638 3822 4690
rect 3846 4638 3892 4690
rect 3892 4638 3902 4690
rect 3926 4638 3956 4690
rect 3956 4638 3968 4690
rect 3968 4638 3982 4690
rect 4006 4638 4020 4690
rect 4020 4638 4032 4690
rect 4032 4638 4062 4690
rect 4086 4638 4096 4690
rect 4096 4638 4142 4690
rect 4166 4638 4212 4690
rect 4212 4638 4222 4690
rect 3766 4636 3822 4638
rect 3846 4636 3902 4638
rect 3926 4636 3982 4638
rect 4006 4636 4062 4638
rect 4086 4636 4142 4638
rect 4166 4636 4222 4638
rect 2520 4172 2576 4174
rect 2520 4120 2522 4172
rect 2522 4120 2574 4172
rect 2574 4120 2576 4172
rect 2520 4118 2576 4120
rect 5704 5228 5760 5230
rect 5784 5228 5840 5230
rect 5864 5228 5920 5230
rect 5944 5228 6000 5230
rect 6024 5228 6080 5230
rect 6104 5228 6160 5230
rect 5704 5176 5714 5228
rect 5714 5176 5760 5228
rect 5784 5176 5830 5228
rect 5830 5176 5840 5228
rect 5864 5176 5894 5228
rect 5894 5176 5906 5228
rect 5906 5176 5920 5228
rect 5944 5176 5958 5228
rect 5958 5176 5970 5228
rect 5970 5176 6000 5228
rect 6024 5176 6034 5228
rect 6034 5176 6080 5228
rect 6104 5176 6150 5228
rect 6150 5176 6160 5228
rect 5704 5174 5760 5176
rect 5784 5174 5840 5176
rect 5864 5174 5920 5176
rect 5944 5174 6000 5176
rect 6024 5174 6080 5176
rect 6104 5174 6160 5176
rect 5724 4690 5780 4692
rect 5804 4690 5860 4692
rect 5884 4690 5940 4692
rect 5964 4690 6020 4692
rect 6044 4690 6100 4692
rect 6124 4690 6180 4692
rect 5724 4638 5734 4690
rect 5734 4638 5780 4690
rect 5804 4638 5850 4690
rect 5850 4638 5860 4690
rect 5884 4638 5914 4690
rect 5914 4638 5926 4690
rect 5926 4638 5940 4690
rect 5964 4638 5978 4690
rect 5978 4638 5990 4690
rect 5990 4638 6020 4690
rect 6044 4638 6054 4690
rect 6054 4638 6100 4690
rect 6124 4638 6170 4690
rect 6170 4638 6180 4690
rect 5724 4636 5780 4638
rect 5804 4636 5860 4638
rect 5884 4636 5940 4638
rect 5964 4636 6020 4638
rect 6044 4636 6100 4638
rect 6124 4636 6180 4638
rect 144 3946 212 4014
rect 1374 3989 1430 3991
rect 1454 3989 1510 3991
rect 1534 3989 1590 3991
rect 1614 3989 1670 3991
rect 1694 3989 1750 3991
rect 1774 3989 1830 3991
rect 1854 3989 1910 3991
rect 1374 3937 1412 3989
rect 1412 3937 1424 3989
rect 1424 3937 1430 3989
rect 1454 3937 1476 3989
rect 1476 3937 1488 3989
rect 1488 3937 1510 3989
rect 1534 3937 1540 3989
rect 1540 3937 1552 3989
rect 1552 3937 1590 3989
rect 1614 3937 1616 3989
rect 1616 3937 1668 3989
rect 1668 3937 1670 3989
rect 1694 3937 1732 3989
rect 1732 3937 1744 3989
rect 1744 3937 1750 3989
rect 1774 3937 1796 3989
rect 1796 3937 1808 3989
rect 1808 3937 1830 3989
rect 1854 3937 1860 3989
rect 1860 3937 1872 3989
rect 1872 3937 1910 3989
rect 1374 3935 1430 3937
rect 1454 3935 1510 3937
rect 1534 3935 1590 3937
rect 1614 3935 1670 3937
rect 1694 3935 1750 3937
rect 1774 3935 1830 3937
rect 1854 3935 1910 3937
rect 3746 4000 3802 4002
rect 3826 4000 3882 4002
rect 3906 4000 3962 4002
rect 3986 4000 4042 4002
rect 4066 4000 4122 4002
rect 4146 4000 4202 4002
rect 3746 3948 3756 4000
rect 3756 3948 3802 4000
rect 3826 3948 3872 4000
rect 3872 3948 3882 4000
rect 3906 3948 3936 4000
rect 3936 3948 3948 4000
rect 3948 3948 3962 4000
rect 3986 3948 4000 4000
rect 4000 3948 4012 4000
rect 4012 3948 4042 4000
rect 4066 3948 4076 4000
rect 4076 3948 4122 4000
rect 4146 3948 4192 4000
rect 4192 3948 4202 4000
rect 3746 3946 3802 3948
rect 3826 3946 3882 3948
rect 3906 3946 3962 3948
rect 3986 3946 4042 3948
rect 4066 3946 4122 3948
rect 4146 3946 4202 3948
rect 1388 3463 1444 3465
rect 1468 3463 1524 3465
rect 1548 3463 1604 3465
rect 1628 3463 1684 3465
rect 1708 3463 1764 3465
rect 1788 3463 1844 3465
rect 1388 3411 1398 3463
rect 1398 3411 1444 3463
rect 1468 3411 1514 3463
rect 1514 3411 1524 3463
rect 1548 3411 1578 3463
rect 1578 3411 1590 3463
rect 1590 3411 1604 3463
rect 1628 3411 1642 3463
rect 1642 3411 1654 3463
rect 1654 3411 1684 3463
rect 1708 3411 1718 3463
rect 1718 3411 1764 3463
rect 1788 3411 1834 3463
rect 1834 3411 1844 3463
rect 1388 3409 1444 3411
rect 1468 3409 1524 3411
rect 1548 3409 1604 3411
rect 1628 3409 1684 3411
rect 1708 3409 1764 3411
rect 1788 3409 1844 3411
rect 1932 3157 1988 3158
rect 1932 3105 1935 3157
rect 1935 3105 1987 3157
rect 1987 3105 1988 3157
rect 1932 3102 1988 3105
rect 3766 3462 3822 3464
rect 3846 3462 3902 3464
rect 3926 3462 3982 3464
rect 4006 3462 4062 3464
rect 4086 3462 4142 3464
rect 4166 3462 4222 3464
rect 3766 3410 3776 3462
rect 3776 3410 3822 3462
rect 3846 3410 3892 3462
rect 3892 3410 3902 3462
rect 3926 3410 3956 3462
rect 3956 3410 3968 3462
rect 3968 3410 3982 3462
rect 4006 3410 4020 3462
rect 4020 3410 4032 3462
rect 4032 3410 4062 3462
rect 4086 3410 4096 3462
rect 4096 3410 4142 3462
rect 4166 3410 4212 3462
rect 4212 3410 4222 3462
rect 3766 3408 3822 3410
rect 3846 3408 3902 3410
rect 3926 3408 3982 3410
rect 4006 3408 4062 3410
rect 4086 3408 4142 3410
rect 4166 3408 4222 3410
rect 2520 2944 2576 2946
rect 2520 2892 2522 2944
rect 2522 2892 2574 2944
rect 2574 2892 2576 2944
rect 2520 2890 2576 2892
rect 5704 4000 5760 4002
rect 5784 4000 5840 4002
rect 5864 4000 5920 4002
rect 5944 4000 6000 4002
rect 6024 4000 6080 4002
rect 6104 4000 6160 4002
rect 5704 3948 5714 4000
rect 5714 3948 5760 4000
rect 5784 3948 5830 4000
rect 5830 3948 5840 4000
rect 5864 3948 5894 4000
rect 5894 3948 5906 4000
rect 5906 3948 5920 4000
rect 5944 3948 5958 4000
rect 5958 3948 5970 4000
rect 5970 3948 6000 4000
rect 6024 3948 6034 4000
rect 6034 3948 6080 4000
rect 6104 3948 6150 4000
rect 6150 3948 6160 4000
rect 5704 3946 5760 3948
rect 5784 3946 5840 3948
rect 5864 3946 5920 3948
rect 5944 3946 6000 3948
rect 6024 3946 6080 3948
rect 6104 3946 6160 3948
rect 5724 3462 5780 3464
rect 5804 3462 5860 3464
rect 5884 3462 5940 3464
rect 5964 3462 6020 3464
rect 6044 3462 6100 3464
rect 6124 3462 6180 3464
rect 5724 3410 5734 3462
rect 5734 3410 5780 3462
rect 5804 3410 5850 3462
rect 5850 3410 5860 3462
rect 5884 3410 5914 3462
rect 5914 3410 5926 3462
rect 5926 3410 5940 3462
rect 5964 3410 5978 3462
rect 5978 3410 5990 3462
rect 5990 3410 6020 3462
rect 6044 3410 6054 3462
rect 6054 3410 6100 3462
rect 6124 3410 6170 3462
rect 6170 3410 6180 3462
rect 5724 3408 5780 3410
rect 5804 3408 5860 3410
rect 5884 3408 5940 3410
rect 5964 3408 6020 3410
rect 6044 3408 6100 3410
rect 6124 3408 6180 3410
rect 144 2710 212 2778
rect 1374 2761 1430 2763
rect 1454 2761 1510 2763
rect 1534 2761 1590 2763
rect 1614 2761 1670 2763
rect 1694 2761 1750 2763
rect 1774 2761 1830 2763
rect 1854 2761 1910 2763
rect 1374 2709 1412 2761
rect 1412 2709 1424 2761
rect 1424 2709 1430 2761
rect 1454 2709 1476 2761
rect 1476 2709 1488 2761
rect 1488 2709 1510 2761
rect 1534 2709 1540 2761
rect 1540 2709 1552 2761
rect 1552 2709 1590 2761
rect 1614 2709 1616 2761
rect 1616 2709 1668 2761
rect 1668 2709 1670 2761
rect 1694 2709 1732 2761
rect 1732 2709 1744 2761
rect 1744 2709 1750 2761
rect 1774 2709 1796 2761
rect 1796 2709 1808 2761
rect 1808 2709 1830 2761
rect 1854 2709 1860 2761
rect 1860 2709 1872 2761
rect 1872 2709 1910 2761
rect 1374 2707 1430 2709
rect 1454 2707 1510 2709
rect 1534 2707 1590 2709
rect 1614 2707 1670 2709
rect 1694 2707 1750 2709
rect 1774 2707 1830 2709
rect 1854 2707 1910 2709
rect 3746 2772 3802 2774
rect 3826 2772 3882 2774
rect 3906 2772 3962 2774
rect 3986 2772 4042 2774
rect 4066 2772 4122 2774
rect 4146 2772 4202 2774
rect 3746 2720 3756 2772
rect 3756 2720 3802 2772
rect 3826 2720 3872 2772
rect 3872 2720 3882 2772
rect 3906 2720 3936 2772
rect 3936 2720 3948 2772
rect 3948 2720 3962 2772
rect 3986 2720 4000 2772
rect 4000 2720 4012 2772
rect 4012 2720 4042 2772
rect 4066 2720 4076 2772
rect 4076 2720 4122 2772
rect 4146 2720 4192 2772
rect 4192 2720 4202 2772
rect 3746 2718 3802 2720
rect 3826 2718 3882 2720
rect 3906 2718 3962 2720
rect 3986 2718 4042 2720
rect 4066 2718 4122 2720
rect 4146 2718 4202 2720
rect 1388 2235 1444 2237
rect 1468 2235 1524 2237
rect 1548 2235 1604 2237
rect 1628 2235 1684 2237
rect 1708 2235 1764 2237
rect 1788 2235 1844 2237
rect 1388 2183 1398 2235
rect 1398 2183 1444 2235
rect 1468 2183 1514 2235
rect 1514 2183 1524 2235
rect 1548 2183 1578 2235
rect 1578 2183 1590 2235
rect 1590 2183 1604 2235
rect 1628 2183 1642 2235
rect 1642 2183 1654 2235
rect 1654 2183 1684 2235
rect 1708 2183 1718 2235
rect 1718 2183 1764 2235
rect 1788 2183 1834 2235
rect 1834 2183 1844 2235
rect 1388 2181 1444 2183
rect 1468 2181 1524 2183
rect 1548 2181 1604 2183
rect 1628 2181 1684 2183
rect 1708 2181 1764 2183
rect 1788 2181 1844 2183
rect 1932 1929 1988 1930
rect 1932 1877 1935 1929
rect 1935 1877 1987 1929
rect 1987 1877 1988 1929
rect 1932 1874 1988 1877
rect 3766 2234 3822 2236
rect 3846 2234 3902 2236
rect 3926 2234 3982 2236
rect 4006 2234 4062 2236
rect 4086 2234 4142 2236
rect 4166 2234 4222 2236
rect 3766 2182 3776 2234
rect 3776 2182 3822 2234
rect 3846 2182 3892 2234
rect 3892 2182 3902 2234
rect 3926 2182 3956 2234
rect 3956 2182 3968 2234
rect 3968 2182 3982 2234
rect 4006 2182 4020 2234
rect 4020 2182 4032 2234
rect 4032 2182 4062 2234
rect 4086 2182 4096 2234
rect 4096 2182 4142 2234
rect 4166 2182 4212 2234
rect 4212 2182 4222 2234
rect 3766 2180 3822 2182
rect 3846 2180 3902 2182
rect 3926 2180 3982 2182
rect 4006 2180 4062 2182
rect 4086 2180 4142 2182
rect 4166 2180 4222 2182
rect 2520 1716 2576 1718
rect 2520 1664 2522 1716
rect 2522 1664 2574 1716
rect 2574 1664 2576 1716
rect 2520 1662 2576 1664
rect 5704 2772 5760 2774
rect 5784 2772 5840 2774
rect 5864 2772 5920 2774
rect 5944 2772 6000 2774
rect 6024 2772 6080 2774
rect 6104 2772 6160 2774
rect 5704 2720 5714 2772
rect 5714 2720 5760 2772
rect 5784 2720 5830 2772
rect 5830 2720 5840 2772
rect 5864 2720 5894 2772
rect 5894 2720 5906 2772
rect 5906 2720 5920 2772
rect 5944 2720 5958 2772
rect 5958 2720 5970 2772
rect 5970 2720 6000 2772
rect 6024 2720 6034 2772
rect 6034 2720 6080 2772
rect 6104 2720 6150 2772
rect 6150 2720 6160 2772
rect 5704 2718 5760 2720
rect 5784 2718 5840 2720
rect 5864 2718 5920 2720
rect 5944 2718 6000 2720
rect 6024 2718 6080 2720
rect 6104 2718 6160 2720
rect 5724 2234 5780 2236
rect 5804 2234 5860 2236
rect 5884 2234 5940 2236
rect 5964 2234 6020 2236
rect 6044 2234 6100 2236
rect 6124 2234 6180 2236
rect 5724 2182 5734 2234
rect 5734 2182 5780 2234
rect 5804 2182 5850 2234
rect 5850 2182 5860 2234
rect 5884 2182 5914 2234
rect 5914 2182 5926 2234
rect 5926 2182 5940 2234
rect 5964 2182 5978 2234
rect 5978 2182 5990 2234
rect 5990 2182 6020 2234
rect 6044 2182 6054 2234
rect 6054 2182 6100 2234
rect 6124 2182 6170 2234
rect 6170 2182 6180 2234
rect 5724 2180 5780 2182
rect 5804 2180 5860 2182
rect 5884 2180 5940 2182
rect 5964 2180 6020 2182
rect 6044 2180 6100 2182
rect 6124 2180 6180 2182
rect 144 1490 212 1558
rect 1374 1533 1430 1535
rect 1454 1533 1510 1535
rect 1534 1533 1590 1535
rect 1614 1533 1670 1535
rect 1694 1533 1750 1535
rect 1774 1533 1830 1535
rect 1854 1533 1910 1535
rect 1374 1481 1412 1533
rect 1412 1481 1424 1533
rect 1424 1481 1430 1533
rect 1454 1481 1476 1533
rect 1476 1481 1488 1533
rect 1488 1481 1510 1533
rect 1534 1481 1540 1533
rect 1540 1481 1552 1533
rect 1552 1481 1590 1533
rect 1614 1481 1616 1533
rect 1616 1481 1668 1533
rect 1668 1481 1670 1533
rect 1694 1481 1732 1533
rect 1732 1481 1744 1533
rect 1744 1481 1750 1533
rect 1774 1481 1796 1533
rect 1796 1481 1808 1533
rect 1808 1481 1830 1533
rect 1854 1481 1860 1533
rect 1860 1481 1872 1533
rect 1872 1481 1910 1533
rect 1374 1479 1430 1481
rect 1454 1479 1510 1481
rect 1534 1479 1590 1481
rect 1614 1479 1670 1481
rect 1694 1479 1750 1481
rect 1774 1479 1830 1481
rect 1854 1479 1910 1481
rect 3746 1544 3802 1546
rect 3826 1544 3882 1546
rect 3906 1544 3962 1546
rect 3986 1544 4042 1546
rect 4066 1544 4122 1546
rect 4146 1544 4202 1546
rect 3746 1492 3756 1544
rect 3756 1492 3802 1544
rect 3826 1492 3872 1544
rect 3872 1492 3882 1544
rect 3906 1492 3936 1544
rect 3936 1492 3948 1544
rect 3948 1492 3962 1544
rect 3986 1492 4000 1544
rect 4000 1492 4012 1544
rect 4012 1492 4042 1544
rect 4066 1492 4076 1544
rect 4076 1492 4122 1544
rect 4146 1492 4192 1544
rect 4192 1492 4202 1544
rect 3746 1490 3802 1492
rect 3826 1490 3882 1492
rect 3906 1490 3962 1492
rect 3986 1490 4042 1492
rect 4066 1490 4122 1492
rect 4146 1490 4202 1492
rect 1388 1007 1444 1009
rect 1468 1007 1524 1009
rect 1548 1007 1604 1009
rect 1628 1007 1684 1009
rect 1708 1007 1764 1009
rect 1788 1007 1844 1009
rect 1388 955 1398 1007
rect 1398 955 1444 1007
rect 1468 955 1514 1007
rect 1514 955 1524 1007
rect 1548 955 1578 1007
rect 1578 955 1590 1007
rect 1590 955 1604 1007
rect 1628 955 1642 1007
rect 1642 955 1654 1007
rect 1654 955 1684 1007
rect 1708 955 1718 1007
rect 1718 955 1764 1007
rect 1788 955 1834 1007
rect 1834 955 1844 1007
rect 1388 953 1444 955
rect 1468 953 1524 955
rect 1548 953 1604 955
rect 1628 953 1684 955
rect 1708 953 1764 955
rect 1788 953 1844 955
rect 1932 701 1988 702
rect 1932 649 1935 701
rect 1935 649 1987 701
rect 1987 649 1988 701
rect 1932 646 1988 649
rect 5704 1544 5760 1546
rect 5784 1544 5840 1546
rect 5864 1544 5920 1546
rect 5944 1544 6000 1546
rect 6024 1544 6080 1546
rect 6104 1544 6160 1546
rect 5704 1492 5714 1544
rect 5714 1492 5760 1544
rect 5784 1492 5830 1544
rect 5830 1492 5840 1544
rect 5864 1492 5894 1544
rect 5894 1492 5906 1544
rect 5906 1492 5920 1544
rect 5944 1492 5958 1544
rect 5958 1492 5970 1544
rect 5970 1492 6000 1544
rect 6024 1492 6034 1544
rect 6034 1492 6080 1544
rect 6104 1492 6150 1544
rect 6150 1492 6160 1544
rect 5704 1490 5760 1492
rect 5784 1490 5840 1492
rect 5864 1490 5920 1492
rect 5944 1490 6000 1492
rect 6024 1490 6080 1492
rect 6104 1490 6160 1492
rect 3766 1006 3822 1008
rect 3846 1006 3902 1008
rect 3926 1006 3982 1008
rect 4006 1006 4062 1008
rect 4086 1006 4142 1008
rect 4166 1006 4222 1008
rect 3766 954 3776 1006
rect 3776 954 3822 1006
rect 3846 954 3892 1006
rect 3892 954 3902 1006
rect 3926 954 3956 1006
rect 3956 954 3968 1006
rect 3968 954 3982 1006
rect 4006 954 4020 1006
rect 4020 954 4032 1006
rect 4032 954 4062 1006
rect 4086 954 4096 1006
rect 4096 954 4142 1006
rect 4166 954 4212 1006
rect 4212 954 4222 1006
rect 3766 952 3822 954
rect 3846 952 3902 954
rect 3926 952 3982 954
rect 4006 952 4062 954
rect 4086 952 4142 954
rect 4166 952 4222 954
rect 2520 488 2576 490
rect 2520 436 2522 488
rect 2522 436 2574 488
rect 2574 436 2576 488
rect 2520 434 2576 436
rect 144 254 212 322
rect 1374 305 1430 307
rect 1454 305 1510 307
rect 1534 305 1590 307
rect 1614 305 1670 307
rect 1694 305 1750 307
rect 1774 305 1830 307
rect 1854 305 1910 307
rect 1374 253 1412 305
rect 1412 253 1424 305
rect 1424 253 1430 305
rect 1454 253 1476 305
rect 1476 253 1488 305
rect 1488 253 1510 305
rect 1534 253 1540 305
rect 1540 253 1552 305
rect 1552 253 1590 305
rect 1614 253 1616 305
rect 1616 253 1668 305
rect 1668 253 1670 305
rect 1694 253 1732 305
rect 1732 253 1744 305
rect 1744 253 1750 305
rect 1774 253 1796 305
rect 1796 253 1808 305
rect 1808 253 1830 305
rect 1854 253 1860 305
rect 1860 253 1872 305
rect 1872 253 1910 305
rect 1374 251 1430 253
rect 1454 251 1510 253
rect 1534 251 1590 253
rect 1614 251 1670 253
rect 1694 251 1750 253
rect 1774 251 1830 253
rect 1854 251 1910 253
rect 3746 316 3802 318
rect 3826 316 3882 318
rect 3906 316 3962 318
rect 3986 316 4042 318
rect 4066 316 4122 318
rect 4146 316 4202 318
rect 3746 264 3756 316
rect 3756 264 3802 316
rect 3826 264 3872 316
rect 3872 264 3882 316
rect 3906 264 3936 316
rect 3936 264 3948 316
rect 3948 264 3962 316
rect 3986 264 4000 316
rect 4000 264 4012 316
rect 4012 264 4042 316
rect 4066 264 4076 316
rect 4076 264 4122 316
rect 4146 264 4192 316
rect 4192 264 4202 316
rect 3746 262 3802 264
rect 3826 262 3882 264
rect 3906 262 3962 264
rect 3986 262 4042 264
rect 4066 262 4122 264
rect 4146 262 4202 264
<< metal3 >>
rect -2 19429 7724 19470
rect -2 19426 1388 19429
rect -2 19358 42 19426
rect 110 19373 1388 19426
rect 1444 19373 1468 19429
rect 1524 19373 1548 19429
rect 1604 19373 1628 19429
rect 1684 19373 1708 19429
rect 1764 19373 1788 19429
rect 1844 19428 7724 19429
rect 1844 19373 3766 19428
rect 110 19372 3766 19373
rect 3822 19372 3846 19428
rect 3902 19372 3926 19428
rect 3982 19372 4006 19428
rect 4062 19372 4086 19428
rect 4142 19372 4166 19428
rect 4222 19372 5724 19428
rect 5780 19372 5804 19428
rect 5860 19372 5884 19428
rect 5940 19372 5964 19428
rect 6020 19372 6044 19428
rect 6100 19372 6124 19428
rect 6180 19372 7724 19428
rect 110 19358 7724 19372
rect -2 19330 7724 19358
rect 1925 19122 1995 19129
rect 1925 19066 1932 19122
rect 1988 19066 1995 19122
rect 1925 19059 1995 19066
rect 1930 18912 1990 19059
rect 2513 18912 2583 18917
rect 1930 18910 2583 18912
rect 1930 18854 2520 18910
rect 2576 18854 2583 18910
rect 1930 18852 2583 18854
rect 2513 18847 2583 18852
rect -2 18750 7724 18780
rect -2 18682 144 18750
rect 212 18738 7724 18750
rect 212 18727 3746 18738
rect 212 18682 1374 18727
rect -2 18671 1374 18682
rect 1430 18671 1454 18727
rect 1510 18671 1534 18727
rect 1590 18671 1614 18727
rect 1670 18671 1694 18727
rect 1750 18671 1774 18727
rect 1830 18671 1854 18727
rect 1910 18682 3746 18727
rect 3802 18682 3826 18738
rect 3882 18682 3906 18738
rect 3962 18682 3986 18738
rect 4042 18682 4066 18738
rect 4122 18682 4146 18738
rect 4202 18682 5704 18738
rect 5760 18682 5784 18738
rect 5840 18682 5864 18738
rect 5920 18682 5944 18738
rect 6000 18682 6024 18738
rect 6080 18682 6104 18738
rect 6160 18682 7724 18738
rect 1910 18671 7724 18682
rect -2 18640 7724 18671
rect -2 18220 7724 18242
rect -2 18152 42 18220
rect 110 18201 7724 18220
rect 110 18152 1388 18201
rect -2 18145 1388 18152
rect 1444 18145 1468 18201
rect 1524 18145 1548 18201
rect 1604 18145 1628 18201
rect 1684 18145 1708 18201
rect 1764 18145 1788 18201
rect 1844 18200 7724 18201
rect 1844 18145 3766 18200
rect -2 18144 3766 18145
rect 3822 18144 3846 18200
rect 3902 18144 3926 18200
rect 3982 18144 4006 18200
rect 4062 18144 4086 18200
rect 4142 18144 4166 18200
rect 4222 18144 5724 18200
rect 5780 18144 5804 18200
rect 5860 18144 5884 18200
rect 5940 18144 5964 18200
rect 6020 18144 6044 18200
rect 6100 18144 6124 18200
rect 6180 18144 7724 18200
rect -2 18102 7724 18144
rect 1925 17894 1995 17901
rect 1925 17838 1932 17894
rect 1988 17838 1995 17894
rect 1925 17831 1995 17838
rect 1930 17684 1990 17831
rect 2513 17684 2583 17689
rect 1930 17682 2583 17684
rect 1930 17626 2520 17682
rect 2576 17626 2583 17682
rect 1930 17624 2583 17626
rect 2513 17619 2583 17624
rect -2 17514 7724 17552
rect -2 17446 144 17514
rect 212 17510 7724 17514
rect 212 17499 3746 17510
rect 212 17446 1374 17499
rect -2 17443 1374 17446
rect 1430 17443 1454 17499
rect 1510 17443 1534 17499
rect 1590 17443 1614 17499
rect 1670 17443 1694 17499
rect 1750 17443 1774 17499
rect 1830 17443 1854 17499
rect 1910 17454 3746 17499
rect 3802 17454 3826 17510
rect 3882 17454 3906 17510
rect 3962 17454 3986 17510
rect 4042 17454 4066 17510
rect 4122 17454 4146 17510
rect 4202 17454 5704 17510
rect 5760 17454 5784 17510
rect 5840 17454 5864 17510
rect 5920 17454 5944 17510
rect 6000 17454 6024 17510
rect 6080 17454 6104 17510
rect 6160 17454 7724 17510
rect 1910 17443 7724 17454
rect -2 17412 7724 17443
rect -2 16973 7724 17014
rect -2 16970 1388 16973
rect -2 16902 42 16970
rect 110 16917 1388 16970
rect 1444 16917 1468 16973
rect 1524 16917 1548 16973
rect 1604 16917 1628 16973
rect 1684 16917 1708 16973
rect 1764 16917 1788 16973
rect 1844 16972 7724 16973
rect 1844 16917 3766 16972
rect 110 16916 3766 16917
rect 3822 16916 3846 16972
rect 3902 16916 3926 16972
rect 3982 16916 4006 16972
rect 4062 16916 4086 16972
rect 4142 16916 4166 16972
rect 4222 16916 5724 16972
rect 5780 16916 5804 16972
rect 5860 16916 5884 16972
rect 5940 16916 5964 16972
rect 6020 16916 6044 16972
rect 6100 16916 6124 16972
rect 6180 16916 7724 16972
rect 110 16902 7724 16916
rect -2 16874 7724 16902
rect 1925 16666 1995 16673
rect 1925 16610 1932 16666
rect 1988 16610 1995 16666
rect 1925 16603 1995 16610
rect 1930 16456 1990 16603
rect 2513 16456 2583 16461
rect 1930 16454 2583 16456
rect 1930 16398 2520 16454
rect 2576 16398 2583 16454
rect 1930 16396 2583 16398
rect 2513 16391 2583 16396
rect -2 16294 7724 16324
rect -2 16226 144 16294
rect 212 16282 7724 16294
rect 212 16271 3746 16282
rect 212 16226 1374 16271
rect -2 16215 1374 16226
rect 1430 16215 1454 16271
rect 1510 16215 1534 16271
rect 1590 16215 1614 16271
rect 1670 16215 1694 16271
rect 1750 16215 1774 16271
rect 1830 16215 1854 16271
rect 1910 16226 3746 16271
rect 3802 16226 3826 16282
rect 3882 16226 3906 16282
rect 3962 16226 3986 16282
rect 4042 16226 4066 16282
rect 4122 16226 4146 16282
rect 4202 16226 5704 16282
rect 5760 16226 5784 16282
rect 5840 16226 5864 16282
rect 5920 16226 5944 16282
rect 6000 16226 6024 16282
rect 6080 16226 6104 16282
rect 6160 16226 7724 16282
rect 1910 16215 7724 16226
rect -2 16184 7724 16215
rect -2 15764 7724 15786
rect -2 15696 42 15764
rect 110 15745 7724 15764
rect 110 15696 1388 15745
rect -2 15689 1388 15696
rect 1444 15689 1468 15745
rect 1524 15689 1548 15745
rect 1604 15689 1628 15745
rect 1684 15689 1708 15745
rect 1764 15689 1788 15745
rect 1844 15744 7724 15745
rect 1844 15689 3766 15744
rect -2 15688 3766 15689
rect 3822 15688 3846 15744
rect 3902 15688 3926 15744
rect 3982 15688 4006 15744
rect 4062 15688 4086 15744
rect 4142 15688 4166 15744
rect 4222 15688 5724 15744
rect 5780 15688 5804 15744
rect 5860 15688 5884 15744
rect 5940 15688 5964 15744
rect 6020 15688 6044 15744
rect 6100 15688 6124 15744
rect 6180 15688 7724 15744
rect -2 15646 7724 15688
rect 1925 15438 1995 15445
rect 1925 15382 1932 15438
rect 1988 15382 1995 15438
rect 1925 15375 1995 15382
rect 1930 15228 1990 15375
rect 2513 15228 2583 15233
rect 1930 15226 2583 15228
rect 1930 15170 2520 15226
rect 2576 15170 2583 15226
rect 1930 15168 2583 15170
rect 2513 15163 2583 15168
rect -2 15058 7724 15096
rect -2 14990 144 15058
rect 212 15054 7724 15058
rect 212 15043 3746 15054
rect 212 14990 1374 15043
rect -2 14987 1374 14990
rect 1430 14987 1454 15043
rect 1510 14987 1534 15043
rect 1590 14987 1614 15043
rect 1670 14987 1694 15043
rect 1750 14987 1774 15043
rect 1830 14987 1854 15043
rect 1910 14998 3746 15043
rect 3802 14998 3826 15054
rect 3882 14998 3906 15054
rect 3962 14998 3986 15054
rect 4042 14998 4066 15054
rect 4122 14998 4146 15054
rect 4202 14998 5704 15054
rect 5760 14998 5784 15054
rect 5840 14998 5864 15054
rect 5920 14998 5944 15054
rect 6000 14998 6024 15054
rect 6080 14998 6104 15054
rect 6160 14998 7724 15054
rect 1910 14987 7724 14998
rect -2 14956 7724 14987
rect -2 14517 7724 14558
rect -2 14514 1388 14517
rect -2 14446 42 14514
rect 110 14461 1388 14514
rect 1444 14461 1468 14517
rect 1524 14461 1548 14517
rect 1604 14461 1628 14517
rect 1684 14461 1708 14517
rect 1764 14461 1788 14517
rect 1844 14516 7724 14517
rect 1844 14461 3766 14516
rect 110 14460 3766 14461
rect 3822 14460 3846 14516
rect 3902 14460 3926 14516
rect 3982 14460 4006 14516
rect 4062 14460 4086 14516
rect 4142 14460 4166 14516
rect 4222 14460 5724 14516
rect 5780 14460 5804 14516
rect 5860 14460 5884 14516
rect 5940 14460 5964 14516
rect 6020 14460 6044 14516
rect 6100 14460 6124 14516
rect 6180 14460 7724 14516
rect 110 14446 7724 14460
rect -2 14418 7724 14446
rect 1925 14210 1995 14217
rect 1925 14154 1932 14210
rect 1988 14154 1995 14210
rect 1925 14147 1995 14154
rect 1930 14000 1990 14147
rect 2513 14000 2583 14005
rect 1930 13998 2583 14000
rect 1930 13942 2520 13998
rect 2576 13942 2583 13998
rect 1930 13940 2583 13942
rect 2513 13935 2583 13940
rect -2 13838 7724 13868
rect -2 13770 144 13838
rect 212 13826 7724 13838
rect 212 13815 3746 13826
rect 212 13770 1374 13815
rect -2 13759 1374 13770
rect 1430 13759 1454 13815
rect 1510 13759 1534 13815
rect 1590 13759 1614 13815
rect 1670 13759 1694 13815
rect 1750 13759 1774 13815
rect 1830 13759 1854 13815
rect 1910 13770 3746 13815
rect 3802 13770 3826 13826
rect 3882 13770 3906 13826
rect 3962 13770 3986 13826
rect 4042 13770 4066 13826
rect 4122 13770 4146 13826
rect 4202 13770 5704 13826
rect 5760 13770 5784 13826
rect 5840 13770 5864 13826
rect 5920 13770 5944 13826
rect 6000 13770 6024 13826
rect 6080 13770 6104 13826
rect 6160 13770 7724 13826
rect 1910 13759 7724 13770
rect -2 13728 7724 13759
rect -2 13308 7724 13330
rect -2 13240 42 13308
rect 110 13289 7724 13308
rect 110 13240 1388 13289
rect -2 13233 1388 13240
rect 1444 13233 1468 13289
rect 1524 13233 1548 13289
rect 1604 13233 1628 13289
rect 1684 13233 1708 13289
rect 1764 13233 1788 13289
rect 1844 13288 7724 13289
rect 1844 13233 3766 13288
rect -2 13232 3766 13233
rect 3822 13232 3846 13288
rect 3902 13232 3926 13288
rect 3982 13232 4006 13288
rect 4062 13232 4086 13288
rect 4142 13232 4166 13288
rect 4222 13232 5724 13288
rect 5780 13232 5804 13288
rect 5860 13232 5884 13288
rect 5940 13232 5964 13288
rect 6020 13232 6044 13288
rect 6100 13232 6124 13288
rect 6180 13232 7724 13288
rect -2 13190 7724 13232
rect 1925 12982 1995 12989
rect 1925 12926 1932 12982
rect 1988 12926 1995 12982
rect 1925 12919 1995 12926
rect 1930 12772 1990 12919
rect 2513 12772 2583 12777
rect 1930 12770 2583 12772
rect 1930 12714 2520 12770
rect 2576 12714 2583 12770
rect 1930 12712 2583 12714
rect 2513 12707 2583 12712
rect -2 12602 7724 12640
rect -2 12534 144 12602
rect 212 12598 7724 12602
rect 212 12587 3746 12598
rect 212 12534 1374 12587
rect -2 12531 1374 12534
rect 1430 12531 1454 12587
rect 1510 12531 1534 12587
rect 1590 12531 1614 12587
rect 1670 12531 1694 12587
rect 1750 12531 1774 12587
rect 1830 12531 1854 12587
rect 1910 12542 3746 12587
rect 3802 12542 3826 12598
rect 3882 12542 3906 12598
rect 3962 12542 3986 12598
rect 4042 12542 4066 12598
rect 4122 12542 4146 12598
rect 4202 12542 5704 12598
rect 5760 12542 5784 12598
rect 5840 12542 5864 12598
rect 5920 12542 5944 12598
rect 6000 12542 6024 12598
rect 6080 12542 6104 12598
rect 6160 12542 7724 12598
rect 1910 12531 7724 12542
rect -2 12500 7724 12531
rect -2 12061 7724 12102
rect -2 12058 1388 12061
rect -2 11990 42 12058
rect 110 12005 1388 12058
rect 1444 12005 1468 12061
rect 1524 12005 1548 12061
rect 1604 12005 1628 12061
rect 1684 12005 1708 12061
rect 1764 12005 1788 12061
rect 1844 12060 7724 12061
rect 1844 12005 3766 12060
rect 110 12004 3766 12005
rect 3822 12004 3846 12060
rect 3902 12004 3926 12060
rect 3982 12004 4006 12060
rect 4062 12004 4086 12060
rect 4142 12004 4166 12060
rect 4222 12004 5724 12060
rect 5780 12004 5804 12060
rect 5860 12004 5884 12060
rect 5940 12004 5964 12060
rect 6020 12004 6044 12060
rect 6100 12004 6124 12060
rect 6180 12004 7724 12060
rect 110 11990 7724 12004
rect -2 11962 7724 11990
rect 1925 11754 1995 11761
rect 1925 11698 1932 11754
rect 1988 11698 1995 11754
rect 1925 11691 1995 11698
rect 1930 11544 1990 11691
rect 2513 11544 2583 11549
rect 1930 11542 2583 11544
rect 1930 11486 2520 11542
rect 2576 11486 2583 11542
rect 1930 11484 2583 11486
rect 2513 11479 2583 11484
rect -2 11382 7724 11412
rect -2 11314 144 11382
rect 212 11370 7724 11382
rect 212 11359 3746 11370
rect 212 11314 1374 11359
rect -2 11303 1374 11314
rect 1430 11303 1454 11359
rect 1510 11303 1534 11359
rect 1590 11303 1614 11359
rect 1670 11303 1694 11359
rect 1750 11303 1774 11359
rect 1830 11303 1854 11359
rect 1910 11314 3746 11359
rect 3802 11314 3826 11370
rect 3882 11314 3906 11370
rect 3962 11314 3986 11370
rect 4042 11314 4066 11370
rect 4122 11314 4146 11370
rect 4202 11314 5704 11370
rect 5760 11314 5784 11370
rect 5840 11314 5864 11370
rect 5920 11314 5944 11370
rect 6000 11314 6024 11370
rect 6080 11314 6104 11370
rect 6160 11314 7724 11370
rect 1910 11303 7724 11314
rect -2 11272 7724 11303
rect -2 10852 7724 10874
rect -2 10784 42 10852
rect 110 10833 7724 10852
rect 110 10784 1388 10833
rect -2 10777 1388 10784
rect 1444 10777 1468 10833
rect 1524 10777 1548 10833
rect 1604 10777 1628 10833
rect 1684 10777 1708 10833
rect 1764 10777 1788 10833
rect 1844 10832 7724 10833
rect 1844 10777 3766 10832
rect -2 10776 3766 10777
rect 3822 10776 3846 10832
rect 3902 10776 3926 10832
rect 3982 10776 4006 10832
rect 4062 10776 4086 10832
rect 4142 10776 4166 10832
rect 4222 10776 5724 10832
rect 5780 10776 5804 10832
rect 5860 10776 5884 10832
rect 5940 10776 5964 10832
rect 6020 10776 6044 10832
rect 6100 10776 6124 10832
rect 6180 10776 7724 10832
rect -2 10734 7724 10776
rect 1925 10526 1995 10533
rect 1925 10470 1932 10526
rect 1988 10470 1995 10526
rect 1925 10463 1995 10470
rect 1930 10316 1990 10463
rect 2513 10316 2583 10321
rect 1930 10314 2583 10316
rect 1930 10258 2520 10314
rect 2576 10258 2583 10314
rect 1930 10256 2583 10258
rect 2513 10251 2583 10256
rect -2 10146 7724 10184
rect -2 10078 144 10146
rect 212 10142 7724 10146
rect 212 10131 3746 10142
rect 212 10078 1374 10131
rect -2 10075 1374 10078
rect 1430 10075 1454 10131
rect 1510 10075 1534 10131
rect 1590 10075 1614 10131
rect 1670 10075 1694 10131
rect 1750 10075 1774 10131
rect 1830 10075 1854 10131
rect 1910 10086 3746 10131
rect 3802 10086 3826 10142
rect 3882 10086 3906 10142
rect 3962 10086 3986 10142
rect 4042 10086 4066 10142
rect 4122 10086 4146 10142
rect 4202 10086 5704 10142
rect 5760 10086 5784 10142
rect 5840 10086 5864 10142
rect 5920 10086 5944 10142
rect 6000 10086 6024 10142
rect 6080 10086 6104 10142
rect 6160 10086 7724 10142
rect 1910 10075 7724 10086
rect -2 10044 7724 10075
rect -2 9605 7724 9646
rect -2 9602 1388 9605
rect -2 9534 42 9602
rect 110 9549 1388 9602
rect 1444 9549 1468 9605
rect 1524 9549 1548 9605
rect 1604 9549 1628 9605
rect 1684 9549 1708 9605
rect 1764 9549 1788 9605
rect 1844 9604 7724 9605
rect 1844 9549 3766 9604
rect 110 9548 3766 9549
rect 3822 9548 3846 9604
rect 3902 9548 3926 9604
rect 3982 9548 4006 9604
rect 4062 9548 4086 9604
rect 4142 9548 4166 9604
rect 4222 9548 5724 9604
rect 5780 9548 5804 9604
rect 5860 9548 5884 9604
rect 5940 9548 5964 9604
rect 6020 9548 6044 9604
rect 6100 9548 6124 9604
rect 6180 9548 7724 9604
rect 110 9534 7724 9548
rect -2 9506 7724 9534
rect 1925 9298 1995 9305
rect 1925 9242 1932 9298
rect 1988 9242 1995 9298
rect 1925 9235 1995 9242
rect 1930 9088 1990 9235
rect 2513 9088 2583 9093
rect 1930 9086 2583 9088
rect 1930 9030 2520 9086
rect 2576 9030 2583 9086
rect 1930 9028 2583 9030
rect 2513 9023 2583 9028
rect -2 8926 7724 8956
rect -2 8858 144 8926
rect 212 8914 7724 8926
rect 212 8903 3746 8914
rect 212 8858 1374 8903
rect -2 8847 1374 8858
rect 1430 8847 1454 8903
rect 1510 8847 1534 8903
rect 1590 8847 1614 8903
rect 1670 8847 1694 8903
rect 1750 8847 1774 8903
rect 1830 8847 1854 8903
rect 1910 8858 3746 8903
rect 3802 8858 3826 8914
rect 3882 8858 3906 8914
rect 3962 8858 3986 8914
rect 4042 8858 4066 8914
rect 4122 8858 4146 8914
rect 4202 8858 5704 8914
rect 5760 8858 5784 8914
rect 5840 8858 5864 8914
rect 5920 8858 5944 8914
rect 6000 8858 6024 8914
rect 6080 8858 6104 8914
rect 6160 8858 7724 8914
rect 1910 8847 7724 8858
rect -2 8816 7724 8847
rect -2 8396 7724 8418
rect -2 8328 42 8396
rect 110 8377 7724 8396
rect 110 8328 1388 8377
rect -2 8321 1388 8328
rect 1444 8321 1468 8377
rect 1524 8321 1548 8377
rect 1604 8321 1628 8377
rect 1684 8321 1708 8377
rect 1764 8321 1788 8377
rect 1844 8376 7724 8377
rect 1844 8321 3766 8376
rect -2 8320 3766 8321
rect 3822 8320 3846 8376
rect 3902 8320 3926 8376
rect 3982 8320 4006 8376
rect 4062 8320 4086 8376
rect 4142 8320 4166 8376
rect 4222 8320 5724 8376
rect 5780 8320 5804 8376
rect 5860 8320 5884 8376
rect 5940 8320 5964 8376
rect 6020 8320 6044 8376
rect 6100 8320 6124 8376
rect 6180 8320 7724 8376
rect -2 8278 7724 8320
rect 1925 8070 1995 8077
rect 1925 8014 1932 8070
rect 1988 8014 1995 8070
rect 1925 8007 1995 8014
rect 1930 7860 1990 8007
rect 2513 7860 2583 7865
rect 1930 7858 2583 7860
rect 1930 7802 2520 7858
rect 2576 7802 2583 7858
rect 1930 7800 2583 7802
rect 2513 7795 2583 7800
rect -2 7690 7724 7728
rect -2 7622 144 7690
rect 212 7686 7724 7690
rect 212 7675 3746 7686
rect 212 7622 1374 7675
rect -2 7619 1374 7622
rect 1430 7619 1454 7675
rect 1510 7619 1534 7675
rect 1590 7619 1614 7675
rect 1670 7619 1694 7675
rect 1750 7619 1774 7675
rect 1830 7619 1854 7675
rect 1910 7630 3746 7675
rect 3802 7630 3826 7686
rect 3882 7630 3906 7686
rect 3962 7630 3986 7686
rect 4042 7630 4066 7686
rect 4122 7630 4146 7686
rect 4202 7630 5704 7686
rect 5760 7630 5784 7686
rect 5840 7630 5864 7686
rect 5920 7630 5944 7686
rect 6000 7630 6024 7686
rect 6080 7630 6104 7686
rect 6160 7630 7724 7686
rect 1910 7619 7724 7630
rect -2 7588 7724 7619
rect -2 7149 7724 7190
rect -2 7146 1388 7149
rect -2 7078 42 7146
rect 110 7093 1388 7146
rect 1444 7093 1468 7149
rect 1524 7093 1548 7149
rect 1604 7093 1628 7149
rect 1684 7093 1708 7149
rect 1764 7093 1788 7149
rect 1844 7148 7724 7149
rect 1844 7093 3766 7148
rect 110 7092 3766 7093
rect 3822 7092 3846 7148
rect 3902 7092 3926 7148
rect 3982 7092 4006 7148
rect 4062 7092 4086 7148
rect 4142 7092 4166 7148
rect 4222 7092 5724 7148
rect 5780 7092 5804 7148
rect 5860 7092 5884 7148
rect 5940 7092 5964 7148
rect 6020 7092 6044 7148
rect 6100 7092 6124 7148
rect 6180 7092 7724 7148
rect 110 7078 7724 7092
rect -2 7050 7724 7078
rect 1925 6842 1995 6849
rect 1925 6786 1932 6842
rect 1988 6786 1995 6842
rect 1925 6779 1995 6786
rect 1930 6632 1990 6779
rect 2513 6632 2583 6637
rect 1930 6630 2583 6632
rect 1930 6574 2520 6630
rect 2576 6574 2583 6630
rect 1930 6572 2583 6574
rect 2513 6567 2583 6572
rect -2 6470 7724 6500
rect -2 6402 144 6470
rect 212 6458 7724 6470
rect 212 6447 3746 6458
rect 212 6402 1374 6447
rect -2 6391 1374 6402
rect 1430 6391 1454 6447
rect 1510 6391 1534 6447
rect 1590 6391 1614 6447
rect 1670 6391 1694 6447
rect 1750 6391 1774 6447
rect 1830 6391 1854 6447
rect 1910 6402 3746 6447
rect 3802 6402 3826 6458
rect 3882 6402 3906 6458
rect 3962 6402 3986 6458
rect 4042 6402 4066 6458
rect 4122 6402 4146 6458
rect 4202 6402 5704 6458
rect 5760 6402 5784 6458
rect 5840 6402 5864 6458
rect 5920 6402 5944 6458
rect 6000 6402 6024 6458
rect 6080 6402 6104 6458
rect 6160 6402 7724 6458
rect 1910 6391 7724 6402
rect -2 6360 7724 6391
rect -2 5940 7724 5962
rect -2 5872 42 5940
rect 110 5921 7724 5940
rect 110 5872 1388 5921
rect -2 5865 1388 5872
rect 1444 5865 1468 5921
rect 1524 5865 1548 5921
rect 1604 5865 1628 5921
rect 1684 5865 1708 5921
rect 1764 5865 1788 5921
rect 1844 5920 7724 5921
rect 1844 5865 3766 5920
rect -2 5864 3766 5865
rect 3822 5864 3846 5920
rect 3902 5864 3926 5920
rect 3982 5864 4006 5920
rect 4062 5864 4086 5920
rect 4142 5864 4166 5920
rect 4222 5864 5724 5920
rect 5780 5864 5804 5920
rect 5860 5864 5884 5920
rect 5940 5864 5964 5920
rect 6020 5864 6044 5920
rect 6100 5864 6124 5920
rect 6180 5864 7724 5920
rect -2 5822 7724 5864
rect 1925 5614 1995 5621
rect 1925 5558 1932 5614
rect 1988 5558 1995 5614
rect 1925 5551 1995 5558
rect 1930 5404 1990 5551
rect 2513 5404 2583 5409
rect 1930 5402 2583 5404
rect 1930 5346 2520 5402
rect 2576 5346 2583 5402
rect 1930 5344 2583 5346
rect 2513 5339 2583 5344
rect -2 5234 7724 5272
rect -2 5166 144 5234
rect 212 5230 7724 5234
rect 212 5219 3746 5230
rect 212 5166 1374 5219
rect -2 5163 1374 5166
rect 1430 5163 1454 5219
rect 1510 5163 1534 5219
rect 1590 5163 1614 5219
rect 1670 5163 1694 5219
rect 1750 5163 1774 5219
rect 1830 5163 1854 5219
rect 1910 5174 3746 5219
rect 3802 5174 3826 5230
rect 3882 5174 3906 5230
rect 3962 5174 3986 5230
rect 4042 5174 4066 5230
rect 4122 5174 4146 5230
rect 4202 5174 5704 5230
rect 5760 5174 5784 5230
rect 5840 5174 5864 5230
rect 5920 5174 5944 5230
rect 6000 5174 6024 5230
rect 6080 5174 6104 5230
rect 6160 5174 7724 5230
rect 1910 5163 7724 5174
rect -2 5132 7724 5163
rect -2 4693 7724 4734
rect -2 4690 1388 4693
rect -2 4622 42 4690
rect 110 4637 1388 4690
rect 1444 4637 1468 4693
rect 1524 4637 1548 4693
rect 1604 4637 1628 4693
rect 1684 4637 1708 4693
rect 1764 4637 1788 4693
rect 1844 4692 7724 4693
rect 1844 4637 3766 4692
rect 110 4636 3766 4637
rect 3822 4636 3846 4692
rect 3902 4636 3926 4692
rect 3982 4636 4006 4692
rect 4062 4636 4086 4692
rect 4142 4636 4166 4692
rect 4222 4636 5724 4692
rect 5780 4636 5804 4692
rect 5860 4636 5884 4692
rect 5940 4636 5964 4692
rect 6020 4636 6044 4692
rect 6100 4636 6124 4692
rect 6180 4636 7724 4692
rect 110 4622 7724 4636
rect -2 4594 7724 4622
rect 1925 4386 1995 4393
rect 1925 4330 1932 4386
rect 1988 4330 1995 4386
rect 1925 4323 1995 4330
rect 1930 4176 1990 4323
rect 2513 4176 2583 4181
rect 1930 4174 2583 4176
rect 1930 4118 2520 4174
rect 2576 4118 2583 4174
rect 1930 4116 2583 4118
rect 2513 4111 2583 4116
rect -2 4014 7724 4044
rect -2 3946 144 4014
rect 212 4002 7724 4014
rect 212 3991 3746 4002
rect 212 3946 1374 3991
rect -2 3935 1374 3946
rect 1430 3935 1454 3991
rect 1510 3935 1534 3991
rect 1590 3935 1614 3991
rect 1670 3935 1694 3991
rect 1750 3935 1774 3991
rect 1830 3935 1854 3991
rect 1910 3946 3746 3991
rect 3802 3946 3826 4002
rect 3882 3946 3906 4002
rect 3962 3946 3986 4002
rect 4042 3946 4066 4002
rect 4122 3946 4146 4002
rect 4202 3946 5704 4002
rect 5760 3946 5784 4002
rect 5840 3946 5864 4002
rect 5920 3946 5944 4002
rect 6000 3946 6024 4002
rect 6080 3946 6104 4002
rect 6160 3946 7724 4002
rect 1910 3935 7724 3946
rect -2 3904 7724 3935
rect -2 3484 7724 3506
rect -2 3416 42 3484
rect 110 3465 7724 3484
rect 110 3416 1388 3465
rect -2 3409 1388 3416
rect 1444 3409 1468 3465
rect 1524 3409 1548 3465
rect 1604 3409 1628 3465
rect 1684 3409 1708 3465
rect 1764 3409 1788 3465
rect 1844 3464 7724 3465
rect 1844 3409 3766 3464
rect -2 3408 3766 3409
rect 3822 3408 3846 3464
rect 3902 3408 3926 3464
rect 3982 3408 4006 3464
rect 4062 3408 4086 3464
rect 4142 3408 4166 3464
rect 4222 3408 5724 3464
rect 5780 3408 5804 3464
rect 5860 3408 5884 3464
rect 5940 3408 5964 3464
rect 6020 3408 6044 3464
rect 6100 3408 6124 3464
rect 6180 3408 7724 3464
rect -2 3366 7724 3408
rect 1925 3158 1995 3165
rect 1925 3102 1932 3158
rect 1988 3102 1995 3158
rect 1925 3095 1995 3102
rect 1930 2948 1990 3095
rect 2513 2948 2583 2953
rect 1930 2946 2583 2948
rect 1930 2890 2520 2946
rect 2576 2890 2583 2946
rect 1930 2888 2583 2890
rect 2513 2883 2583 2888
rect -2 2778 7724 2816
rect -2 2710 144 2778
rect 212 2774 7724 2778
rect 212 2763 3746 2774
rect 212 2710 1374 2763
rect -2 2707 1374 2710
rect 1430 2707 1454 2763
rect 1510 2707 1534 2763
rect 1590 2707 1614 2763
rect 1670 2707 1694 2763
rect 1750 2707 1774 2763
rect 1830 2707 1854 2763
rect 1910 2718 3746 2763
rect 3802 2718 3826 2774
rect 3882 2718 3906 2774
rect 3962 2718 3986 2774
rect 4042 2718 4066 2774
rect 4122 2718 4146 2774
rect 4202 2718 5704 2774
rect 5760 2718 5784 2774
rect 5840 2718 5864 2774
rect 5920 2718 5944 2774
rect 6000 2718 6024 2774
rect 6080 2718 6104 2774
rect 6160 2718 7724 2774
rect 1910 2707 7724 2718
rect -2 2676 7724 2707
rect -2 2237 7724 2278
rect -2 2234 1388 2237
rect -2 2166 42 2234
rect 110 2181 1388 2234
rect 1444 2181 1468 2237
rect 1524 2181 1548 2237
rect 1604 2181 1628 2237
rect 1684 2181 1708 2237
rect 1764 2181 1788 2237
rect 1844 2236 7724 2237
rect 1844 2181 3766 2236
rect 110 2180 3766 2181
rect 3822 2180 3846 2236
rect 3902 2180 3926 2236
rect 3982 2180 4006 2236
rect 4062 2180 4086 2236
rect 4142 2180 4166 2236
rect 4222 2180 5724 2236
rect 5780 2180 5804 2236
rect 5860 2180 5884 2236
rect 5940 2180 5964 2236
rect 6020 2180 6044 2236
rect 6100 2180 6124 2236
rect 6180 2180 7724 2236
rect 110 2166 7724 2180
rect -2 2138 7724 2166
rect 1925 1930 1995 1937
rect 1925 1874 1932 1930
rect 1988 1874 1995 1930
rect 1925 1867 1995 1874
rect 1930 1720 1990 1867
rect 2513 1720 2583 1725
rect 1930 1718 2583 1720
rect 1930 1662 2520 1718
rect 2576 1662 2583 1718
rect 1930 1660 2583 1662
rect 2513 1655 2583 1660
rect -2 1558 7724 1588
rect -2 1490 144 1558
rect 212 1546 7724 1558
rect 212 1535 3746 1546
rect 212 1490 1374 1535
rect -2 1479 1374 1490
rect 1430 1479 1454 1535
rect 1510 1479 1534 1535
rect 1590 1479 1614 1535
rect 1670 1479 1694 1535
rect 1750 1479 1774 1535
rect 1830 1479 1854 1535
rect 1910 1490 3746 1535
rect 3802 1490 3826 1546
rect 3882 1490 3906 1546
rect 3962 1490 3986 1546
rect 4042 1490 4066 1546
rect 4122 1490 4146 1546
rect 4202 1490 5704 1546
rect 5760 1490 5784 1546
rect 5840 1490 5864 1546
rect 5920 1490 5944 1546
rect 6000 1490 6024 1546
rect 6080 1490 6104 1546
rect 6160 1490 7724 1546
rect 1910 1479 7724 1490
rect -2 1448 7724 1479
rect -2 1028 7724 1050
rect -2 960 42 1028
rect 110 1009 7724 1028
rect 110 960 1388 1009
rect -2 953 1388 960
rect 1444 953 1468 1009
rect 1524 953 1548 1009
rect 1604 953 1628 1009
rect 1684 953 1708 1009
rect 1764 953 1788 1009
rect 1844 1008 7724 1009
rect 1844 953 3766 1008
rect -2 952 3766 953
rect 3822 952 3846 1008
rect 3902 952 3926 1008
rect 3982 952 4006 1008
rect 4062 952 4086 1008
rect 4142 952 4166 1008
rect 4222 952 7724 1008
rect -2 910 7724 952
rect 1925 702 1995 709
rect 1925 646 1932 702
rect 1988 646 1995 702
rect 1925 639 1995 646
rect 1930 492 1990 639
rect 2513 492 2583 497
rect 1930 490 2583 492
rect 1930 434 2520 490
rect 2576 434 2583 490
rect 1930 432 2583 434
rect 2513 427 2583 432
rect -2 322 7724 360
rect -2 254 144 322
rect 212 318 7724 322
rect 212 307 3746 318
rect 212 254 1374 307
rect -2 251 1374 254
rect 1430 251 1454 307
rect 1510 251 1534 307
rect 1590 251 1614 307
rect 1670 251 1694 307
rect 1750 251 1774 307
rect 1830 251 1854 307
rect 1910 262 3746 307
rect 3802 262 3826 318
rect 3882 262 3906 318
rect 3962 262 3986 318
rect 4042 262 4066 318
rect 4122 262 4146 318
rect 4202 262 7724 318
rect 1910 251 7724 262
rect -2 220 7724 251
<< labels >>
rlabel metal2 82 9906 82 9906 3 VCC
port 1 e
rlabel metal2 180 9904 180 9904 3 VSS
port 2 e
rlabel metal2 290 19592 290 19592 3 D0
port 3 e
rlabel metal2 392 19600 392 19600 3 VREFL
port 4 e
rlabel metal2 3576 19606 3576 19606 3 D1
port 5 e
rlabel metal2 5136 19622 5136 19622 3 D2
port 6 e
rlabel metal2 5230 19628 5230 19628 3 D3
port 7 e
rlabel metal2 5310 19634 5310 19634 3 D4
port 8 e
rlabel metal2 5386 19634 5386 19634 3 D5
port 9 e
rlabel metal2 282 42 282 42 3 D0_BUF
port 10 e
rlabel metal2 418 36 418 36 3 VREFH
port 11 e
rlabel metal2 3588 24 3588 24 3 D1_BUF
port 12 e
rlabel metal2 5128 1298 5128 1298 3 D2_BUF
port 13 e
rlabel metal2 5210 1312 5210 1312 3 D3_BUF
port 14 e
rlabel metal2 5288 1292 5288 1292 3 D4_BUF
port 15 e
rlabel metal2 5374 1294 5374 1294 3 D5_BUF
port 16 e
rlabel metal2 7344 10781 7344 10781 3 VOUT
port 17 e
flabel metal1 5562 10400 5582 10438 7 FreeSans 600 0 0 0 switch_n_3v3_0.DX
flabel metal1 5534 9946 5562 9984 7 FreeSans 600 0 0 0 switch_n_3v3_0.DX_BUF
flabel metal3 7052 10734 7082 10874 3 FreeSans 600 0 0 0 switch_n_3v3_0.VCC
flabel metal3 7052 10044 7082 10184 3 FreeSans 600 0 0 0 switch_n_3v3_0.VSS
flabel metal3 5072 10044 5102 10184 7 FreeSans 600 0 0 0 switch_n_3v3_0.VSS
flabel metal3 5072 10734 5102 10874 7 FreeSans 600 0 0 0 switch_n_3v3_0.VCC
flabel metal2 5142 10950 5142 10950 1 FreeSans 400 0 0 0 switch_n_3v3_0.D2
flabel metal2 5222 10954 5222 10954 1 FreeSans 400 0 0 0 switch_n_3v3_0.D3
flabel metal2 5304 10954 5304 10954 1 FreeSans 400 0 0 0 switch_n_3v3_0.D4
flabel metal2 5384 10956 5384 10956 1 FreeSans 400 0 0 0 switch_n_3v3_0.D5
flabel metal2 5462 10956 5462 10956 1 FreeSans 400 0 0 0 switch_n_3v3_0.D6
flabel metal2 5542 10954 5542 10954 1 FreeSans 400 0 0 0 switch_n_3v3_0.D7
flabel metal1 6516 10898 6556 10922 3 FreeSans 600 0 0 0 switch_n_3v3_0.VOUT
flabel metal2 6518 9976 6556 10000 7 FreeSans 600 0 0 0 switch_n_3v3_0.VOUT
flabel metal1 5872 10374 5872 10374 7 FreeSans 600 0 0 0 switch_n_3v3_0.DX_
flabel metal1 6908 9970 6936 9994 3 FreeSans 600 0 0 0 switch_n_3v3_0.VREFH
flabel metal1 6986 10894 7016 10914 3 FreeSans 600 0 0 0 switch_n_3v3_0.VREFL
rlabel metal2 72 4824 72 4824 7 5_bit_dac_0[0].VCC
rlabel metal2 170 4830 170 4830 7 5_bit_dac_0[0].VSS
rlabel metal2 308 9780 308 9780 7 5_bit_dac_0[0].D0
rlabel metal2 416 9768 416 9768 7 5_bit_dac_0[0].VREFL
rlabel metal2 312 44 312 44 7 5_bit_dac_0[0].D0_BUF
rlabel metal2 402 34 402 34 7 5_bit_dac_0[0].VREFH
rlabel metal2 3574 22 3574 22 7 5_bit_dac_0[0].D1_BUF
rlabel metal2 3586 9790 3586 9790 7 5_bit_dac_0[0].D1
rlabel metal2 5150 9800 5150 9800 7 5_bit_dac_0[0].D2
rlabel metal2 5222 9798 5222 9798 7 5_bit_dac_0[0].D3
rlabel metal2 5302 9806 5302 9806 7 5_bit_dac_0[0].D4
rlabel metal2 5152 1296 5152 1296 3 5_bit_dac_0[0].D2_BUF
rlabel metal2 5220 1306 5220 1306 3 5_bit_dac_0[0].D3_BUF
rlabel metal2 5294 1284 5294 1284 3 5_bit_dac_0[0].D4_BUF
rlabel metal2 7176 5084 7176 5084 3 5_bit_dac_0[0].VOUT
flabel metal1 5562 5488 5582 5526 7 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.DX
flabel metal1 5534 5034 5562 5072 7 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.DX_BUF
flabel metal3 7052 5822 7082 5962 3 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VCC
flabel metal3 7052 5132 7082 5272 3 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VSS
flabel metal3 5072 5132 5102 5272 7 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VSS
flabel metal3 5072 5822 5102 5962 7 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VCC
flabel metal2 5142 6038 5142 6038 1 FreeSans 400 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.D2
flabel metal2 5222 6042 5222 6042 1 FreeSans 400 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.D3
flabel metal2 5304 6042 5304 6042 1 FreeSans 400 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.D4
flabel metal2 5384 6044 5384 6044 1 FreeSans 400 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.D5
flabel metal2 5462 6044 5462 6044 1 FreeSans 400 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.D6
flabel metal2 5542 6042 5542 6042 1 FreeSans 400 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.D7
flabel metal1 6516 5986 6556 6010 3 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VOUT
flabel metal2 6518 5064 6556 5088 7 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VOUT
flabel metal1 5872 5462 5872 5462 7 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.DX_
flabel metal1 6908 5058 6936 5082 3 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VREFH
flabel metal1 6986 5982 7016 6002 3 FreeSans 600 0 0 0 5_bit_dac_0[0].switch_n_3v3_0.VREFL
rlabel metal2 74 4472 74 4472 7 5_bit_dac_0[0].4_bit_dac_0[0].VCC
rlabel metal2 182 3754 182 3754 7 5_bit_dac_0[0].4_bit_dac_0[0].VSS
rlabel metal2 312 4878 312 4878 7 5_bit_dac_0[0].4_bit_dac_0[0].D0
rlabel metal2 420 4878 420 4878 7 5_bit_dac_0[0].4_bit_dac_0[0].VREFL
rlabel metal2 316 22 316 22 7 5_bit_dac_0[0].4_bit_dac_0[0].D0_BUF
rlabel metal2 416 16 416 16 3 5_bit_dac_0[0].4_bit_dac_0[0].VREFH
rlabel metal2 3592 4898 3592 4898 3 5_bit_dac_0[0].4_bit_dac_0[0].D1
rlabel metal2 3574 8 3574 8 3 5_bit_dac_0[0].4_bit_dac_0[0].D1_BUF
rlabel metal2 5150 4900 5150 4900 3 5_bit_dac_0[0].4_bit_dac_0[0].D2
rlabel metal2 5222 4898 5222 4898 3 5_bit_dac_0[0].4_bit_dac_0[0].D3
rlabel metal2 5140 1282 5140 1282 3 5_bit_dac_0[0].4_bit_dac_0[0].D2_BUF
rlabel metal2 5212 1290 5212 1290 3 5_bit_dac_0[0].4_bit_dac_0[0].D3_BUF
rlabel metal2 7142 3534 7142 3534 3 5_bit_dac_0[0].4_bit_dac_0[0].VOUT
flabel metal1 5562 3032 5582 3070 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX
flabel metal1 5534 2578 5562 2616 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_BUF
flabel metal3 7052 3366 7082 3506 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VCC
flabel metal3 7052 2676 7082 2816 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VSS
flabel metal3 5072 2676 5102 2816 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VSS
flabel metal3 5072 3366 5102 3506 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VCC
flabel metal2 5142 3582 5142 3582 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2
flabel metal2 5222 3586 5222 3586 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D3
flabel metal2 5304 3586 5304 3586 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D4
flabel metal2 5384 3588 5384 3588 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D5
flabel metal2 5462 3588 5462 3588 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D6
flabel metal2 5542 3586 5542 3586 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D7
flabel metal1 6516 3530 6556 3554 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VOUT
flabel metal2 6518 2608 6556 2632 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VOUT
flabel metal1 5872 3006 5872 3006 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_
flabel metal1 6908 2602 6936 2626 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VREFH
flabel metal1 6986 3526 7016 3546 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.VREFL
rlabel metal3 18 2234 18 2234 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VCC
rlabel metal3 26 1522 26 1522 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VSS
rlabel metal2 302 2430 302 2430 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0
rlabel metal2 406 2432 406 2432 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VREFL
rlabel metal2 304 20 304 20 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0_BUF
rlabel metal2 400 12 400 12 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VREFH
rlabel metal2 3586 2450 3586 2450 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1
rlabel metal2 3586 12 3586 12 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1_BUF
rlabel metal2 5141 2436 5141 2436 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D2
rlabel metal2 5141 1290 5141 1290 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D2_BUF
rlabel metal2 7139 2310 7139 2310 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT
flabel metal1 5562 1804 5582 1842 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX
flabel metal1 5534 1350 5562 1388 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_BUF
flabel metal3 7052 2138 7082 2278 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal3 7052 1448 7082 1588 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 1448 5102 1588 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 2138 5102 2278 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal2 5142 2354 5142 2354 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D2
flabel metal2 5222 2358 5222 2358 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D3
flabel metal2 5304 2358 5304 2358 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D4
flabel metal2 5384 2360 5384 2360 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D5
flabel metal2 5462 2360 5462 2360 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D6
flabel metal2 5542 2358 5542 2358 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D7
flabel metal1 6516 2302 6556 2326 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal2 6518 1380 6556 1404 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal1 5872 1778 5872 1778 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_
flabel metal1 6908 1374 6936 1398 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VREFH
flabel metal1 6986 2298 7016 2318 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VREFL
rlabel metal3 148 991 148 991 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VCC
rlabel metal3 166 286 166 286 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VSS
rlabel metal2 295 1186 295 1186 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0
rlabel metal2 406 1186 406 1186 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VREFL
rlabel metal2 301 36 301 36 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 19 409 19 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VREFH
rlabel metal2 5056 1077 5056 1077 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT
rlabel metal2 3586 18 3586 18 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 1204 3584 1204 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1
flabel metal1 3492 966 3492 966 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 252 3478 252 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 662 1254 662 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 930 2662 930 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 756 1266 756 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 578 624 578 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 464 614 464 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 902 634 902 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 220 528 360 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 910 528 1050 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 575 3624 614 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 121 3603 160 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 910 5124 1050 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 220 5124 360 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 1074 4597 1099 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 151 4598 175 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 550 3914 550 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 220 3462 360 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 910 3462 1050 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 1107 4888 1107 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 141 5041 141 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 2219 148 2219 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VCC
rlabel metal3 166 1514 166 1514 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VSS
rlabel metal2 295 2414 295 2414 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D0
rlabel metal2 406 2414 406 2414 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFL
rlabel metal2 301 1264 301 1264 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 1247 409 1247 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH
rlabel metal2 5056 2305 5056 2305 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT
rlabel metal2 3586 1246 3586 1246 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 2432 3584 2432 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D1
flabel metal1 3492 2194 3492 2194 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 1480 3478 1480 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 1890 1254 1890 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 2158 2662 2158 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 1984 1266 1984 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 1806 624 1806 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 1692 614 1692 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 2130 634 2130 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 1448 528 1588 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 2138 528 2278 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 1803 3624 1842 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 1349 3603 1388 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 2138 5124 2278 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 1448 5124 1588 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 2302 4597 2327 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 1379 4598 1403 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 1778 3914 1778 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 1448 3462 1588 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 2138 3462 2278 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 2335 4888 2335 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 1369 5041 1369 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal3 18 4690 18 4690 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VCC
rlabel metal3 26 3978 26 3978 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VSS
rlabel metal2 302 4886 302 4886 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].D0
rlabel metal2 406 4888 406 4888 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFL
rlabel metal2 304 2476 304 2476 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].D0_BUF
rlabel metal2 400 2468 400 2468 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH
rlabel metal2 3586 4906 3586 4906 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].D1
rlabel metal2 3586 2468 3586 2468 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].D1_BUF
rlabel metal2 5141 4892 5141 4892 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].D2
rlabel metal2 5141 3746 5141 3746 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].D2_BUF
rlabel metal2 7139 4766 7139 4766 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT
flabel metal1 5562 4260 5582 4298 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX
flabel metal1 5534 3806 5562 3844 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_BUF
flabel metal3 7052 4594 7082 4734 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal3 7052 3904 7082 4044 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 3904 5102 4044 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 4594 5102 4734 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal2 5142 4810 5142 4810 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D2
flabel metal2 5222 4814 5222 4814 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D3
flabel metal2 5304 4814 5304 4814 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D4
flabel metal2 5384 4816 5384 4816 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D5
flabel metal2 5462 4816 5462 4816 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D6
flabel metal2 5542 4814 5542 4814 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D7
flabel metal1 6516 4758 6556 4782 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal2 6518 3836 6556 3860 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal1 5872 4234 5872 4234 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_
flabel metal1 6908 3830 6936 3854 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VREFH
flabel metal1 6986 4754 7016 4774 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VREFL
rlabel metal3 148 3447 148 3447 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VCC
rlabel metal3 166 2742 166 2742 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VSS
rlabel metal2 295 3642 295 3642 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0
rlabel metal2 406 3642 406 3642 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VREFL
rlabel metal2 301 2492 301 2492 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 2475 409 2475 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VREFH
rlabel metal2 5056 3533 5056 3533 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT
rlabel metal2 3586 2474 3586 2474 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 3660 3584 3660 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1
flabel metal1 3492 3422 3492 3422 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 2708 3478 2708 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 3118 1254 3118 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 3386 2662 3386 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 3212 1266 3212 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 3034 624 3034 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 2920 614 2920 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 3358 634 3358 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 2676 528 2816 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 3366 528 3506 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 3031 3624 3070 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 2577 3603 2616 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 3366 5124 3506 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 2676 5124 2816 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 3530 4597 3555 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 2607 4598 2631 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 3006 3914 3006 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 2676 3462 2816 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 3366 3462 3506 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 3563 4888 3563 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 2597 5041 2597 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 4675 148 4675 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VCC
rlabel metal3 166 3970 166 3970 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VSS
rlabel metal2 295 4870 295 4870 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D0
rlabel metal2 406 4870 406 4870 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFL
rlabel metal2 301 3720 301 3720 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 3703 409 3703 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH
rlabel metal2 5056 4761 5056 4761 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT
rlabel metal2 3586 3702 3586 3702 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 4888 3584 4888 7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D1
flabel metal1 3492 4650 3492 4650 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 3936 3478 3936 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 4346 1254 4346 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 4614 2662 4614 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 4440 1266 4440 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 4262 624 4262 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 4148 614 4148 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 4586 634 4586 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 3904 528 4044 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 4594 528 4734 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 4259 3624 4298 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 3805 3603 3844 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 4594 5124 4734 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 3904 5124 4044 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 4758 4597 4783 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 3835 4598 3859 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 4234 3914 4234 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 3904 3462 4044 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 4594 3462 4734 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 4791 4888 4791 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 3825 5041 3825 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal2 74 9384 74 9384 7 5_bit_dac_0[0].4_bit_dac_0[1].VCC
rlabel metal2 182 8666 182 8666 7 5_bit_dac_0[0].4_bit_dac_0[1].VSS
rlabel metal2 312 9790 312 9790 7 5_bit_dac_0[0].4_bit_dac_0[1].D0
rlabel metal2 420 9790 420 9790 7 5_bit_dac_0[0].4_bit_dac_0[1].VREFL
rlabel metal2 316 4934 316 4934 7 5_bit_dac_0[0].4_bit_dac_0[1].D0_BUF
rlabel metal2 416 4928 416 4928 3 5_bit_dac_0[0].4_bit_dac_0[1].VREFH
rlabel metal2 3592 9810 3592 9810 3 5_bit_dac_0[0].4_bit_dac_0[1].D1
rlabel metal2 3574 4920 3574 4920 3 5_bit_dac_0[0].4_bit_dac_0[1].D1_BUF
rlabel metal2 5150 9812 5150 9812 3 5_bit_dac_0[0].4_bit_dac_0[1].D2
rlabel metal2 5222 9810 5222 9810 3 5_bit_dac_0[0].4_bit_dac_0[1].D3
rlabel metal2 5140 6194 5140 6194 3 5_bit_dac_0[0].4_bit_dac_0[1].D2_BUF
rlabel metal2 5212 6202 5212 6202 3 5_bit_dac_0[0].4_bit_dac_0[1].D3_BUF
rlabel metal2 7142 8446 7142 8446 3 5_bit_dac_0[0].4_bit_dac_0[1].VOUT
flabel metal1 5562 7944 5582 7982 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX
flabel metal1 5534 7490 5562 7528 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_BUF
flabel metal3 7052 8278 7082 8418 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VCC
flabel metal3 7052 7588 7082 7728 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VSS
flabel metal3 5072 7588 5102 7728 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VSS
flabel metal3 5072 8278 5102 8418 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VCC
flabel metal2 5142 8494 5142 8494 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2
flabel metal2 5222 8498 5222 8498 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D3
flabel metal2 5304 8498 5304 8498 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D4
flabel metal2 5384 8500 5384 8500 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D5
flabel metal2 5462 8500 5462 8500 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D6
flabel metal2 5542 8498 5542 8498 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D7
flabel metal1 6516 8442 6556 8466 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VOUT
flabel metal2 6518 7520 6556 7544 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VOUT
flabel metal1 5872 7918 5872 7918 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_
flabel metal1 6908 7514 6936 7538 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VREFH
flabel metal1 6986 8438 7016 8458 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.VREFL
rlabel metal3 18 7146 18 7146 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VCC
rlabel metal3 26 6434 26 6434 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VSS
rlabel metal2 302 7342 302 7342 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0
rlabel metal2 406 7344 406 7344 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VREFL
rlabel metal2 304 4932 304 4932 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0_BUF
rlabel metal2 400 4924 400 4924 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VREFH
rlabel metal2 3586 7362 3586 7362 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1
rlabel metal2 3586 4924 3586 4924 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1_BUF
rlabel metal2 5141 7348 5141 7348 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D2
rlabel metal2 5141 6202 5141 6202 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D2_BUF
rlabel metal2 7139 7222 7139 7222 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT
flabel metal1 5562 6716 5582 6754 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX
flabel metal1 5534 6262 5562 6300 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_BUF
flabel metal3 7052 7050 7082 7190 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal3 7052 6360 7082 6500 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 6360 5102 6500 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 7050 5102 7190 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal2 5142 7266 5142 7266 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D2
flabel metal2 5222 7270 5222 7270 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D3
flabel metal2 5304 7270 5304 7270 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D4
flabel metal2 5384 7272 5384 7272 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D5
flabel metal2 5462 7272 5462 7272 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D6
flabel metal2 5542 7270 5542 7270 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D7
flabel metal1 6516 7214 6556 7238 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal2 6518 6292 6556 6316 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal1 5872 6690 5872 6690 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_
flabel metal1 6908 6286 6936 6310 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VREFH
flabel metal1 6986 7210 7016 7230 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VREFL
rlabel metal3 148 5903 148 5903 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VCC
rlabel metal3 166 5198 166 5198 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VSS
rlabel metal2 295 6098 295 6098 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0
rlabel metal2 406 6098 406 6098 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VREFL
rlabel metal2 301 4948 301 4948 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 4931 409 4931 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VREFH
rlabel metal2 5056 5989 5056 5989 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT
rlabel metal2 3586 4930 3586 4930 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 6116 3584 6116 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1
flabel metal1 3492 5878 3492 5878 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 5164 3478 5164 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 5574 1254 5574 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 5842 2662 5842 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 5668 1266 5668 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 5490 624 5490 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 5376 614 5376 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 5814 634 5814 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 5132 528 5272 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 5822 528 5962 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 5487 3624 5526 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 5033 3603 5072 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 5822 5124 5962 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 5132 5124 5272 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 5986 4597 6011 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 5063 4598 5087 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 5462 3914 5462 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 5132 3462 5272 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 5822 3462 5962 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 6019 4888 6019 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 5053 5041 5053 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 7131 148 7131 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VCC
rlabel metal3 166 6426 166 6426 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VSS
rlabel metal2 295 7326 295 7326 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D0
rlabel metal2 406 7326 406 7326 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFL
rlabel metal2 301 6176 301 6176 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 6159 409 6159 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH
rlabel metal2 5056 7217 5056 7217 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT
rlabel metal2 3586 6158 3586 6158 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 7344 3584 7344 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D1
flabel metal1 3492 7106 3492 7106 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 6392 3478 6392 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 6802 1254 6802 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 7070 2662 7070 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 6896 1266 6896 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 6718 624 6718 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 6604 614 6604 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 7042 634 7042 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 6360 528 6500 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 7050 528 7190 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 6715 3624 6754 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 6261 3603 6300 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 7050 5124 7190 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 6360 5124 6500 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 7214 4597 7239 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 6291 4598 6315 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 6690 3914 6690 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 6360 3462 6500 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 7050 3462 7190 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 7247 4888 7247 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 6281 5041 6281 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal3 18 9602 18 9602 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VCC
rlabel metal3 26 8890 26 8890 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VSS
rlabel metal2 302 9798 302 9798 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].D0
rlabel metal2 406 9800 406 9800 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFL
rlabel metal2 304 7388 304 7388 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].D0_BUF
rlabel metal2 400 7380 400 7380 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH
rlabel metal2 3586 9818 3586 9818 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].D1
rlabel metal2 3586 7380 3586 7380 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].D1_BUF
rlabel metal2 5141 9804 5141 9804 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].D2
rlabel metal2 5141 8658 5141 8658 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].D2_BUF
rlabel metal2 7139 9678 7139 9678 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT
flabel metal1 5562 9172 5582 9210 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX
flabel metal1 5534 8718 5562 8756 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_BUF
flabel metal3 7052 9506 7082 9646 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal3 7052 8816 7082 8956 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 8816 5102 8956 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 9506 5102 9646 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal2 5142 9722 5142 9722 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D2
flabel metal2 5222 9726 5222 9726 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D3
flabel metal2 5304 9726 5304 9726 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D4
flabel metal2 5384 9728 5384 9728 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D5
flabel metal2 5462 9728 5462 9728 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D6
flabel metal2 5542 9726 5542 9726 1 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D7
flabel metal1 6516 9670 6556 9694 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal2 6518 8748 6556 8772 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal1 5872 9146 5872 9146 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_
flabel metal1 6908 8742 6936 8766 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VREFH
flabel metal1 6986 9666 7016 9686 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VREFL
rlabel metal3 148 8359 148 8359 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VCC
rlabel metal3 166 7654 166 7654 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VSS
rlabel metal2 295 8554 295 8554 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0
rlabel metal2 406 8554 406 8554 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VREFL
rlabel metal2 301 7404 301 7404 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 7387 409 7387 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VREFH
rlabel metal2 5056 8445 5056 8445 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT
rlabel metal2 3586 7386 3586 7386 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 8572 3584 8572 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1
flabel metal1 3492 8334 3492 8334 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 7620 3478 7620 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 8030 1254 8030 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 8298 2662 8298 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 8124 1266 8124 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 7946 624 7946 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 7832 614 7832 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 8270 634 8270 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 7588 528 7728 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 8278 528 8418 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 7943 3624 7982 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 7489 3603 7528 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 8278 5124 8418 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 7588 5124 7728 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 8442 4597 8467 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 7519 4598 7543 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 7918 3914 7918 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 7588 3462 7728 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 8278 3462 8418 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 8475 4888 8475 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 7509 5041 7509 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 9587 148 9587 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VCC
rlabel metal3 166 8882 166 8882 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VSS
rlabel metal2 295 9782 295 9782 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D0
rlabel metal2 406 9782 406 9782 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFL
rlabel metal2 301 8632 301 8632 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 8615 409 8615 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH
rlabel metal2 5056 9673 5056 9673 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT
rlabel metal2 3586 8614 3586 8614 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 9800 3584 9800 7 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D1
flabel metal1 3492 9562 3492 9562 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 8848 3478 8848 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 9258 1254 9258 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 9526 2662 9526 3 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 9352 1266 9352 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 9174 624 9174 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 9060 614 9060 7 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 9498 634 9498 5 FreeSans 400 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 8816 528 8956 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 9506 528 9646 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 9171 3624 9210 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 8717 3603 8756 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 9506 5124 9646 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 8816 5124 8956 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 9670 4597 9695 3 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 8747 4598 8771 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 9146 3914 9146 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 8816 3462 8956 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 9506 3462 9646 7 FreeSans 600 0 0 0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 9703 4888 9703 1 FreeSans 480 0 0 40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 8737 5041 8737 5 FreeSans 480 0 0 -40 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal2 72 14648 72 14648 7 5_bit_dac_0[1].VCC
rlabel metal2 170 14654 170 14654 7 5_bit_dac_0[1].VSS
rlabel metal2 308 19604 308 19604 7 5_bit_dac_0[1].D0
rlabel metal2 416 19592 416 19592 7 5_bit_dac_0[1].VREFL
rlabel metal2 312 9868 312 9868 7 5_bit_dac_0[1].D0_BUF
rlabel metal2 402 9858 402 9858 7 5_bit_dac_0[1].VREFH
rlabel metal2 3574 9846 3574 9846 7 5_bit_dac_0[1].D1_BUF
rlabel metal2 3586 19614 3586 19614 7 5_bit_dac_0[1].D1
rlabel metal2 5150 19624 5150 19624 7 5_bit_dac_0[1].D2
rlabel metal2 5222 19622 5222 19622 7 5_bit_dac_0[1].D3
rlabel metal2 5302 19630 5302 19630 7 5_bit_dac_0[1].D4
rlabel metal2 5152 11120 5152 11120 3 5_bit_dac_0[1].D2_BUF
rlabel metal2 5220 11130 5220 11130 3 5_bit_dac_0[1].D3_BUF
rlabel metal2 5294 11108 5294 11108 3 5_bit_dac_0[1].D4_BUF
rlabel metal2 7176 14908 7176 14908 3 5_bit_dac_0[1].VOUT
flabel metal1 5562 15312 5582 15350 7 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.DX
flabel metal1 5534 14858 5562 14896 7 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.DX_BUF
flabel metal3 7052 15646 7082 15786 3 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VCC
flabel metal3 7052 14956 7082 15096 3 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VSS
flabel metal3 5072 14956 5102 15096 7 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VSS
flabel metal3 5072 15646 5102 15786 7 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VCC
flabel metal2 5142 15862 5142 15862 1 FreeSans 400 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.D2
flabel metal2 5222 15866 5222 15866 1 FreeSans 400 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.D3
flabel metal2 5304 15866 5304 15866 1 FreeSans 400 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.D4
flabel metal2 5384 15868 5384 15868 1 FreeSans 400 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.D5
flabel metal2 5462 15868 5462 15868 1 FreeSans 400 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.D6
flabel metal2 5542 15866 5542 15866 1 FreeSans 400 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.D7
flabel metal1 6516 15810 6556 15834 3 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VOUT
flabel metal2 6518 14888 6556 14912 7 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VOUT
flabel metal1 5872 15286 5872 15286 7 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.DX_
flabel metal1 6908 14882 6936 14906 3 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VREFH
flabel metal1 6986 15806 7016 15826 3 FreeSans 600 0 0 0 5_bit_dac_0[1].switch_n_3v3_0.VREFL
rlabel metal2 74 14296 74 14296 7 5_bit_dac_0[1].4_bit_dac_0[0].VCC
rlabel metal2 182 13578 182 13578 7 5_bit_dac_0[1].4_bit_dac_0[0].VSS
rlabel metal2 312 14702 312 14702 7 5_bit_dac_0[1].4_bit_dac_0[0].D0
rlabel metal2 420 14702 420 14702 7 5_bit_dac_0[1].4_bit_dac_0[0].VREFL
rlabel metal2 316 9846 316 9846 7 5_bit_dac_0[1].4_bit_dac_0[0].D0_BUF
rlabel metal2 416 9840 416 9840 3 5_bit_dac_0[1].4_bit_dac_0[0].VREFH
rlabel metal2 3592 14722 3592 14722 3 5_bit_dac_0[1].4_bit_dac_0[0].D1
rlabel metal2 3574 9832 3574 9832 3 5_bit_dac_0[1].4_bit_dac_0[0].D1_BUF
rlabel metal2 5150 14724 5150 14724 3 5_bit_dac_0[1].4_bit_dac_0[0].D2
rlabel metal2 5222 14722 5222 14722 3 5_bit_dac_0[1].4_bit_dac_0[0].D3
rlabel metal2 5140 11106 5140 11106 3 5_bit_dac_0[1].4_bit_dac_0[0].D2_BUF
rlabel metal2 5212 11114 5212 11114 3 5_bit_dac_0[1].4_bit_dac_0[0].D3_BUF
rlabel metal2 7142 13358 7142 13358 3 5_bit_dac_0[1].4_bit_dac_0[0].VOUT
flabel metal1 5562 12856 5582 12894 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX
flabel metal1 5534 12402 5562 12440 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_BUF
flabel metal3 7052 13190 7082 13330 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VCC
flabel metal3 7052 12500 7082 12640 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VSS
flabel metal3 5072 12500 5102 12640 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VSS
flabel metal3 5072 13190 5102 13330 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VCC
flabel metal2 5142 13406 5142 13406 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2
flabel metal2 5222 13410 5222 13410 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D3
flabel metal2 5304 13410 5304 13410 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D4
flabel metal2 5384 13412 5384 13412 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D5
flabel metal2 5462 13412 5462 13412 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D6
flabel metal2 5542 13410 5542 13410 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D7
flabel metal1 6516 13354 6556 13378 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VOUT
flabel metal2 6518 12432 6556 12456 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VOUT
flabel metal1 5872 12830 5872 12830 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_
flabel metal1 6908 12426 6936 12450 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VREFH
flabel metal1 6986 13350 7016 13370 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.VREFL
rlabel metal3 18 12058 18 12058 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VCC
rlabel metal3 26 11346 26 11346 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VSS
rlabel metal2 302 12254 302 12254 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0
rlabel metal2 406 12256 406 12256 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VREFL
rlabel metal2 304 9844 304 9844 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0_BUF
rlabel metal2 400 9836 400 9836 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VREFH
rlabel metal2 3586 12274 3586 12274 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1
rlabel metal2 3586 9836 3586 9836 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1_BUF
rlabel metal2 5141 12260 5141 12260 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D2
rlabel metal2 5141 11114 5141 11114 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D2_BUF
rlabel metal2 7139 12134 7139 12134 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT
flabel metal1 5562 11628 5582 11666 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX
flabel metal1 5534 11174 5562 11212 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_BUF
flabel metal3 7052 11962 7082 12102 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal3 7052 11272 7082 11412 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 11272 5102 11412 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 11962 5102 12102 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal2 5142 12178 5142 12178 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D2
flabel metal2 5222 12182 5222 12182 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D3
flabel metal2 5304 12182 5304 12182 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D4
flabel metal2 5384 12184 5384 12184 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D5
flabel metal2 5462 12184 5462 12184 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D6
flabel metal2 5542 12182 5542 12182 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.D7
flabel metal1 6516 12126 6556 12150 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal2 6518 11204 6556 11228 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal1 5872 11602 5872 11602 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_
flabel metal1 6908 11198 6936 11222 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VREFH
flabel metal1 6986 12122 7016 12142 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.VREFL
rlabel metal3 148 10815 148 10815 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VCC
rlabel metal3 166 10110 166 10110 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VSS
rlabel metal2 295 11010 295 11010 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0
rlabel metal2 406 11010 406 11010 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VREFL
rlabel metal2 301 9860 301 9860 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 9843 409 9843 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VREFH
rlabel metal2 5056 10901 5056 10901 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT
rlabel metal2 3586 9842 3586 9842 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 11028 3584 11028 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1
flabel metal1 3492 10790 3492 10790 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 10076 3478 10076 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 10486 1254 10486 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 10754 2662 10754 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 10580 1266 10580 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 10402 624 10402 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 10288 614 10288 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 10726 634 10726 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 10044 528 10184 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 10734 528 10874 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 10399 3624 10438 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 9945 3603 9984 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 10734 5124 10874 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 10044 5124 10184 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 10898 4597 10923 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 9975 4598 9999 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 10374 3914 10374 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 10044 3462 10184 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 10734 3462 10874 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 10931 4888 10931 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 9965 5041 9965 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 12043 148 12043 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VCC
rlabel metal3 166 11338 166 11338 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VSS
rlabel metal2 295 12238 295 12238 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D0
rlabel metal2 406 12238 406 12238 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFL
rlabel metal2 301 11088 301 11088 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 11071 409 11071 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH
rlabel metal2 5056 12129 5056 12129 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT
rlabel metal2 3586 11070 3586 11070 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 12256 3584 12256 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].D1
flabel metal1 3492 12018 3492 12018 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 11304 3478 11304 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 11714 1254 11714 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 11982 2662 11982 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 11808 1266 11808 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 11630 624 11630 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 11516 614 11516 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 11954 634 11954 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 11272 528 11412 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 11962 528 12102 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 11627 3624 11666 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 11173 3603 11212 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 11962 5124 12102 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 11272 5124 11412 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 12126 4597 12151 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 11203 4598 11227 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 11602 3914 11602 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 11272 3462 11412 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 11962 3462 12102 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 12159 4888 12159 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 11193 5041 11193 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal3 18 14514 18 14514 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VCC
rlabel metal3 26 13802 26 13802 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VSS
rlabel metal2 302 14710 302 14710 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].D0
rlabel metal2 406 14712 406 14712 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFL
rlabel metal2 304 12300 304 12300 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].D0_BUF
rlabel metal2 400 12292 400 12292 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH
rlabel metal2 3586 14730 3586 14730 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].D1
rlabel metal2 3586 12292 3586 12292 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].D1_BUF
rlabel metal2 5141 14716 5141 14716 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].D2
rlabel metal2 5141 13570 5141 13570 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].D2_BUF
rlabel metal2 7139 14590 7139 14590 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT
flabel metal1 5562 14084 5582 14122 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX
flabel metal1 5534 13630 5562 13668 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_BUF
flabel metal3 7052 14418 7082 14558 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal3 7052 13728 7082 13868 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 13728 5102 13868 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 14418 5102 14558 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal2 5142 14634 5142 14634 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D2
flabel metal2 5222 14638 5222 14638 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D3
flabel metal2 5304 14638 5304 14638 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D4
flabel metal2 5384 14640 5384 14640 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D5
flabel metal2 5462 14640 5462 14640 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D6
flabel metal2 5542 14638 5542 14638 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.D7
flabel metal1 6516 14582 6556 14606 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal2 6518 13660 6556 13684 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal1 5872 14058 5872 14058 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_
flabel metal1 6908 13654 6936 13678 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VREFH
flabel metal1 6986 14578 7016 14598 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.VREFL
rlabel metal3 148 13271 148 13271 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VCC
rlabel metal3 166 12566 166 12566 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VSS
rlabel metal2 295 13466 295 13466 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0
rlabel metal2 406 13466 406 13466 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VREFL
rlabel metal2 301 12316 301 12316 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 12299 409 12299 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VREFH
rlabel metal2 5056 13357 5056 13357 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT
rlabel metal2 3586 12298 3586 12298 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 13484 3584 13484 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1
flabel metal1 3492 13246 3492 13246 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 12532 3478 12532 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 12942 1254 12942 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 13210 2662 13210 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 13036 1266 13036 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 12858 624 12858 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 12744 614 12744 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 13182 634 13182 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 12500 528 12640 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 13190 528 13330 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 12855 3624 12894 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 12401 3603 12440 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 13190 5124 13330 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 12500 5124 12640 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 13354 4597 13379 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 12431 4598 12455 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 12830 3914 12830 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 12500 3462 12640 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 13190 3462 13330 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 13387 4888 13387 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 12421 5041 12421 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 14499 148 14499 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VCC
rlabel metal3 166 13794 166 13794 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VSS
rlabel metal2 295 14694 295 14694 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D0
rlabel metal2 406 14694 406 14694 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFL
rlabel metal2 301 13544 301 13544 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 13527 409 13527 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH
rlabel metal2 5056 14585 5056 14585 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT
rlabel metal2 3586 13526 3586 13526 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 14712 3584 14712 7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].D1
flabel metal1 3492 14474 3492 14474 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 13760 3478 13760 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 14170 1254 14170 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 14438 2662 14438 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 14264 1266 14264 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 14086 624 14086 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 13972 614 13972 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 14410 634 14410 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 13728 528 13868 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 14418 528 14558 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 14083 3624 14122 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 13629 3603 13668 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 14418 5124 14558 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 13728 5124 13868 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 14582 4597 14607 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 13659 4598 13683 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 14058 3914 14058 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 13728 3462 13868 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 14418 3462 14558 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 14615 4888 14615 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 13649 5041 13649 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal2 74 19208 74 19208 7 5_bit_dac_0[1].4_bit_dac_0[1].VCC
rlabel metal2 182 18490 182 18490 7 5_bit_dac_0[1].4_bit_dac_0[1].VSS
rlabel metal2 312 19614 312 19614 7 5_bit_dac_0[1].4_bit_dac_0[1].D0
rlabel metal2 420 19614 420 19614 7 5_bit_dac_0[1].4_bit_dac_0[1].VREFL
rlabel metal2 316 14758 316 14758 7 5_bit_dac_0[1].4_bit_dac_0[1].D0_BUF
rlabel metal2 416 14752 416 14752 3 5_bit_dac_0[1].4_bit_dac_0[1].VREFH
rlabel metal2 3592 19634 3592 19634 3 5_bit_dac_0[1].4_bit_dac_0[1].D1
rlabel metal2 3574 14744 3574 14744 3 5_bit_dac_0[1].4_bit_dac_0[1].D1_BUF
rlabel metal2 5150 19636 5150 19636 3 5_bit_dac_0[1].4_bit_dac_0[1].D2
rlabel metal2 5222 19634 5222 19634 3 5_bit_dac_0[1].4_bit_dac_0[1].D3
rlabel metal2 5140 16018 5140 16018 3 5_bit_dac_0[1].4_bit_dac_0[1].D2_BUF
rlabel metal2 5212 16026 5212 16026 3 5_bit_dac_0[1].4_bit_dac_0[1].D3_BUF
rlabel metal2 7142 18270 7142 18270 3 5_bit_dac_0[1].4_bit_dac_0[1].VOUT
flabel metal1 5562 17768 5582 17806 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX
flabel metal1 5534 17314 5562 17352 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_BUF
flabel metal3 7052 18102 7082 18242 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VCC
flabel metal3 7052 17412 7082 17552 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VSS
flabel metal3 5072 17412 5102 17552 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VSS
flabel metal3 5072 18102 5102 18242 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VCC
flabel metal2 5142 18318 5142 18318 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2
flabel metal2 5222 18322 5222 18322 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D3
flabel metal2 5304 18322 5304 18322 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D4
flabel metal2 5384 18324 5384 18324 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D5
flabel metal2 5462 18324 5462 18324 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D6
flabel metal2 5542 18322 5542 18322 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D7
flabel metal1 6516 18266 6556 18290 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VOUT
flabel metal2 6518 17344 6556 17368 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VOUT
flabel metal1 5872 17742 5872 17742 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_
flabel metal1 6908 17338 6936 17362 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VREFH
flabel metal1 6986 18262 7016 18282 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.VREFL
rlabel metal3 18 16970 18 16970 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VCC
rlabel metal3 26 16258 26 16258 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VSS
rlabel metal2 302 17166 302 17166 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0
rlabel metal2 406 17168 406 17168 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VREFL
rlabel metal2 304 14756 304 14756 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0_BUF
rlabel metal2 400 14748 400 14748 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VREFH
rlabel metal2 3586 17186 3586 17186 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1
rlabel metal2 3586 14748 3586 14748 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1_BUF
rlabel metal2 5141 17172 5141 17172 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D2
rlabel metal2 5141 16026 5141 16026 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D2_BUF
rlabel metal2 7139 17046 7139 17046 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT
flabel metal1 5562 16540 5582 16578 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX
flabel metal1 5534 16086 5562 16124 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_BUF
flabel metal3 7052 16874 7082 17014 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal3 7052 16184 7082 16324 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 16184 5102 16324 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VSS
flabel metal3 5072 16874 5102 17014 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VCC
flabel metal2 5142 17090 5142 17090 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D2
flabel metal2 5222 17094 5222 17094 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D3
flabel metal2 5304 17094 5304 17094 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D4
flabel metal2 5384 17096 5384 17096 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D5
flabel metal2 5462 17096 5462 17096 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D6
flabel metal2 5542 17094 5542 17094 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.D7
flabel metal1 6516 17038 6556 17062 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal2 6518 16116 6556 16140 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VOUT
flabel metal1 5872 16514 5872 16514 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_
flabel metal1 6908 16110 6936 16134 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VREFH
flabel metal1 6986 17034 7016 17054 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.VREFL
rlabel metal3 148 15727 148 15727 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VCC
rlabel metal3 166 15022 166 15022 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VSS
rlabel metal2 295 15922 295 15922 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0
rlabel metal2 406 15922 406 15922 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VREFL
rlabel metal2 301 14772 301 14772 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 14755 409 14755 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VREFH
rlabel metal2 5056 15813 5056 15813 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT
rlabel metal2 3586 14754 3586 14754 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 15940 3584 15940 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1
flabel metal1 3492 15702 3492 15702 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 14988 3478 14988 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 15398 1254 15398 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 15666 2662 15666 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 15492 1266 15492 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 15314 624 15314 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 15200 614 15200 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 15638 634 15638 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 14956 528 15096 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 15646 528 15786 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 15311 3624 15350 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 14857 3603 14896 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 15646 5124 15786 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 14956 5124 15096 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 15810 4597 15835 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 14887 4598 14911 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 15286 3914 15286 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 14956 3462 15096 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 15646 3462 15786 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 15843 4888 15843 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 14877 5041 14877 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 16955 148 16955 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VCC
rlabel metal3 166 16250 166 16250 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VSS
rlabel metal2 295 17150 295 17150 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D0
rlabel metal2 406 17150 406 17150 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFL
rlabel metal2 301 16000 301 16000 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 15983 409 15983 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH
rlabel metal2 5056 17041 5056 17041 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT
rlabel metal2 3586 15982 3586 15982 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 17168 3584 17168 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].D1
flabel metal1 3492 16930 3492 16930 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 16216 3478 16216 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 16626 1254 16626 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 16894 2662 16894 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 16720 1266 16720 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 16542 624 16542 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 16428 614 16428 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 16866 634 16866 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 16184 528 16324 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 16874 528 17014 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 16539 3624 16578 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 16085 3603 16124 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 16874 5124 17014 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 16184 5124 16324 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 17038 4597 17063 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 16115 4598 16139 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 16514 3914 16514 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 16184 3462 16324 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 16874 3462 17014 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 17071 4888 17071 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 16105 5041 16105 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
rlabel metal3 18 19426 18 19426 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VCC
rlabel metal3 26 18714 26 18714 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VSS
rlabel metal2 302 19622 302 19622 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].D0
rlabel metal2 406 19624 406 19624 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFL
rlabel metal2 304 17212 304 17212 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].D0_BUF
rlabel metal2 400 17204 400 17204 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH
rlabel metal2 3586 19642 3586 19642 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].D1
rlabel metal2 3586 17204 3586 17204 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].D1_BUF
rlabel metal2 5141 19628 5141 19628 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].D2
rlabel metal2 5141 18482 5141 18482 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].D2_BUF
rlabel metal2 7139 19502 7139 19502 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT
flabel metal1 5562 18996 5582 19034 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX
flabel metal1 5534 18542 5562 18580 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_BUF
flabel metal3 7052 19330 7082 19470 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal3 7052 18640 7082 18780 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 18640 5102 18780 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VSS
flabel metal3 5072 19330 5102 19470 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VCC
flabel metal2 5142 19546 5142 19546 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D2
flabel metal2 5222 19550 5222 19550 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D3
flabel metal2 5304 19550 5304 19550 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D4
flabel metal2 5384 19552 5384 19552 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D5
flabel metal2 5462 19552 5462 19552 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D6
flabel metal2 5542 19550 5542 19550 1 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.D7
flabel metal1 6516 19494 6556 19518 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal2 6518 18572 6556 18596 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VOUT
flabel metal1 5872 18970 5872 18970 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_
flabel metal1 6908 18566 6936 18590 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VREFH
flabel metal1 6986 19490 7016 19510 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.VREFL
rlabel metal3 148 18183 148 18183 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VCC
rlabel metal3 166 17478 166 17478 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VSS
rlabel metal2 295 18378 295 18378 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0
rlabel metal2 406 18378 406 18378 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VREFL
rlabel metal2 301 17228 301 17228 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0_BUF
rlabel metal2 409 17211 409 17211 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VREFH
rlabel metal2 5056 18269 5056 18269 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT
rlabel metal2 3586 17210 3586 17210 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1_BUF
rlabel metal2 3584 18396 3584 18396 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1
flabel metal1 3492 18158 3492 18158 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3478 17444 3478 17444 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1254 17854 1254 17854 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2662 18122 2662 18122 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1266 17948 1266 17948 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 624 17770 624 17770 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 614 17656 614 17656 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 634 18094 634 18094 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 498 17412 528 17552 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 498 18102 528 18242 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3604 17767 3624 17806 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3575 17313 3603 17352 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 18102 5124 18242 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 5094 17412 5124 17552 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4558 18266 4597 18291 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 17343 4598 17367 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 17742 3914 17742 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3432 17412 3462 17552 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3432 18102 3462 18242 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4888 18299 4888 18299 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 17333 5041 17333 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 148 19411 148 19411 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VCC
rlabel metal3 166 18706 166 18706 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VSS
rlabel metal2 295 19606 295 19606 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D0
rlabel metal2 406 19606 406 19606 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFL
rlabel metal2 301 18456 301 18456 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D0_BUF
rlabel metal2 409 18439 409 18439 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH
rlabel metal2 5056 19497 5056 19497 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT
rlabel metal2 3586 18438 3586 18438 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D1_BUF
rlabel metal2 3584 19624 3584 19624 7 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].D1
flabel metal1 3492 19386 3492 19386 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3478 18672 3478 18672 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1254 19082 1254 19082 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2662 19350 2662 19350 3 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1266 19176 1266 19176 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 624 18998 624 18998 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 614 18884 614 18884 7 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 634 19322 634 19322 5 FreeSans 400 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 498 18640 528 18780 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 498 19330 528 19470 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3604 18995 3624 19034 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3575 18541 3603 18580 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 5094 19330 5124 19470 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 5094 18640 5124 18780 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4558 19494 4597 19519 3 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4559 18571 4598 18595 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3914 18970 3914 18970 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3432 18640 3462 18780 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3432 19330 3462 19470 7 FreeSans 600 0 0 0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4888 19527 4888 19527 1 FreeSans 480 0 0 40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 5041 18561 5041 18561 5 FreeSans 480 0 0 -40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
<< end >>
