* SPICE3 file created from 3_bit_dac.ext - technology: sky130A

.subckt x3_bit_dac VCC VSS D0 VREFL D0_BUF VREFH D1 D1_BUF D2 D2_BUF VOUT
X0 2_bit_dac_0[0]/VOUT D1_BUF 2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 D1_BUF 2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 2_bit_dac_0[0]/VOUT D1_BUF 2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 D1_BUF 2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X9 2_bit_dac_0[0]/switch2n_3v3_0/VREFH D0_BUF 2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X10 2_bit_dac_0[0]/switch2n_3v3_0/VREFH 2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X11 D0_BUF 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X12 2_bit_dac_0[1]/VREFH D0_BUF 2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X13 2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X14 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X15 2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X16 2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X17 2_bit_dac_0[0]/switch2n_3v3_0/R_H D0_BUF 2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 2_bit_dac_0[0]/switch2n_3v3_0/R_H 2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X19 2_bit_dac_0[0]/switch2n_3v3_0/R_L 2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X20 2_bit_dac_0[0]/switch2n_3v3_0/R_L D0_BUF 2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X21 D0_BUF 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X22 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X23 2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X24 2_bit_dac_0[1]/VOUT 2_bit_dac_0[0]/D1 2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X25 2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.9 ps=25.8 w=1 l=0.5
X26 2_bit_dac_0[0]/D1 2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X27 2_bit_dac_0[1]/VOUT 2_bit_dac_0[0]/D1 2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X28 2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=1.45 ps=15.8 w=0.5 l=0.5
X29 2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X30 2_bit_dac_0[0]/D1 2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X31 2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X32 2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X33 2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2_bit_dac_0[0]/D0 2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X34 2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X35 2_bit_dac_0[0]/D0 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X36 VREFL 2_bit_dac_0[0]/D0 2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X37 2_bit_dac_0[1]/switch2n_3v3_0/VREFH 2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X38 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X39 2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.361 ps=3.45 w=0.5 l=0.5
X40 2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X41 2_bit_dac_0[1]/switch2n_3v3_0/R_H 2_bit_dac_0[0]/D0 2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X42 2_bit_dac_0[1]/switch2n_3v3_0/R_H 2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X43 2_bit_dac_0[1]/switch2n_3v3_0/R_L VREFL VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X44 2_bit_dac_0[1]/switch2n_3v3_0/R_L 2_bit_dac_0[0]/D0 2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X45 2_bit_dac_0[0]/D0 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X46 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X47 2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X48 VOUT D2_BUF 2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X49 switch_n_3v3_0/DX_ D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X50 D2_BUF switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X51 VOUT D2_BUF 2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X52 switch_n_3v3_0/DX_ D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X53 2_bit_dac_0[1]/VOUT switch_n_3v3_0/DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X54 D2_BUF switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X55 2_bit_dac_0[0]/VOUT switch_n_3v3_0/DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends



X1 VCC VSS D0 VREFL D0_BUF VREFH D1 D1_BUF D2 D2_BUF VOUT x3_bit_dac

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


V1 VSS 0 dc 0
V2 VCC 0 dc 3.3

V3 VREFH 0 dc 2
V4 VREFL 0 dc 0

V5 D0 0 PULSE(0 1.8 0 1n 1n 1u 2u)
V6 D1 0 PULSE(0 1.8 0 1n 1n 2u 4u)
V7 D2 0 PULSE(0 1.8 0 1n 1n 4u 8u)

.tran 100n 10u
.control
run
plot VOUT
.endc
.end
