magic
tech sky130A
timestamp 1687027365
<< nwell >>
rect 165 916 2345 1140
rect 365 70 2345 916
<< mvnmos >>
rect 540 -457 590 -57
rect 679 -177 729 23
rect 838 -167 888 33
rect 759 -417 809 -217
rect 838 -417 888 -217
rect 979 -387 1079 -187
rect 1108 -387 1208 -187
rect 1299 -382 1399 18
rect 1494 -387 1544 -187
rect 1573 -387 1623 -187
rect 1757 -464 1857 -64
rect 1886 -464 1986 -64
rect 2015 -464 2115 -64
rect 2144 -464 2244 -64
<< mvpmos >>
rect 432 113 532 913
rect 561 113 661 913
rect 882 708 982 908
rect 752 188 852 588
rect 881 188 981 588
rect 1072 113 1172 913
rect 1201 113 1301 913
rect 1412 513 1512 913
rect 1541 513 1641 913
rect 1397 146 1447 346
rect 1602 146 1652 346
rect 1757 112 1857 912
rect 1886 112 1986 912
rect 2015 112 2115 912
rect 2144 112 2244 912
<< mvndiff >>
rect 208 433 250 461
rect 208 416 214 433
rect 244 416 250 433
rect 208 410 250 416
rect 280 433 322 461
rect 280 416 286 433
rect 316 416 322 433
rect 280 410 322 416
rect 204 321 252 327
rect 204 304 210 321
rect 246 304 252 321
rect 204 276 252 304
rect 282 321 330 327
rect 282 304 288 321
rect 324 304 330 321
rect 282 276 330 304
rect 809 27 838 33
rect 650 17 679 23
rect 197 -437 239 -408
rect 197 -454 203 -437
rect 233 -454 239 -437
rect 197 -460 239 -454
rect 413 -437 455 -408
rect 413 -454 419 -437
rect 449 -454 455 -437
rect 413 -460 455 -454
rect 511 -63 540 -57
rect 511 -451 517 -63
rect 534 -451 540 -63
rect 511 -457 540 -451
rect 590 -63 619 -57
rect 590 -451 596 -63
rect 613 -451 619 -63
rect 650 -171 656 17
rect 673 -171 679 17
rect 650 -177 679 -171
rect 729 17 758 23
rect 729 -171 735 17
rect 752 -171 758 17
rect 809 -161 815 27
rect 832 -161 838 27
rect 809 -167 838 -161
rect 888 27 917 33
rect 888 -161 894 27
rect 911 -161 917 27
rect 888 -167 917 -161
rect 1270 12 1299 18
rect 729 -177 758 -171
rect 950 -193 979 -187
rect 730 -223 759 -217
rect 730 -411 736 -223
rect 753 -411 759 -223
rect 730 -417 759 -411
rect 809 -223 838 -217
rect 809 -411 815 -223
rect 832 -411 838 -223
rect 809 -417 838 -411
rect 888 -223 917 -217
rect 888 -411 894 -223
rect 911 -411 917 -223
rect 950 -381 956 -193
rect 973 -381 979 -193
rect 950 -387 979 -381
rect 1079 -193 1108 -187
rect 1079 -381 1085 -193
rect 1102 -381 1108 -193
rect 1079 -387 1108 -381
rect 1208 -193 1237 -187
rect 1208 -381 1214 -193
rect 1231 -381 1237 -193
rect 1208 -387 1237 -381
rect 1270 -376 1276 12
rect 1293 -376 1299 12
rect 1270 -382 1299 -376
rect 1399 12 1428 18
rect 1399 -376 1405 12
rect 1422 -376 1428 12
rect 1728 -70 1757 -64
rect 1399 -382 1428 -376
rect 1465 -193 1494 -187
rect 1465 -381 1471 -193
rect 1488 -381 1494 -193
rect 1465 -387 1494 -381
rect 1544 -193 1573 -187
rect 1544 -381 1550 -193
rect 1567 -381 1573 -193
rect 1544 -387 1573 -381
rect 1623 -193 1652 -187
rect 1623 -381 1629 -193
rect 1646 -381 1652 -193
rect 1623 -387 1652 -381
rect 888 -417 917 -411
rect 590 -457 619 -451
rect 1728 -458 1734 -70
rect 1751 -458 1757 -70
rect 1728 -464 1757 -458
rect 1857 -70 1886 -64
rect 1857 -458 1863 -70
rect 1880 -458 1886 -70
rect 1857 -464 1886 -458
rect 1986 -70 2015 -64
rect 1986 -458 1992 -70
rect 2009 -458 2015 -70
rect 1986 -464 2015 -458
rect 2115 -70 2144 -64
rect 2115 -458 2121 -70
rect 2138 -458 2144 -70
rect 2115 -464 2144 -458
rect 2244 -70 2273 -64
rect 2244 -458 2250 -70
rect 2267 -458 2273 -70
rect 2244 -464 2273 -458
<< mvpdiff >>
rect 403 907 432 913
rect 403 119 409 907
rect 426 119 432 907
rect 403 113 432 119
rect 532 907 561 913
rect 532 119 538 907
rect 555 119 561 907
rect 532 113 561 119
rect 661 907 690 913
rect 661 119 667 907
rect 684 119 690 907
rect 853 902 882 908
rect 853 714 859 902
rect 876 714 882 902
rect 853 708 882 714
rect 982 902 1011 908
rect 982 714 988 902
rect 1005 714 1011 902
rect 982 708 1011 714
rect 1043 907 1072 913
rect 723 582 752 588
rect 723 194 729 582
rect 746 194 752 582
rect 723 188 752 194
rect 852 582 881 588
rect 852 194 858 582
rect 875 194 881 582
rect 852 188 881 194
rect 981 582 1010 588
rect 981 194 987 582
rect 1004 194 1010 582
rect 981 188 1010 194
rect 661 113 690 119
rect 1043 119 1049 907
rect 1066 119 1072 907
rect 1043 113 1072 119
rect 1172 907 1201 913
rect 1172 119 1178 907
rect 1195 119 1201 907
rect 1172 113 1201 119
rect 1301 907 1330 913
rect 1301 119 1307 907
rect 1324 119 1330 907
rect 1383 907 1412 913
rect 1383 519 1389 907
rect 1406 519 1412 907
rect 1383 513 1412 519
rect 1512 907 1541 913
rect 1512 519 1518 907
rect 1535 519 1541 907
rect 1512 513 1541 519
rect 1641 907 1670 913
rect 1641 519 1647 907
rect 1664 519 1670 907
rect 1641 513 1670 519
rect 1728 906 1757 912
rect 1368 340 1397 346
rect 1368 152 1374 340
rect 1391 152 1397 340
rect 1368 146 1397 152
rect 1447 340 1476 346
rect 1447 152 1453 340
rect 1470 152 1476 340
rect 1447 146 1476 152
rect 1573 340 1602 346
rect 1573 152 1579 340
rect 1596 152 1602 340
rect 1573 146 1602 152
rect 1652 340 1681 346
rect 1652 152 1658 340
rect 1675 152 1681 340
rect 1652 146 1681 152
rect 1301 113 1330 119
rect 1728 118 1734 906
rect 1751 118 1757 906
rect 1728 112 1757 118
rect 1857 906 1886 912
rect 1857 118 1863 906
rect 1880 118 1886 906
rect 1857 112 1886 118
rect 1986 906 2015 912
rect 1986 118 1992 906
rect 2009 118 2015 906
rect 1986 112 2015 118
rect 2115 906 2144 912
rect 2115 118 2121 906
rect 2138 118 2144 906
rect 2115 112 2144 118
rect 2244 906 2273 912
rect 2244 118 2250 906
rect 2267 118 2273 906
rect 2244 112 2273 118
<< mvndiffc >>
rect 214 416 244 433
rect 286 416 316 433
rect 210 304 246 321
rect 288 304 324 321
rect 203 -454 233 -437
rect 419 -454 449 -437
rect 517 -451 534 -63
rect 596 -451 613 -63
rect 656 -171 673 17
rect 735 -171 752 17
rect 815 -161 832 27
rect 894 -161 911 27
rect 736 -411 753 -223
rect 815 -411 832 -223
rect 894 -411 911 -223
rect 956 -381 973 -193
rect 1085 -381 1102 -193
rect 1214 -381 1231 -193
rect 1276 -376 1293 12
rect 1405 -376 1422 12
rect 1471 -381 1488 -193
rect 1550 -381 1567 -193
rect 1629 -381 1646 -193
rect 1734 -458 1751 -70
rect 1863 -458 1880 -70
rect 1992 -458 2009 -70
rect 2121 -458 2138 -70
rect 2250 -458 2267 -70
<< mvpdiffc >>
rect 409 119 426 907
rect 538 119 555 907
rect 667 119 684 907
rect 859 714 876 902
rect 988 714 1005 902
rect 729 194 746 582
rect 858 194 875 582
rect 987 194 1004 582
rect 1049 119 1066 907
rect 1178 119 1195 907
rect 1307 119 1324 907
rect 1389 519 1406 907
rect 1518 519 1535 907
rect 1647 519 1664 907
rect 1374 152 1391 340
rect 1453 152 1470 340
rect 1579 152 1596 340
rect 1658 152 1675 340
rect 1734 118 1751 906
rect 1863 118 1880 906
rect 1992 118 2009 906
rect 2121 118 2138 906
rect 2250 118 2267 906
<< mvpsubdiff >>
rect 535 -530 2100 -505
rect 535 -630 595 -530
rect 2055 -630 2100 -530
rect 535 -655 2100 -630
<< mvnsubdiff >>
rect 255 1070 2020 1100
rect 255 980 305 1070
rect 815 980 875 1070
rect 1380 980 1460 1070
rect 1970 980 2020 1070
rect 255 950 2020 980
<< mvpsubdiffcont >>
rect 595 -630 2055 -530
<< mvnsubdiffcont >>
rect 305 980 815 1070
rect 875 980 1380 1070
rect 1460 980 1970 1070
<< poly >>
rect 432 913 532 926
rect 561 913 661 926
rect 882 908 982 921
rect 1072 913 1172 926
rect 1201 913 1301 926
rect 1412 913 1512 926
rect 1541 913 1641 926
rect 882 695 982 708
rect 920 669 948 695
rect 917 664 951 669
rect 917 646 925 664
rect 943 646 951 664
rect 917 641 951 646
rect 752 588 852 601
rect 881 588 981 601
rect 752 175 852 188
rect 881 175 981 188
rect 796 149 824 175
rect 921 149 949 175
rect 793 144 827 149
rect 793 121 801 144
rect 819 121 827 144
rect 793 116 827 121
rect 918 144 952 149
rect 918 121 926 144
rect 944 121 952 144
rect 918 116 952 121
rect 1757 912 1857 925
rect 1886 912 1986 925
rect 2015 912 2115 925
rect 2144 912 2244 925
rect 1412 500 1512 513
rect 1541 500 1641 513
rect 1451 474 1479 500
rect 1581 474 1609 500
rect 1448 469 1482 474
rect 1448 451 1456 469
rect 1474 451 1482 469
rect 1448 446 1482 451
rect 1578 469 1612 474
rect 1578 451 1586 469
rect 1604 451 1612 469
rect 1578 446 1612 451
rect 1397 346 1447 359
rect 1602 346 1652 359
rect 1397 133 1447 146
rect 1602 133 1652 146
rect 432 100 532 113
rect 561 100 661 113
rect 1072 100 1172 113
rect 1201 100 1301 113
rect 1406 109 1434 133
rect 1606 109 1634 133
rect 1403 104 1437 109
rect 476 74 504 100
rect 606 74 634 100
rect 848 89 881 94
rect 675 79 708 84
rect 473 69 507 74
rect 473 51 481 69
rect 499 51 507 69
rect 473 46 507 51
rect 603 69 637 74
rect 603 51 611 69
rect 629 51 637 69
rect 675 62 683 79
rect 700 62 708 79
rect 848 72 856 89
rect 873 72 881 89
rect 1111 74 1139 100
rect 1241 74 1269 100
rect 1403 81 1411 104
rect 1429 81 1437 104
rect 1403 76 1437 81
rect 1603 104 1637 109
rect 1603 81 1611 104
rect 1629 81 1637 104
rect 1757 99 1857 112
rect 1886 99 1986 112
rect 2015 99 2115 112
rect 2144 99 2244 112
rect 1603 76 1637 81
rect 1791 74 1819 99
rect 1921 74 1949 99
rect 2051 74 2079 99
rect 2176 74 2204 99
rect 848 67 881 72
rect 1108 69 1142 74
rect 675 57 708 62
rect 603 46 637 51
rect 683 36 699 57
rect 856 46 872 67
rect 1108 51 1116 69
rect 1134 51 1142 69
rect 1108 46 1142 51
rect 1238 69 1272 74
rect 1238 51 1246 69
rect 1264 51 1272 69
rect 1238 46 1272 51
rect 1788 69 1822 74
rect 1788 46 1796 69
rect 1814 46 1822 69
rect 679 23 729 36
rect 838 33 888 46
rect 1788 41 1822 46
rect 1918 69 1952 74
rect 1918 46 1926 69
rect 1944 46 1952 69
rect 1918 41 1952 46
rect 2048 69 2082 74
rect 2048 46 2056 69
rect 2074 46 2082 69
rect 2048 41 2082 46
rect 2173 69 2207 74
rect 2173 46 2181 69
rect 2199 46 2207 69
rect 2173 41 2207 46
rect 557 -1 590 4
rect 557 -18 565 -1
rect 582 -18 590 -1
rect 557 -23 590 -18
rect 566 -44 582 -23
rect 540 -57 590 -44
rect 1299 18 1399 31
rect 679 -190 729 -177
rect 838 -180 888 -167
rect 979 -187 1079 -174
rect 1108 -187 1208 -174
rect 759 -217 809 -204
rect 838 -217 888 -204
rect 1788 -8 1821 -3
rect 1788 -25 1796 -8
rect 1813 -25 1821 -8
rect 1788 -30 1821 -25
rect 1921 -8 1954 -3
rect 1921 -25 1929 -8
rect 1946 -25 1954 -8
rect 1921 -30 1954 -25
rect 2048 -8 2081 -3
rect 2048 -25 2056 -8
rect 2073 -25 2081 -8
rect 2048 -30 2081 -25
rect 2179 -8 2212 -3
rect 2179 -25 2187 -8
rect 2204 -25 2212 -8
rect 2179 -30 2212 -25
rect 1796 -51 1812 -30
rect 1930 -51 1946 -30
rect 2056 -51 2072 -30
rect 2188 -51 2204 -30
rect 1757 -64 1857 -51
rect 1886 -64 1986 -51
rect 2015 -64 2115 -51
rect 2144 -64 2244 -51
rect 1507 -121 1542 -116
rect 1507 -144 1515 -121
rect 1534 -144 1542 -121
rect 1507 -149 1542 -144
rect 1572 -121 1607 -116
rect 1572 -144 1580 -121
rect 1599 -144 1607 -121
rect 1572 -149 1607 -144
rect 1510 -174 1539 -149
rect 1575 -174 1604 -149
rect 1494 -187 1544 -174
rect 1573 -187 1623 -174
rect 979 -400 1079 -387
rect 1108 -400 1208 -387
rect 1299 -395 1399 -382
rect 759 -430 809 -417
rect 838 -430 888 -417
rect 1011 -421 1039 -400
rect 1008 -426 1042 -421
rect 1153 -422 1181 -400
rect 1336 -420 1364 -395
rect 1494 -400 1544 -387
rect 1573 -400 1623 -387
rect 761 -451 789 -430
rect 856 -451 884 -430
rect 1008 -449 1016 -426
rect 1034 -449 1042 -426
rect 758 -456 792 -451
rect 540 -470 590 -457
rect 758 -480 766 -456
rect 784 -480 792 -456
rect 758 -485 792 -480
rect 853 -456 887 -451
rect 1008 -454 1042 -449
rect 1150 -427 1184 -422
rect 1150 -450 1158 -427
rect 1176 -450 1184 -427
rect 1150 -455 1184 -450
rect 1333 -425 1367 -420
rect 1333 -449 1341 -425
rect 1359 -449 1367 -425
rect 1333 -454 1367 -449
rect 853 -480 861 -456
rect 879 -480 887 -456
rect 1757 -477 1857 -464
rect 1886 -477 1986 -464
rect 2015 -477 2115 -464
rect 2144 -477 2244 -464
rect 853 -485 887 -480
<< polycont >>
rect 925 646 943 664
rect 801 121 819 144
rect 926 121 944 144
rect 1456 451 1474 469
rect 1586 451 1604 469
rect 481 51 499 69
rect 611 51 629 69
rect 683 62 700 79
rect 856 72 873 89
rect 1411 81 1429 104
rect 1611 81 1629 104
rect 1116 51 1134 69
rect 1246 51 1264 69
rect 1796 46 1814 69
rect 1926 46 1944 69
rect 2056 46 2074 69
rect 2181 46 2199 69
rect 565 -18 582 -1
rect 1796 -25 1813 -8
rect 1929 -25 1946 -8
rect 2056 -25 2073 -8
rect 2187 -25 2204 -8
rect 1515 -144 1534 -121
rect 1580 -144 1599 -121
rect 1016 -449 1034 -426
rect 766 -480 784 -456
rect 1158 -450 1176 -427
rect 1341 -449 1359 -425
rect 861 -480 879 -456
<< mvndiffres >>
rect 208 841 322 883
rect 208 461 250 841
rect 280 461 322 841
rect 204 92 252 276
rect 282 92 330 276
rect 204 44 330 92
rect 197 -28 311 13
rect 197 -408 239 -28
rect 269 -344 311 -28
rect 341 -28 455 13
rect 341 -344 383 -28
rect 269 -386 383 -344
rect 413 -408 455 -28
<< locali >>
rect 255 1070 2020 1100
rect 255 980 305 1070
rect 815 980 875 1070
rect 1380 980 1460 1070
rect 1970 980 2020 1070
rect 255 950 2020 980
rect 409 907 426 915
rect 283 548 319 551
rect 283 518 286 548
rect 316 518 319 548
rect 212 433 248 487
rect 283 433 319 518
rect 206 416 214 433
rect 244 416 252 433
rect 278 416 286 433
rect 316 416 324 433
rect 212 382 248 416
rect 283 412 319 416
rect 335 382 357 383
rect 212 380 357 382
rect 212 360 335 380
rect 354 360 357 380
rect 212 358 357 360
rect 212 357 355 358
rect 212 321 248 357
rect 294 321 330 331
rect 202 304 210 321
rect 246 304 254 321
rect 280 304 288 321
rect 324 304 332 321
rect 212 298 248 304
rect 294 -410 330 304
rect 409 111 426 119
rect 538 907 555 915
rect 538 111 555 119
rect 667 907 684 915
rect 859 902 876 910
rect 855 714 859 747
rect 988 902 1005 910
rect 876 714 880 747
rect 729 582 746 590
rect 855 582 880 714
rect 988 706 1005 714
rect 1049 907 1066 915
rect 925 669 943 672
rect 925 638 943 641
rect 855 547 858 582
rect 729 186 746 194
rect 875 547 880 582
rect 987 582 1004 590
rect 858 186 875 194
rect 801 149 819 152
rect 926 149 944 152
rect 667 111 684 119
rect 801 113 819 116
rect 926 113 944 116
rect 856 89 873 97
rect 683 85 700 87
rect 481 74 499 77
rect 611 74 629 77
rect 702 72 856 85
rect 987 88 1004 194
rect 1049 111 1066 119
rect 1178 907 1195 915
rect 1178 111 1195 119
rect 1307 907 1324 915
rect 1389 907 1406 915
rect 1389 511 1406 519
rect 1518 907 1535 915
rect 1518 511 1535 519
rect 1647 907 1664 915
rect 1647 511 1664 519
rect 1734 906 1751 914
rect 1456 474 1474 477
rect 1586 474 1604 477
rect 1456 443 1474 446
rect 1586 443 1604 446
rect 1374 340 1391 348
rect 1374 144 1391 152
rect 1453 340 1470 348
rect 1579 340 1596 348
rect 1470 152 1520 170
rect 1453 145 1520 152
rect 1453 144 1470 145
rect 1307 111 1324 119
rect 1411 109 1429 112
rect 873 72 875 85
rect 702 60 875 72
rect 894 71 1004 88
rect 1116 74 1134 77
rect 1246 74 1264 77
rect 683 54 700 60
rect 481 43 499 46
rect 611 43 629 46
rect 815 27 832 35
rect 656 17 673 25
rect 565 -1 582 7
rect 565 -26 582 -18
rect 224 -437 238 -436
rect 195 -454 203 -437
rect 233 -454 241 -437
rect 517 -63 534 -55
rect 415 -437 440 -430
rect 411 -454 419 -437
rect 415 -460 440 -454
rect 517 -459 534 -451
rect 596 -63 613 -55
rect 656 -179 673 -171
rect 735 17 752 25
rect 815 -169 832 -161
rect 894 27 911 71
rect 1052 49 1069 54
rect 953 32 1069 49
rect 1305 73 1340 75
rect 1411 73 1429 76
rect 1305 56 1306 73
rect 1323 56 1340 73
rect 1495 62 1520 145
rect 1579 144 1596 152
rect 1658 340 1675 348
rect 1658 144 1675 152
rect 1611 109 1629 112
rect 1734 110 1751 118
rect 1863 906 1880 914
rect 1863 110 1880 118
rect 1992 906 2009 914
rect 1992 110 2009 118
rect 2121 906 2138 914
rect 2121 110 2138 118
rect 2250 906 2267 914
rect 2250 110 2267 118
rect 1611 73 1629 76
rect 1796 74 1814 77
rect 1926 74 1944 77
rect 2056 74 2074 77
rect 2181 74 2199 77
rect 1305 55 1340 56
rect 1116 43 1134 46
rect 1246 43 1264 46
rect 1276 12 1293 20
rect 1140 5 1161 9
rect 1140 4 1180 5
rect 994 -17 1035 2
rect 1140 -13 1141 4
rect 1158 -13 1180 4
rect 1140 -15 1180 -13
rect 894 -169 911 -161
rect 735 -179 752 -171
rect 956 -193 973 -185
rect 736 -223 753 -215
rect 736 -419 753 -411
rect 815 -223 832 -215
rect 815 -419 832 -411
rect 894 -223 911 -215
rect 956 -389 973 -381
rect 1015 -285 1035 -17
rect 894 -419 911 -411
rect 1015 -421 1035 -305
rect 1085 -193 1102 -185
rect 1085 -389 1102 -381
rect 1160 -355 1180 -15
rect 1160 -419 1180 -375
rect 1214 -193 1231 -185
rect 1214 -389 1231 -381
rect 1320 -40 1340 55
rect 1467 37 1520 62
rect 1683 45 1791 70
rect 1405 12 1422 20
rect 1276 -384 1293 -376
rect 1467 -122 1492 37
rect 1683 -40 1703 45
rect 1819 45 1921 70
rect 1949 45 2051 70
rect 2079 45 2176 70
rect 2204 45 2205 70
rect 1796 38 1814 41
rect 1926 38 1944 41
rect 2056 38 2074 41
rect 2181 38 2199 41
rect 1796 -5 1813 0
rect 1929 -5 1946 0
rect 2056 -5 2073 0
rect 2187 -5 2204 0
rect 1815 -8 2204 -5
rect 1815 -25 1929 -8
rect 1946 -25 2056 -8
rect 2073 -25 2187 -8
rect 1796 -33 1813 -25
rect 1929 -33 1946 -25
rect 2056 -33 2073 -25
rect 2187 -33 2204 -25
rect 1540 -60 1703 -40
rect 1734 -70 1751 -62
rect 1515 -116 1534 -113
rect 1580 -116 1599 -113
rect 1467 -147 1510 -122
rect 1467 -193 1492 -147
rect 1515 -152 1534 -149
rect 1580 -152 1599 -149
rect 1467 -202 1471 -193
rect 1405 -384 1422 -376
rect 1488 -202 1492 -193
rect 1550 -193 1567 -185
rect 1471 -389 1488 -381
rect 1550 -389 1567 -381
rect 1629 -193 1646 -185
rect 1629 -389 1646 -381
rect 1158 -422 1180 -419
rect 1341 -420 1359 -417
rect 766 -451 784 -448
rect 861 -451 879 -448
rect 596 -459 613 -451
rect 789 -481 856 -456
rect 1016 -457 1034 -454
rect 1158 -458 1176 -455
rect 1341 -457 1359 -454
rect 1734 -466 1751 -458
rect 1863 -70 1880 -62
rect 1863 -466 1880 -458
rect 1992 -70 2009 -62
rect 1992 -466 2009 -458
rect 2121 -70 2138 -62
rect 2121 -466 2138 -458
rect 2250 -70 2267 -62
rect 2250 -466 2267 -458
rect 766 -488 784 -485
rect 861 -488 879 -485
rect 535 -530 2100 -505
rect 535 -630 595 -530
rect 2055 -630 2100 -530
rect 535 -655 2100 -630
<< viali >>
rect 305 980 815 1070
rect 875 980 1380 1070
rect 1460 980 1970 1070
rect 286 518 316 548
rect 335 360 354 380
rect 409 119 426 907
rect 538 119 555 907
rect 667 119 684 907
rect 859 714 876 902
rect 729 194 746 582
rect 988 714 1005 902
rect 920 664 948 669
rect 920 646 925 664
rect 925 646 943 664
rect 943 646 948 664
rect 920 641 948 646
rect 858 194 875 582
rect 987 194 1004 582
rect 796 144 824 149
rect 796 121 801 144
rect 801 121 819 144
rect 819 121 824 144
rect 796 116 824 121
rect 921 144 949 149
rect 921 121 926 144
rect 926 121 944 144
rect 944 121 949 144
rect 921 116 949 121
rect 677 79 702 85
rect 476 69 504 74
rect 476 51 481 69
rect 481 51 499 69
rect 499 51 504 69
rect 476 46 504 51
rect 606 69 634 74
rect 606 51 611 69
rect 611 51 629 69
rect 629 51 634 69
rect 677 62 683 79
rect 683 62 700 79
rect 700 62 702 79
rect 856 72 873 89
rect 1049 119 1066 907
rect 1178 119 1195 907
rect 1307 119 1324 907
rect 1389 519 1406 907
rect 1518 519 1535 907
rect 1647 519 1664 907
rect 1451 469 1479 474
rect 1451 451 1456 469
rect 1456 451 1474 469
rect 1474 451 1479 469
rect 1451 446 1479 451
rect 1581 469 1609 474
rect 1581 451 1586 469
rect 1586 451 1604 469
rect 1604 451 1609 469
rect 1581 446 1609 451
rect 1374 152 1391 340
rect 1453 152 1470 340
rect 677 60 702 62
rect 1406 104 1434 109
rect 1406 81 1411 104
rect 1411 81 1429 104
rect 1429 81 1434 104
rect 1406 76 1434 81
rect 606 46 634 51
rect 565 -18 582 -1
rect 207 -437 224 -436
rect 207 -453 224 -437
rect 294 -446 330 -410
rect 440 -437 470 -430
rect 440 -454 449 -437
rect 449 -454 470 -437
rect 440 -460 470 -454
rect 517 -451 534 -63
rect 596 -451 613 -63
rect 656 -171 673 17
rect 735 -171 752 17
rect 815 -161 832 27
rect 1052 54 1069 71
rect 936 32 953 49
rect 1111 69 1139 74
rect 1111 51 1116 69
rect 1116 51 1134 69
rect 1134 51 1139 69
rect 1111 46 1139 51
rect 1241 69 1269 74
rect 1241 51 1246 69
rect 1246 51 1264 69
rect 1264 51 1269 69
rect 1306 56 1323 73
rect 1579 152 1596 340
rect 1658 152 1675 340
rect 1734 118 1751 906
rect 1863 118 1880 906
rect 1992 118 2009 906
rect 2121 118 2138 906
rect 2250 118 2267 906
rect 1606 104 1634 109
rect 1606 81 1611 104
rect 1611 81 1629 104
rect 1629 81 1634 104
rect 1606 76 1634 81
rect 1241 46 1269 51
rect 894 -161 911 27
rect 974 -17 994 2
rect 1141 -13 1158 4
rect 736 -411 753 -223
rect 815 -411 832 -223
rect 894 -411 911 -223
rect 956 -381 973 -193
rect 1015 -305 1035 -285
rect 1085 -381 1102 -193
rect 1160 -375 1180 -355
rect 1214 -381 1231 -193
rect 1276 -376 1293 12
rect 1791 69 1819 74
rect 1791 46 1796 69
rect 1796 46 1814 69
rect 1814 46 1819 69
rect 1320 -60 1340 -40
rect 1405 -376 1422 12
rect 1791 41 1819 46
rect 1921 69 1949 74
rect 1921 46 1926 69
rect 1926 46 1944 69
rect 1944 46 1949 69
rect 1921 41 1949 46
rect 2051 69 2079 74
rect 2051 46 2056 69
rect 2056 46 2074 69
rect 2074 46 2079 69
rect 2051 41 2079 46
rect 2176 69 2204 74
rect 2176 46 2181 69
rect 2181 46 2199 69
rect 2199 46 2204 69
rect 2176 41 2204 46
rect 1795 -8 1815 -5
rect 1795 -25 1796 -8
rect 1796 -25 1813 -8
rect 1813 -25 1815 -8
rect 1929 -25 1946 -8
rect 2056 -25 2073 -8
rect 2187 -25 2204 -8
rect 1523 -60 1540 -40
rect 1510 -121 1539 -116
rect 1510 -144 1515 -121
rect 1515 -144 1534 -121
rect 1534 -144 1539 -121
rect 1510 -149 1539 -144
rect 1575 -121 1604 -116
rect 1575 -144 1580 -121
rect 1580 -144 1599 -121
rect 1599 -144 1604 -121
rect 1575 -149 1604 -144
rect 1471 -381 1488 -193
rect 1550 -381 1567 -193
rect 1629 -381 1646 -193
rect 1011 -426 1039 -421
rect 1011 -449 1016 -426
rect 1016 -449 1034 -426
rect 1034 -449 1039 -426
rect 761 -456 789 -451
rect 856 -456 884 -451
rect 1011 -454 1039 -449
rect 1153 -427 1181 -422
rect 1153 -450 1158 -427
rect 1158 -450 1176 -427
rect 1176 -450 1181 -427
rect 761 -480 766 -456
rect 766 -480 784 -456
rect 784 -480 789 -456
rect 761 -485 789 -480
rect 856 -480 861 -456
rect 861 -480 879 -456
rect 879 -480 884 -456
rect 1153 -455 1181 -450
rect 1336 -425 1364 -420
rect 1336 -449 1341 -425
rect 1341 -449 1359 -425
rect 1359 -449 1364 -425
rect 1336 -454 1364 -449
rect 1734 -458 1751 -70
rect 1863 -458 1880 -70
rect 1992 -458 2009 -70
rect 2121 -458 2138 -70
rect 2250 -458 2267 -70
rect 856 -485 884 -480
rect 595 -630 2055 -530
<< metal1 >>
rect 255 1070 2280 1100
rect 255 980 305 1070
rect 815 980 875 1070
rect 1380 980 1460 1070
rect 1970 980 2280 1070
rect 255 950 2280 980
rect 283 548 319 950
rect 283 518 286 548
rect 316 518 319 548
rect 283 512 319 518
rect 406 907 429 913
rect 332 383 358 386
rect 329 357 332 383
rect 358 357 360 383
rect 332 354 358 357
rect 406 119 409 907
rect 426 119 429 907
rect 406 113 429 119
rect 535 907 560 950
rect 665 913 685 930
rect 535 119 538 907
rect 555 900 560 907
rect 664 907 687 913
rect 555 119 558 900
rect 664 798 667 907
rect 684 798 687 907
rect 856 902 879 908
rect 659 772 662 798
rect 688 772 691 798
rect 603 136 606 164
rect 634 136 637 164
rect 535 113 558 119
rect 412 68 428 113
rect 606 80 634 136
rect 664 119 667 772
rect 684 119 687 772
rect 856 714 859 902
rect 876 714 879 902
rect 856 708 879 714
rect 985 902 1010 950
rect 985 714 988 902
rect 1005 895 1010 902
rect 1046 907 1069 913
rect 1005 714 1008 895
rect 985 708 1008 714
rect 917 669 951 675
rect 753 641 756 669
rect 784 641 920 669
rect 950 641 953 669
rect 917 635 951 641
rect 726 582 749 588
rect 726 194 729 582
rect 746 194 749 582
rect 726 188 749 194
rect 855 582 878 588
rect 855 194 858 582
rect 875 194 878 582
rect 855 188 878 194
rect 984 582 1007 588
rect 984 194 987 582
rect 1004 194 1007 582
rect 984 188 1007 194
rect 728 145 748 188
rect 793 149 827 155
rect 728 125 755 145
rect 793 143 796 149
rect 664 113 687 119
rect 674 88 705 91
rect 473 74 507 80
rect 473 68 476 74
rect 412 52 476 68
rect 412 -366 428 52
rect 473 46 476 52
rect 504 68 507 74
rect 603 74 637 80
rect 603 68 606 74
rect 504 52 606 68
rect 504 46 507 52
rect 473 40 507 46
rect 603 46 606 52
rect 634 46 637 74
rect 671 62 674 88
rect 705 85 708 88
rect 705 62 710 85
rect 671 60 677 62
rect 702 60 710 62
rect 671 57 710 60
rect 675 56 710 57
rect 603 40 637 46
rect 735 23 755 125
rect 790 122 796 143
rect 824 143 827 149
rect 918 149 952 155
rect 918 143 921 149
rect 824 122 830 143
rect 915 122 921 143
rect 793 116 796 122
rect 824 116 827 122
rect 793 110 827 116
rect 918 116 921 122
rect 949 143 952 149
rect 949 122 955 143
rect 949 116 952 122
rect 918 110 952 116
rect 1046 119 1049 907
rect 1066 119 1069 907
rect 1046 113 1069 119
rect 1175 907 1200 950
rect 1175 119 1178 907
rect 1195 900 1200 907
rect 1304 907 1327 913
rect 1195 119 1198 900
rect 1175 113 1198 119
rect 1304 119 1307 907
rect 1324 119 1327 907
rect 1386 907 1409 913
rect 1386 520 1389 907
rect 1385 519 1389 520
rect 1406 520 1409 907
rect 1515 907 1540 950
rect 1406 519 1410 520
rect 1385 417 1410 519
rect 1515 519 1518 907
rect 1535 890 1540 907
rect 1644 907 1667 913
rect 1535 519 1538 890
rect 1515 513 1538 519
rect 1644 519 1647 907
rect 1664 567 1667 907
rect 1730 906 1755 950
rect 1985 912 2010 950
rect 1730 895 1734 906
rect 1664 519 1670 567
rect 1644 513 1670 519
rect 1448 479 1482 480
rect 1444 476 1482 479
rect 1472 474 1488 476
rect 1479 468 1488 474
rect 1578 474 1612 480
rect 1578 468 1581 474
rect 1479 452 1581 468
rect 1479 447 1488 452
rect 1444 446 1451 447
rect 1479 446 1482 447
rect 1444 444 1482 446
rect 1448 440 1482 444
rect 1578 446 1581 452
rect 1609 468 1612 474
rect 1609 452 1615 468
rect 1609 446 1612 452
rect 1578 440 1612 446
rect 1645 422 1670 513
rect 1367 392 1410 417
rect 1572 397 1670 422
rect 1367 346 1392 392
rect 1572 346 1597 397
rect 1367 340 1394 346
rect 1367 203 1374 340
rect 1391 203 1394 340
rect 1393 177 1394 203
rect 1367 174 1374 177
rect 1371 152 1374 174
rect 1391 152 1394 177
rect 1371 146 1394 152
rect 1450 340 1473 346
rect 1450 152 1453 340
rect 1470 152 1473 340
rect 1572 340 1599 346
rect 1572 313 1579 340
rect 1596 313 1599 340
rect 1655 340 1678 346
rect 1569 287 1572 313
rect 1598 287 1601 313
rect 1450 146 1473 152
rect 1576 152 1579 287
rect 1596 152 1599 287
rect 1576 146 1599 152
rect 1655 152 1658 340
rect 1675 152 1678 340
rect 1655 146 1678 152
rect 1304 113 1327 119
rect 925 95 945 110
rect 848 89 883 95
rect 848 72 856 89
rect 873 72 883 89
rect 925 75 1035 95
rect 1052 77 1068 113
rect 848 66 883 72
rect 933 53 956 55
rect 653 17 676 23
rect 653 14 656 17
rect 649 11 656 14
rect 673 14 676 17
rect 732 17 755 23
rect 673 11 681 14
rect 544 0 547 6
rect 515 -20 547 0
rect 573 5 576 6
rect 573 -1 592 5
rect 582 -18 592 -1
rect 649 -15 652 11
rect 678 -15 681 11
rect 649 -18 656 -15
rect 573 -20 592 -18
rect 515 -57 535 -20
rect 558 -23 592 -20
rect 562 -24 585 -23
rect 207 -383 428 -366
rect 514 -63 537 -57
rect 207 -433 223 -383
rect 288 -410 336 -407
rect 201 -436 230 -433
rect 201 -453 207 -436
rect 224 -453 230 -436
rect 288 -446 294 -410
rect 330 -446 336 -410
rect 288 -449 336 -446
rect 437 -430 473 -424
rect 201 -456 230 -453
rect 294 -521 330 -449
rect 437 -460 440 -430
rect 470 -460 473 -430
rect 514 -451 517 -63
rect 534 -451 537 -63
rect 514 -457 537 -451
rect 593 -63 616 -57
rect 593 -451 596 -63
rect 613 -451 616 -63
rect 653 -171 656 -18
rect 673 -18 681 -15
rect 673 -171 676 -18
rect 732 -170 735 17
rect 653 -177 676 -171
rect 730 -171 735 -170
rect 752 -171 755 17
rect 812 27 835 33
rect 812 -67 815 27
rect 832 -67 835 27
rect 891 27 914 33
rect 929 27 932 53
rect 958 27 961 53
rect 809 -70 812 -67
rect 808 -90 812 -70
rect 809 -93 812 -90
rect 838 -93 841 -67
rect 812 -161 815 -93
rect 832 -161 835 -93
rect 812 -167 835 -161
rect 891 -161 894 27
rect 911 -150 914 27
rect 933 26 956 27
rect 968 6 1000 9
rect 968 -20 971 6
rect 997 -20 1000 6
rect 968 -23 1000 -20
rect 1015 5 1035 75
rect 1049 71 1072 77
rect 1049 54 1052 71
rect 1069 68 1072 71
rect 1108 74 1142 80
rect 1108 68 1111 74
rect 1069 54 1111 68
rect 1049 52 1111 54
rect 1049 48 1072 52
rect 1108 46 1111 52
rect 1139 68 1142 74
rect 1238 74 1272 80
rect 1305 79 1325 113
rect 1403 111 1437 115
rect 1403 109 1438 111
rect 1403 103 1406 109
rect 1434 108 1438 109
rect 1400 82 1406 103
rect 1603 109 1637 115
rect 1603 105 1606 109
rect 1438 82 1606 105
rect 1238 68 1241 74
rect 1139 52 1241 68
rect 1139 46 1142 52
rect 1108 40 1142 46
rect 1238 46 1241 52
rect 1269 46 1272 74
rect 1303 73 1326 79
rect 1303 56 1306 73
rect 1323 56 1326 73
rect 1403 76 1406 82
rect 1434 80 1606 82
rect 1434 79 1438 80
rect 1434 76 1437 79
rect 1403 70 1437 76
rect 1603 76 1606 80
rect 1634 103 1637 109
rect 1634 82 1640 103
rect 1634 76 1637 82
rect 1603 70 1637 76
rect 1303 50 1326 56
rect 1238 40 1272 46
rect 1655 35 1675 146
rect 1731 118 1734 895
rect 1751 895 1755 906
rect 1860 906 1883 912
rect 1751 118 1754 895
rect 1731 112 1754 118
rect 1860 118 1863 906
rect 1880 125 1883 906
rect 1985 906 2012 912
rect 1985 900 1992 906
rect 1880 118 1885 125
rect 1788 74 1822 80
rect 1788 68 1791 74
rect 1785 47 1791 68
rect 1788 41 1791 47
rect 1819 68 1822 74
rect 1860 68 1885 118
rect 1989 118 1992 900
rect 2009 118 2012 906
rect 2118 906 2141 912
rect 2118 132 2121 906
rect 1989 112 2012 118
rect 2117 118 2121 132
rect 2138 132 2141 906
rect 2245 906 2270 950
rect 2245 900 2250 906
rect 2138 118 2142 132
rect 1918 74 1952 80
rect 1918 68 1921 74
rect 1819 47 1825 68
rect 1819 41 1822 47
rect 1856 42 1859 68
rect 1885 42 1888 68
rect 1915 47 1921 68
rect 1788 35 1822 41
rect 1273 12 1296 18
rect 1138 5 1164 10
rect 1015 4 1164 5
rect 1015 -13 1141 4
rect 1158 -13 1164 4
rect 1015 -15 1164 -13
rect 1015 -25 1035 -15
rect 1138 -19 1164 -15
rect 1097 -37 1123 -34
rect 1217 -37 1243 -34
rect 1123 -60 1217 -40
rect 1097 -66 1123 -63
rect 1217 -66 1243 -63
rect 1152 -92 1178 -89
rect 952 -117 1152 -92
rect 911 -161 915 -150
rect 730 -217 755 -171
rect 730 -223 756 -217
rect 730 -230 736 -223
rect 733 -411 736 -230
rect 753 -411 756 -223
rect 733 -417 756 -411
rect 812 -223 835 -217
rect 812 -411 815 -223
rect 832 -411 835 -223
rect 812 -417 835 -411
rect 891 -223 915 -161
rect 952 -193 977 -117
rect 1152 -121 1178 -118
rect 1273 -137 1276 12
rect 1080 -162 1276 -137
rect 1080 -190 1105 -162
rect 952 -212 956 -193
rect 891 -411 894 -223
rect 911 -228 915 -223
rect 911 -411 914 -228
rect 953 -381 956 -212
rect 973 -212 977 -193
rect 1082 -193 1105 -190
rect 973 -381 976 -212
rect 1012 -282 1038 -279
rect 1009 -308 1012 -282
rect 1038 -308 1041 -282
rect 1012 -311 1038 -308
rect 953 -387 976 -381
rect 1082 -381 1085 -193
rect 1102 -381 1105 -193
rect 1211 -193 1234 -187
rect 1211 -207 1214 -193
rect 1231 -207 1234 -193
rect 1209 -233 1212 -207
rect 1238 -233 1241 -207
rect 1157 -352 1183 -349
rect 1154 -378 1157 -352
rect 1183 -378 1186 -352
rect 1157 -381 1183 -378
rect 1211 -381 1214 -233
rect 1231 -287 1237 -233
rect 1231 -381 1234 -287
rect 1082 -387 1105 -381
rect 1211 -387 1234 -381
rect 1273 -376 1276 -162
rect 1293 -376 1296 12
rect 1402 12 1425 18
rect 1317 -37 1343 -34
rect 1314 -63 1317 -37
rect 1343 -63 1346 -37
rect 1317 -66 1343 -63
rect 1402 -357 1405 12
rect 1273 -382 1296 -376
rect 1400 -376 1405 -357
rect 1422 -376 1425 12
rect 1630 15 1675 35
rect 1630 -5 1650 15
rect 1792 -1 1818 1
rect 1788 -5 1823 -1
rect 1630 -25 1795 -5
rect 1815 -25 1823 -5
rect 1517 -37 1543 -34
rect 1543 -63 1546 -37
rect 1517 -66 1543 -63
rect 1507 -116 1542 -110
rect 1507 -122 1510 -116
rect 1505 -143 1510 -122
rect 1507 -149 1510 -143
rect 1539 -120 1542 -116
rect 1572 -116 1607 -110
rect 1572 -120 1575 -116
rect 1539 -145 1575 -120
rect 1539 -149 1542 -145
rect 1507 -155 1542 -149
rect 1572 -149 1575 -145
rect 1604 -122 1607 -116
rect 1604 -143 1610 -122
rect 1604 -149 1607 -143
rect 1572 -155 1607 -149
rect 1630 -187 1650 -25
rect 1788 -30 1823 -25
rect 1792 -31 1818 -30
rect 891 -417 914 -411
rect 593 -457 616 -451
rect 657 -452 683 -449
rect 437 -466 473 -460
rect 440 -521 470 -466
rect 595 -505 615 -457
rect 758 -451 792 -445
rect 758 -455 761 -451
rect 683 -475 761 -455
rect 657 -481 683 -478
rect 755 -479 761 -475
rect 758 -485 761 -479
rect 789 -457 792 -451
rect 789 -479 795 -457
rect 789 -485 792 -479
rect 758 -491 792 -485
rect 815 -505 835 -417
rect 1008 -421 1042 -415
rect 1008 -427 1011 -421
rect 853 -451 887 -445
rect 1005 -448 1011 -427
rect 853 -457 856 -451
rect 850 -479 856 -457
rect 853 -485 856 -479
rect 884 -453 887 -451
rect 962 -451 988 -448
rect 884 -475 962 -453
rect 884 -479 890 -475
rect 1008 -454 1011 -448
rect 1039 -427 1042 -421
rect 1150 -422 1184 -416
rect 1039 -448 1045 -427
rect 1150 -428 1153 -422
rect 1039 -454 1042 -448
rect 1147 -449 1153 -428
rect 1008 -460 1042 -454
rect 1150 -455 1153 -449
rect 1181 -428 1184 -422
rect 1333 -420 1367 -414
rect 1181 -449 1187 -428
rect 1181 -455 1184 -449
rect 1254 -450 1257 -424
rect 1283 -426 1286 -424
rect 1333 -426 1336 -420
rect 1283 -448 1336 -426
rect 1283 -450 1286 -448
rect 1150 -461 1184 -455
rect 1333 -454 1336 -448
rect 1364 -426 1367 -420
rect 1364 -448 1370 -426
rect 1364 -454 1367 -448
rect 1333 -460 1367 -454
rect 884 -485 887 -479
rect 962 -480 988 -477
rect 853 -491 887 -485
rect 1400 -505 1425 -376
rect 1468 -193 1491 -187
rect 1468 -381 1471 -193
rect 1488 -381 1491 -193
rect 1547 -193 1570 -187
rect 1547 -380 1550 -193
rect 1468 -387 1491 -381
rect 1545 -381 1550 -380
rect 1567 -381 1570 -193
rect 1545 -505 1570 -381
rect 1626 -193 1650 -187
rect 1626 -381 1629 -193
rect 1646 -215 1650 -193
rect 1731 -70 1754 -64
rect 1646 -381 1649 -215
rect 1626 -387 1649 -381
rect 1731 -413 1734 -70
rect 1730 -458 1734 -413
rect 1751 -413 1754 -70
rect 1860 -70 1885 42
rect 1918 41 1921 47
rect 1949 68 1952 74
rect 2048 74 2082 80
rect 2048 68 2051 74
rect 1949 47 1955 68
rect 2045 47 2051 68
rect 1949 41 1952 47
rect 1918 35 1952 41
rect 2048 41 2051 47
rect 2079 68 2082 74
rect 2117 68 2142 118
rect 2247 118 2250 900
rect 2267 118 2270 906
rect 2247 112 2270 118
rect 2173 74 2207 80
rect 2173 68 2176 74
rect 2079 47 2085 68
rect 2079 41 2082 47
rect 2114 42 2117 68
rect 2143 42 2146 68
rect 2170 47 2176 68
rect 2048 35 2082 41
rect 1922 -8 1956 -1
rect 1922 -25 1929 -8
rect 1946 -25 1956 -8
rect 1922 -30 1956 -25
rect 2048 -8 2083 -1
rect 2048 -25 2056 -8
rect 2073 -25 2083 -8
rect 2048 -30 2083 -25
rect 1926 -31 1949 -30
rect 2053 -31 2076 -30
rect 2120 -64 2145 42
rect 2173 41 2176 47
rect 2204 68 2207 74
rect 2204 47 2210 68
rect 2204 41 2207 47
rect 2173 35 2207 41
rect 2180 -8 2214 -1
rect 2180 -25 2187 -8
rect 2204 -25 2214 -8
rect 2180 -30 2214 -25
rect 2184 -31 2207 -30
rect 1860 -282 1863 -70
rect 1880 -282 1885 -70
rect 1989 -70 2012 -64
rect 1859 -308 1862 -282
rect 1888 -308 1891 -282
rect 1751 -458 1755 -413
rect 1730 -505 1755 -458
rect 1860 -458 1863 -308
rect 1880 -458 1883 -308
rect 1860 -464 1883 -458
rect 1989 -458 1992 -70
rect 2009 -408 2012 -70
rect 2118 -70 2145 -64
rect 2009 -458 2015 -408
rect 1989 -464 2015 -458
rect 2118 -458 2121 -70
rect 2138 -75 2145 -70
rect 2247 -70 2270 -64
rect 2138 -458 2141 -75
rect 2247 -393 2250 -70
rect 2118 -464 2141 -458
rect 2245 -458 2250 -393
rect 2267 -458 2270 -70
rect 1990 -505 2015 -464
rect 535 -521 2100 -505
rect 294 -527 2100 -521
rect 2245 -527 2270 -458
rect 294 -530 2270 -527
rect 294 -557 595 -530
rect 535 -630 595 -557
rect 2055 -552 2270 -530
rect 2055 -630 2100 -552
rect 535 -655 2100 -630
<< via1 >>
rect 305 980 815 1070
rect 875 980 1380 1070
rect 1460 980 1970 1070
rect 332 380 358 383
rect 332 360 335 380
rect 335 360 354 380
rect 354 360 358 380
rect 332 357 358 360
rect 662 772 667 798
rect 667 772 684 798
rect 684 772 688 798
rect 606 136 634 164
rect 756 641 784 669
rect 921 641 948 669
rect 948 641 950 669
rect 674 85 705 88
rect 674 62 677 85
rect 677 62 702 85
rect 702 62 705 85
rect 797 122 823 148
rect 1444 474 1472 476
rect 1444 447 1451 474
rect 1451 447 1472 474
rect 1367 177 1374 203
rect 1374 177 1391 203
rect 1391 177 1393 203
rect 1572 287 1579 313
rect 1579 287 1596 313
rect 1596 287 1598 313
rect 547 -1 573 6
rect 547 -18 565 -1
rect 565 -18 573 -1
rect 652 -15 656 11
rect 656 -15 673 11
rect 673 -15 678 11
rect 547 -20 573 -18
rect 932 49 958 53
rect 932 32 936 49
rect 936 32 953 49
rect 953 32 958 49
rect 932 27 958 32
rect 812 -93 815 -67
rect 815 -93 832 -67
rect 832 -93 838 -67
rect 971 2 997 6
rect 971 -17 974 2
rect 974 -17 994 2
rect 994 -17 997 2
rect 971 -20 997 -17
rect 1412 82 1434 108
rect 1434 82 1438 108
rect 1859 42 1885 68
rect 1097 -63 1123 -37
rect 1217 -63 1243 -37
rect 1152 -118 1178 -92
rect 1012 -285 1038 -282
rect 1012 -305 1015 -285
rect 1015 -305 1035 -285
rect 1035 -305 1038 -285
rect 1012 -308 1038 -305
rect 1212 -233 1214 -207
rect 1214 -233 1231 -207
rect 1231 -233 1238 -207
rect 1157 -355 1183 -352
rect 1157 -375 1160 -355
rect 1160 -375 1180 -355
rect 1180 -375 1183 -355
rect 1157 -378 1183 -375
rect 1317 -40 1343 -37
rect 1317 -60 1320 -40
rect 1320 -60 1340 -40
rect 1340 -60 1343 -40
rect 1317 -63 1343 -60
rect 1517 -40 1543 -37
rect 1517 -60 1523 -40
rect 1523 -60 1540 -40
rect 1540 -60 1543 -40
rect 1517 -63 1543 -60
rect 657 -478 683 -452
rect 962 -477 988 -451
rect 1257 -450 1283 -424
rect 2117 42 2143 68
rect 1862 -308 1863 -282
rect 1863 -308 1880 -282
rect 1880 -308 1888 -282
rect 595 -630 2055 -530
<< metal2 >>
rect 255 1070 2020 1100
rect 255 980 305 1070
rect 815 980 875 1070
rect 1380 980 1460 1070
rect 1970 980 2020 1070
rect 255 950 2020 980
rect 461 826 1540 851
rect 461 383 486 826
rect 662 798 688 801
rect 329 357 332 383
rect 358 358 486 383
rect 550 775 662 795
rect 358 357 361 358
rect 550 9 570 775
rect 662 769 688 772
rect 756 669 784 672
rect 606 641 756 669
rect 606 164 634 641
rect 756 638 784 641
rect 921 669 950 672
rect 950 641 1472 669
rect 921 638 950 641
rect 1444 476 1472 641
rect 1441 447 1444 476
rect 1472 447 1475 476
rect 1515 391 1540 826
rect 1412 366 1540 391
rect 1412 292 1437 366
rect 606 133 634 136
rect 677 267 1437 292
rect 677 88 702 267
rect 1364 177 1367 203
rect 1393 177 1396 203
rect 794 122 797 148
rect 823 145 826 148
rect 823 125 994 145
rect 823 122 826 125
rect 671 62 674 88
rect 705 62 708 88
rect 932 55 958 56
rect 930 53 960 55
rect 930 47 932 53
rect 657 30 932 47
rect 657 14 680 30
rect 930 27 932 30
rect 958 27 960 53
rect 930 25 960 27
rect 932 24 958 25
rect 649 11 681 14
rect 547 6 573 9
rect 573 -20 630 0
rect 649 -15 652 11
rect 678 -15 681 11
rect 974 9 994 125
rect 1367 17 1392 177
rect 1412 108 1437 267
rect 1572 313 1598 316
rect 1572 284 1598 287
rect 1409 82 1412 108
rect 1438 82 1441 108
rect 649 -18 681 -15
rect 968 6 1000 9
rect 547 -23 573 -20
rect 610 -250 630 -20
rect 968 -20 971 6
rect 997 -20 1000 6
rect 968 -23 1000 -20
rect 1152 -7 1392 17
rect 1094 -40 1097 -37
rect 940 -60 1097 -40
rect 812 -67 838 -64
rect 940 -70 960 -60
rect 1094 -63 1097 -60
rect 1123 -63 1126 -37
rect 838 -90 960 -70
rect 1152 -92 1177 -7
rect 1317 -37 1343 -34
rect 1214 -63 1217 -37
rect 1243 -40 1246 -37
rect 1243 -60 1317 -40
rect 1243 -63 1246 -60
rect 1514 -40 1517 -37
rect 1343 -60 1517 -40
rect 1514 -63 1517 -60
rect 1543 -63 1546 -37
rect 1317 -66 1343 -63
rect 812 -96 838 -93
rect 1149 -118 1152 -92
rect 1178 -118 1181 -92
rect 1572 -123 1597 284
rect 1859 68 1885 71
rect 2117 68 2143 71
rect 1885 42 2117 67
rect 2143 42 2270 67
rect 1859 39 1885 42
rect 2117 39 2143 42
rect 2245 24 2270 42
rect 2245 0 2344 24
rect 1212 -148 1597 -123
rect 1212 -204 1237 -148
rect 1212 -207 1238 -204
rect 1212 -236 1238 -233
rect 610 -270 680 -250
rect 660 -452 680 -270
rect 1012 -282 1038 -279
rect 1862 -282 1888 -279
rect 1038 -305 1862 -285
rect 1012 -311 1038 -308
rect 1862 -311 1888 -308
rect 1157 -352 1183 -349
rect 1183 -375 2348 -355
rect 1157 -381 1183 -378
rect 1257 -424 1283 -421
rect 1094 -447 1257 -426
rect 654 -478 657 -452
rect 683 -478 686 -452
rect 959 -477 962 -451
rect 988 -454 991 -451
rect 1094 -454 1116 -447
rect 1257 -453 1283 -450
rect 988 -475 1116 -454
rect 988 -477 991 -475
rect 535 -530 2100 -505
rect 535 -630 595 -530
rect 2055 -630 2100 -530
rect 535 -655 2100 -630
<< via2 >>
rect 305 980 815 1070
rect 875 980 1380 1070
rect 1460 980 1970 1070
rect 595 -630 2055 -530
<< metal3 >>
rect 136 1070 2370 1100
rect 136 980 305 1070
rect 815 980 875 1070
rect 1380 980 1460 1070
rect 1970 980 2370 1070
rect 136 950 2370 980
rect 136 -530 2370 -505
rect 136 -630 595 -530
rect 2055 -630 2370 -530
rect 136 -655 2370 -630
<< labels >>
flabel metal3 s 170 -595 170 -595 0 FreeSans 320 0 0 0 VSSA
flabel metal2 s 2334 -366 2334 -366 0 FreeSans 400 0 0 0 VIN
flabel metal2 s 2330 13 2330 13 0 FreeSans 400 0 0 0 VOUT
flabel metal3 s 195 1031 195 1031 0 FreeSans 320 0 0 0 VDDA
<< end >>
