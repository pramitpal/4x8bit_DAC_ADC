magic
tech sky130A
magscale 1 2
timestamp 1687970707
<< nwell >>
rect 1162 2140 1828 2346
rect 3260 2328 4174 2336
rect 5504 2328 6132 2336
rect 3260 2140 4866 2328
rect 1162 2068 4866 2140
rect 1210 1816 4866 2068
rect 5504 1816 6824 2328
rect 1210 1808 3362 1816
rect 1210 1806 3290 1808
rect 2714 1802 3028 1806
rect 1162 912 1828 1118
rect 3260 1100 4174 1108
rect 3260 912 4866 1100
rect 1162 840 4866 912
rect 1210 588 4866 840
rect 1210 580 3362 588
rect 1210 578 3290 580
rect 2714 574 3028 578
<< pwell >>
rect 690 2194 980 2200
rect 400 1522 980 2194
rect 4246 1770 4822 1772
rect 6204 1770 6780 1772
rect 1254 1608 3232 1760
rect 3586 1620 4822 1770
rect 5544 1620 6780 1770
rect 3586 1618 4162 1620
rect 5544 1618 6120 1620
rect 3586 1614 4152 1618
rect 5544 1614 6110 1618
rect 1254 1602 1867 1608
rect 400 1516 682 1522
rect 1180 1422 1867 1602
rect 3560 1422 4152 1614
rect 5518 1422 6110 1614
rect 690 966 980 972
rect 400 294 980 966
rect 4246 542 4822 544
rect 1254 380 3232 532
rect 3586 392 4822 542
rect 3586 390 4162 392
rect 3586 386 4152 390
rect 1254 374 1867 380
rect 400 288 682 294
rect 1180 194 1867 374
rect 3560 194 4152 386
<< mvnmos >>
rect 1338 1634 1438 1734
rect 1626 1634 1726 1734
rect 1958 1634 2058 1734
rect 2300 1634 2400 1734
rect 2704 1634 2804 1734
rect 3048 1634 3148 1734
rect 3670 1644 3770 1744
rect 3978 1644 4078 1744
rect 4330 1646 4430 1746
rect 4638 1646 4738 1746
rect 5628 1644 5728 1744
rect 5936 1644 6036 1744
rect 6288 1646 6388 1746
rect 6596 1646 6696 1746
rect 1338 406 1438 506
rect 1626 406 1726 506
rect 1958 406 2058 506
rect 2300 406 2400 506
rect 2704 406 2804 506
rect 3048 406 3148 506
rect 3670 416 3770 516
rect 3978 416 4078 516
rect 4330 418 4430 518
rect 4638 418 4738 518
<< mvpmos >>
rect 1338 1872 1438 2072
rect 1626 1872 1726 2072
rect 1958 1872 2058 2072
rect 2300 1872 2400 2072
rect 2704 1872 2804 2072
rect 3048 1872 3148 2072
rect 3670 1882 3770 2082
rect 3978 1882 4078 2082
rect 4330 1882 4430 2082
rect 4638 1882 4738 2082
rect 5628 1882 5728 2082
rect 5936 1882 6036 2082
rect 6288 1882 6388 2082
rect 6596 1882 6696 2082
rect 1338 644 1438 844
rect 1626 644 1726 844
rect 1958 644 2058 844
rect 2300 644 2400 844
rect 2704 644 2804 844
rect 3048 644 3148 844
rect 3670 654 3770 854
rect 3978 654 4078 854
rect 4330 654 4430 854
rect 4638 654 4738 854
<< mvndiff >>
rect 426 2156 510 2168
rect 426 2122 451 2156
rect 485 2122 510 2156
rect 426 2065 510 2122
rect 426 1588 510 1645
rect 426 1554 451 1588
rect 485 1554 510 1588
rect 426 1542 510 1554
rect 572 2156 656 2168
rect 572 2122 597 2156
rect 631 2122 656 2156
rect 572 2065 656 2122
rect 572 1588 656 1645
rect 572 1554 597 1588
rect 631 1554 656 1588
rect 572 1542 656 1554
rect 716 2162 800 2174
rect 716 2128 741 2162
rect 775 2128 800 2162
rect 716 2071 800 2128
rect 716 1594 800 1651
rect 716 1560 741 1594
rect 775 1560 800 1594
rect 716 1548 800 1560
rect 870 2162 954 2174
rect 870 2128 895 2162
rect 929 2128 954 2162
rect 870 2071 954 2128
rect 870 1594 954 1651
rect 1280 1701 1338 1734
rect 1280 1667 1292 1701
rect 1326 1667 1338 1701
rect 1280 1634 1338 1667
rect 1438 1701 1496 1734
rect 1438 1667 1450 1701
rect 1484 1667 1496 1701
rect 1438 1634 1496 1667
rect 1568 1701 1626 1734
rect 1568 1667 1580 1701
rect 1614 1667 1626 1701
rect 1568 1634 1626 1667
rect 1726 1701 1784 1734
rect 1726 1667 1738 1701
rect 1772 1667 1784 1701
rect 1726 1634 1784 1667
rect 1900 1701 1958 1734
rect 1900 1667 1912 1701
rect 1946 1667 1958 1701
rect 1900 1634 1958 1667
rect 2058 1701 2116 1734
rect 2058 1667 2070 1701
rect 2104 1667 2116 1701
rect 2058 1634 2116 1667
rect 2242 1701 2300 1734
rect 2242 1667 2254 1701
rect 2288 1667 2300 1701
rect 2242 1634 2300 1667
rect 2400 1701 2458 1734
rect 2400 1667 2412 1701
rect 2446 1667 2458 1701
rect 2400 1634 2458 1667
rect 2646 1701 2704 1734
rect 2646 1667 2658 1701
rect 2692 1667 2704 1701
rect 2646 1634 2704 1667
rect 2804 1701 2862 1734
rect 2804 1667 2816 1701
rect 2850 1667 2862 1701
rect 2804 1634 2862 1667
rect 2990 1701 3048 1734
rect 2990 1667 3002 1701
rect 3036 1667 3048 1701
rect 2990 1634 3048 1667
rect 3148 1701 3206 1734
rect 3148 1667 3160 1701
rect 3194 1667 3206 1701
rect 3148 1634 3206 1667
rect 3612 1711 3670 1744
rect 3612 1677 3624 1711
rect 3658 1677 3670 1711
rect 3612 1644 3670 1677
rect 3770 1711 3828 1744
rect 3770 1677 3782 1711
rect 3816 1677 3828 1711
rect 3770 1644 3828 1677
rect 3920 1711 3978 1744
rect 3920 1677 3932 1711
rect 3966 1677 3978 1711
rect 3920 1644 3978 1677
rect 4078 1711 4136 1744
rect 4078 1677 4090 1711
rect 4124 1677 4136 1711
rect 4078 1644 4136 1677
rect 4272 1713 4330 1746
rect 4272 1679 4284 1713
rect 4318 1679 4330 1713
rect 4272 1646 4330 1679
rect 4430 1713 4488 1746
rect 4430 1679 4442 1713
rect 4476 1679 4488 1713
rect 4430 1646 4488 1679
rect 4580 1713 4638 1746
rect 4580 1679 4592 1713
rect 4626 1679 4638 1713
rect 4580 1646 4638 1679
rect 4738 1713 4796 1746
rect 4738 1679 4750 1713
rect 4784 1679 4796 1713
rect 4738 1646 4796 1679
rect 5570 1712 5628 1744
rect 5570 1678 5582 1712
rect 5616 1678 5628 1712
rect 5570 1644 5628 1678
rect 5728 1712 5786 1744
rect 5728 1678 5740 1712
rect 5774 1678 5786 1712
rect 5728 1644 5786 1678
rect 5878 1712 5936 1744
rect 5878 1678 5890 1712
rect 5924 1678 5936 1712
rect 5878 1644 5936 1678
rect 6036 1712 6094 1744
rect 6036 1678 6048 1712
rect 6082 1678 6094 1712
rect 6036 1644 6094 1678
rect 6230 1714 6288 1746
rect 6230 1680 6242 1714
rect 6276 1680 6288 1714
rect 6230 1646 6288 1680
rect 6388 1714 6446 1746
rect 6388 1680 6400 1714
rect 6434 1680 6446 1714
rect 6388 1646 6446 1680
rect 6538 1714 6596 1746
rect 6538 1680 6550 1714
rect 6584 1680 6596 1714
rect 6538 1646 6596 1680
rect 6696 1714 6754 1746
rect 6696 1680 6708 1714
rect 6742 1680 6754 1714
rect 6696 1646 6754 1680
rect 870 1560 895 1594
rect 929 1560 954 1594
rect 870 1548 954 1560
rect 426 928 510 940
rect 426 894 451 928
rect 485 894 510 928
rect 426 837 510 894
rect 426 360 510 417
rect 426 326 451 360
rect 485 326 510 360
rect 426 314 510 326
rect 572 928 656 940
rect 572 894 597 928
rect 631 894 656 928
rect 572 837 656 894
rect 572 360 656 417
rect 572 326 597 360
rect 631 326 656 360
rect 572 314 656 326
rect 716 934 800 946
rect 716 900 741 934
rect 775 900 800 934
rect 716 843 800 900
rect 716 366 800 423
rect 716 332 741 366
rect 775 332 800 366
rect 716 320 800 332
rect 870 934 954 946
rect 870 900 895 934
rect 929 900 954 934
rect 870 843 954 900
rect 870 366 954 423
rect 1280 473 1338 506
rect 1280 439 1292 473
rect 1326 439 1338 473
rect 1280 406 1338 439
rect 1438 473 1496 506
rect 1438 439 1450 473
rect 1484 439 1496 473
rect 1438 406 1496 439
rect 1568 473 1626 506
rect 1568 439 1580 473
rect 1614 439 1626 473
rect 1568 406 1626 439
rect 1726 473 1784 506
rect 1726 439 1738 473
rect 1772 439 1784 473
rect 1726 406 1784 439
rect 1900 473 1958 506
rect 1900 439 1912 473
rect 1946 439 1958 473
rect 1900 406 1958 439
rect 2058 473 2116 506
rect 2058 439 2070 473
rect 2104 439 2116 473
rect 2058 406 2116 439
rect 2242 473 2300 506
rect 2242 439 2254 473
rect 2288 439 2300 473
rect 2242 406 2300 439
rect 2400 473 2458 506
rect 2400 439 2412 473
rect 2446 439 2458 473
rect 2400 406 2458 439
rect 2646 473 2704 506
rect 2646 439 2658 473
rect 2692 439 2704 473
rect 2646 406 2704 439
rect 2804 473 2862 506
rect 2804 439 2816 473
rect 2850 439 2862 473
rect 2804 406 2862 439
rect 2990 473 3048 506
rect 2990 439 3002 473
rect 3036 439 3048 473
rect 2990 406 3048 439
rect 3148 473 3206 506
rect 3148 439 3160 473
rect 3194 439 3206 473
rect 3148 406 3206 439
rect 3612 483 3670 516
rect 3612 449 3624 483
rect 3658 449 3670 483
rect 3612 416 3670 449
rect 3770 483 3828 516
rect 3770 449 3782 483
rect 3816 449 3828 483
rect 3770 416 3828 449
rect 3920 483 3978 516
rect 3920 449 3932 483
rect 3966 449 3978 483
rect 3920 416 3978 449
rect 4078 483 4136 516
rect 4078 449 4090 483
rect 4124 449 4136 483
rect 4078 416 4136 449
rect 4272 485 4330 518
rect 4272 451 4284 485
rect 4318 451 4330 485
rect 4272 418 4330 451
rect 4430 485 4488 518
rect 4430 451 4442 485
rect 4476 451 4488 485
rect 4430 418 4488 451
rect 4580 485 4638 518
rect 4580 451 4592 485
rect 4626 451 4638 485
rect 4580 418 4638 451
rect 4738 485 4796 518
rect 4738 451 4750 485
rect 4784 451 4796 485
rect 4738 418 4796 451
rect 870 332 895 366
rect 929 332 954 366
rect 870 320 954 332
<< mvpdiff >>
rect 1280 2057 1338 2072
rect 1280 2023 1292 2057
rect 1326 2023 1338 2057
rect 1280 1989 1338 2023
rect 1280 1955 1292 1989
rect 1326 1955 1338 1989
rect 1280 1921 1338 1955
rect 1280 1887 1292 1921
rect 1326 1887 1338 1921
rect 1280 1872 1338 1887
rect 1438 2057 1496 2072
rect 1438 2023 1450 2057
rect 1484 2023 1496 2057
rect 1438 1989 1496 2023
rect 1438 1955 1450 1989
rect 1484 1955 1496 1989
rect 1438 1921 1496 1955
rect 1438 1887 1450 1921
rect 1484 1887 1496 1921
rect 1438 1872 1496 1887
rect 1568 2057 1626 2072
rect 1568 2023 1580 2057
rect 1614 2023 1626 2057
rect 1568 1989 1626 2023
rect 1568 1955 1580 1989
rect 1614 1955 1626 1989
rect 1568 1921 1626 1955
rect 1568 1887 1580 1921
rect 1614 1887 1626 1921
rect 1568 1872 1626 1887
rect 1726 2057 1784 2072
rect 1726 2023 1738 2057
rect 1772 2023 1784 2057
rect 1726 1989 1784 2023
rect 1726 1955 1738 1989
rect 1772 1955 1784 1989
rect 1726 1921 1784 1955
rect 1726 1887 1738 1921
rect 1772 1887 1784 1921
rect 1726 1872 1784 1887
rect 1900 2057 1958 2072
rect 1900 2023 1912 2057
rect 1946 2023 1958 2057
rect 1900 1989 1958 2023
rect 1900 1955 1912 1989
rect 1946 1955 1958 1989
rect 1900 1921 1958 1955
rect 1900 1887 1912 1921
rect 1946 1887 1958 1921
rect 1900 1872 1958 1887
rect 2058 2057 2116 2072
rect 2058 2023 2070 2057
rect 2104 2023 2116 2057
rect 2058 1989 2116 2023
rect 2058 1955 2070 1989
rect 2104 1955 2116 1989
rect 2058 1921 2116 1955
rect 2058 1887 2070 1921
rect 2104 1887 2116 1921
rect 2058 1872 2116 1887
rect 2242 2057 2300 2072
rect 2242 2023 2254 2057
rect 2288 2023 2300 2057
rect 2242 1989 2300 2023
rect 2242 1955 2254 1989
rect 2288 1955 2300 1989
rect 2242 1921 2300 1955
rect 2242 1887 2254 1921
rect 2288 1887 2300 1921
rect 2242 1872 2300 1887
rect 2400 2057 2458 2072
rect 2400 2023 2412 2057
rect 2446 2023 2458 2057
rect 2400 1989 2458 2023
rect 2400 1955 2412 1989
rect 2446 1955 2458 1989
rect 2400 1921 2458 1955
rect 2400 1887 2412 1921
rect 2446 1887 2458 1921
rect 2400 1872 2458 1887
rect 2646 2057 2704 2072
rect 2646 2023 2658 2057
rect 2692 2023 2704 2057
rect 2646 1989 2704 2023
rect 2646 1955 2658 1989
rect 2692 1955 2704 1989
rect 2646 1921 2704 1955
rect 2646 1887 2658 1921
rect 2692 1887 2704 1921
rect 2646 1872 2704 1887
rect 2804 2057 2862 2072
rect 2804 2023 2816 2057
rect 2850 2023 2862 2057
rect 2804 1989 2862 2023
rect 2804 1955 2816 1989
rect 2850 1955 2862 1989
rect 2804 1921 2862 1955
rect 2804 1887 2816 1921
rect 2850 1887 2862 1921
rect 2804 1872 2862 1887
rect 2990 2057 3048 2072
rect 2990 2023 3002 2057
rect 3036 2023 3048 2057
rect 2990 1989 3048 2023
rect 2990 1955 3002 1989
rect 3036 1955 3048 1989
rect 2990 1921 3048 1955
rect 2990 1887 3002 1921
rect 3036 1887 3048 1921
rect 2990 1872 3048 1887
rect 3148 2057 3206 2072
rect 3148 2023 3160 2057
rect 3194 2023 3206 2057
rect 3148 1989 3206 2023
rect 3148 1955 3160 1989
rect 3194 1955 3206 1989
rect 3148 1921 3206 1955
rect 3148 1887 3160 1921
rect 3194 1887 3206 1921
rect 3148 1872 3206 1887
rect 3612 2067 3670 2082
rect 3612 2033 3624 2067
rect 3658 2033 3670 2067
rect 3612 1999 3670 2033
rect 3612 1965 3624 1999
rect 3658 1965 3670 1999
rect 3612 1931 3670 1965
rect 3612 1897 3624 1931
rect 3658 1897 3670 1931
rect 3612 1882 3670 1897
rect 3770 2067 3828 2082
rect 3770 2033 3782 2067
rect 3816 2033 3828 2067
rect 3770 1999 3828 2033
rect 3770 1965 3782 1999
rect 3816 1965 3828 1999
rect 3770 1931 3828 1965
rect 3770 1897 3782 1931
rect 3816 1897 3828 1931
rect 3770 1882 3828 1897
rect 3920 2067 3978 2082
rect 3920 2033 3932 2067
rect 3966 2033 3978 2067
rect 3920 1999 3978 2033
rect 3920 1965 3932 1999
rect 3966 1965 3978 1999
rect 3920 1931 3978 1965
rect 3920 1897 3932 1931
rect 3966 1897 3978 1931
rect 3920 1882 3978 1897
rect 4078 2067 4136 2082
rect 4078 2033 4090 2067
rect 4124 2033 4136 2067
rect 4078 1999 4136 2033
rect 4078 1965 4090 1999
rect 4124 1965 4136 1999
rect 4078 1931 4136 1965
rect 4078 1897 4090 1931
rect 4124 1897 4136 1931
rect 4078 1882 4136 1897
rect 4272 2067 4330 2082
rect 4272 2033 4284 2067
rect 4318 2033 4330 2067
rect 4272 1999 4330 2033
rect 4272 1965 4284 1999
rect 4318 1965 4330 1999
rect 4272 1931 4330 1965
rect 4272 1897 4284 1931
rect 4318 1897 4330 1931
rect 4272 1882 4330 1897
rect 4430 2067 4488 2082
rect 4430 2033 4442 2067
rect 4476 2033 4488 2067
rect 4430 1999 4488 2033
rect 4430 1965 4442 1999
rect 4476 1965 4488 1999
rect 4430 1931 4488 1965
rect 4430 1897 4442 1931
rect 4476 1897 4488 1931
rect 4430 1882 4488 1897
rect 4580 2067 4638 2082
rect 4580 2033 4592 2067
rect 4626 2033 4638 2067
rect 4580 1999 4638 2033
rect 4580 1965 4592 1999
rect 4626 1965 4638 1999
rect 4580 1931 4638 1965
rect 4580 1897 4592 1931
rect 4626 1897 4638 1931
rect 4580 1882 4638 1897
rect 4738 2067 4796 2082
rect 4738 2033 4750 2067
rect 4784 2033 4796 2067
rect 4738 1999 4796 2033
rect 4738 1965 4750 1999
rect 4784 1965 4796 1999
rect 4738 1931 4796 1965
rect 4738 1897 4750 1931
rect 4784 1897 4796 1931
rect 4738 1882 4796 1897
rect 5570 2068 5628 2082
rect 5570 2034 5582 2068
rect 5616 2034 5628 2068
rect 5570 2000 5628 2034
rect 5570 1966 5582 2000
rect 5616 1966 5628 2000
rect 5570 1932 5628 1966
rect 5570 1898 5582 1932
rect 5616 1898 5628 1932
rect 5570 1882 5628 1898
rect 5728 2068 5786 2082
rect 5728 2034 5740 2068
rect 5774 2034 5786 2068
rect 5728 2000 5786 2034
rect 5728 1966 5740 2000
rect 5774 1966 5786 2000
rect 5728 1932 5786 1966
rect 5728 1898 5740 1932
rect 5774 1898 5786 1932
rect 5728 1882 5786 1898
rect 5878 2068 5936 2082
rect 5878 2034 5890 2068
rect 5924 2034 5936 2068
rect 5878 2000 5936 2034
rect 5878 1966 5890 2000
rect 5924 1966 5936 2000
rect 5878 1932 5936 1966
rect 5878 1898 5890 1932
rect 5924 1898 5936 1932
rect 5878 1882 5936 1898
rect 6036 2068 6094 2082
rect 6036 2034 6048 2068
rect 6082 2034 6094 2068
rect 6036 2000 6094 2034
rect 6036 1966 6048 2000
rect 6082 1966 6094 2000
rect 6036 1932 6094 1966
rect 6036 1898 6048 1932
rect 6082 1898 6094 1932
rect 6036 1882 6094 1898
rect 6230 2068 6288 2082
rect 6230 2034 6242 2068
rect 6276 2034 6288 2068
rect 6230 2000 6288 2034
rect 6230 1966 6242 2000
rect 6276 1966 6288 2000
rect 6230 1932 6288 1966
rect 6230 1898 6242 1932
rect 6276 1898 6288 1932
rect 6230 1882 6288 1898
rect 6388 2068 6446 2082
rect 6388 2034 6400 2068
rect 6434 2034 6446 2068
rect 6388 2000 6446 2034
rect 6388 1966 6400 2000
rect 6434 1966 6446 2000
rect 6388 1932 6446 1966
rect 6388 1898 6400 1932
rect 6434 1898 6446 1932
rect 6388 1882 6446 1898
rect 6538 2068 6596 2082
rect 6538 2034 6550 2068
rect 6584 2034 6596 2068
rect 6538 2000 6596 2034
rect 6538 1966 6550 2000
rect 6584 1966 6596 2000
rect 6538 1932 6596 1966
rect 6538 1898 6550 1932
rect 6584 1898 6596 1932
rect 6538 1882 6596 1898
rect 6696 2068 6754 2082
rect 6696 2034 6708 2068
rect 6742 2034 6754 2068
rect 6696 2000 6754 2034
rect 6696 1966 6708 2000
rect 6742 1966 6754 2000
rect 6696 1932 6754 1966
rect 6696 1898 6708 1932
rect 6742 1898 6754 1932
rect 6696 1882 6754 1898
rect 1280 829 1338 844
rect 1280 795 1292 829
rect 1326 795 1338 829
rect 1280 761 1338 795
rect 1280 727 1292 761
rect 1326 727 1338 761
rect 1280 693 1338 727
rect 1280 659 1292 693
rect 1326 659 1338 693
rect 1280 644 1338 659
rect 1438 829 1496 844
rect 1438 795 1450 829
rect 1484 795 1496 829
rect 1438 761 1496 795
rect 1438 727 1450 761
rect 1484 727 1496 761
rect 1438 693 1496 727
rect 1438 659 1450 693
rect 1484 659 1496 693
rect 1438 644 1496 659
rect 1568 829 1626 844
rect 1568 795 1580 829
rect 1614 795 1626 829
rect 1568 761 1626 795
rect 1568 727 1580 761
rect 1614 727 1626 761
rect 1568 693 1626 727
rect 1568 659 1580 693
rect 1614 659 1626 693
rect 1568 644 1626 659
rect 1726 829 1784 844
rect 1726 795 1738 829
rect 1772 795 1784 829
rect 1726 761 1784 795
rect 1726 727 1738 761
rect 1772 727 1784 761
rect 1726 693 1784 727
rect 1726 659 1738 693
rect 1772 659 1784 693
rect 1726 644 1784 659
rect 1900 829 1958 844
rect 1900 795 1912 829
rect 1946 795 1958 829
rect 1900 761 1958 795
rect 1900 727 1912 761
rect 1946 727 1958 761
rect 1900 693 1958 727
rect 1900 659 1912 693
rect 1946 659 1958 693
rect 1900 644 1958 659
rect 2058 829 2116 844
rect 2058 795 2070 829
rect 2104 795 2116 829
rect 2058 761 2116 795
rect 2058 727 2070 761
rect 2104 727 2116 761
rect 2058 693 2116 727
rect 2058 659 2070 693
rect 2104 659 2116 693
rect 2058 644 2116 659
rect 2242 829 2300 844
rect 2242 795 2254 829
rect 2288 795 2300 829
rect 2242 761 2300 795
rect 2242 727 2254 761
rect 2288 727 2300 761
rect 2242 693 2300 727
rect 2242 659 2254 693
rect 2288 659 2300 693
rect 2242 644 2300 659
rect 2400 829 2458 844
rect 2400 795 2412 829
rect 2446 795 2458 829
rect 2400 761 2458 795
rect 2400 727 2412 761
rect 2446 727 2458 761
rect 2400 693 2458 727
rect 2400 659 2412 693
rect 2446 659 2458 693
rect 2400 644 2458 659
rect 2646 829 2704 844
rect 2646 795 2658 829
rect 2692 795 2704 829
rect 2646 761 2704 795
rect 2646 727 2658 761
rect 2692 727 2704 761
rect 2646 693 2704 727
rect 2646 659 2658 693
rect 2692 659 2704 693
rect 2646 644 2704 659
rect 2804 829 2862 844
rect 2804 795 2816 829
rect 2850 795 2862 829
rect 2804 761 2862 795
rect 2804 727 2816 761
rect 2850 727 2862 761
rect 2804 693 2862 727
rect 2804 659 2816 693
rect 2850 659 2862 693
rect 2804 644 2862 659
rect 2990 829 3048 844
rect 2990 795 3002 829
rect 3036 795 3048 829
rect 2990 761 3048 795
rect 2990 727 3002 761
rect 3036 727 3048 761
rect 2990 693 3048 727
rect 2990 659 3002 693
rect 3036 659 3048 693
rect 2990 644 3048 659
rect 3148 829 3206 844
rect 3148 795 3160 829
rect 3194 795 3206 829
rect 3148 761 3206 795
rect 3148 727 3160 761
rect 3194 727 3206 761
rect 3148 693 3206 727
rect 3148 659 3160 693
rect 3194 659 3206 693
rect 3148 644 3206 659
rect 3612 839 3670 854
rect 3612 805 3624 839
rect 3658 805 3670 839
rect 3612 771 3670 805
rect 3612 737 3624 771
rect 3658 737 3670 771
rect 3612 703 3670 737
rect 3612 669 3624 703
rect 3658 669 3670 703
rect 3612 654 3670 669
rect 3770 839 3828 854
rect 3770 805 3782 839
rect 3816 805 3828 839
rect 3770 771 3828 805
rect 3770 737 3782 771
rect 3816 737 3828 771
rect 3770 703 3828 737
rect 3770 669 3782 703
rect 3816 669 3828 703
rect 3770 654 3828 669
rect 3920 839 3978 854
rect 3920 805 3932 839
rect 3966 805 3978 839
rect 3920 771 3978 805
rect 3920 737 3932 771
rect 3966 737 3978 771
rect 3920 703 3978 737
rect 3920 669 3932 703
rect 3966 669 3978 703
rect 3920 654 3978 669
rect 4078 839 4136 854
rect 4078 805 4090 839
rect 4124 805 4136 839
rect 4078 771 4136 805
rect 4078 737 4090 771
rect 4124 737 4136 771
rect 4078 703 4136 737
rect 4078 669 4090 703
rect 4124 669 4136 703
rect 4078 654 4136 669
rect 4272 839 4330 854
rect 4272 805 4284 839
rect 4318 805 4330 839
rect 4272 771 4330 805
rect 4272 737 4284 771
rect 4318 737 4330 771
rect 4272 703 4330 737
rect 4272 669 4284 703
rect 4318 669 4330 703
rect 4272 654 4330 669
rect 4430 839 4488 854
rect 4430 805 4442 839
rect 4476 805 4488 839
rect 4430 771 4488 805
rect 4430 737 4442 771
rect 4476 737 4488 771
rect 4430 703 4488 737
rect 4430 669 4442 703
rect 4476 669 4488 703
rect 4430 654 4488 669
rect 4580 839 4638 854
rect 4580 805 4592 839
rect 4626 805 4638 839
rect 4580 771 4638 805
rect 4580 737 4592 771
rect 4626 737 4638 771
rect 4580 703 4638 737
rect 4580 669 4592 703
rect 4626 669 4638 703
rect 4580 654 4638 669
rect 4738 839 4796 854
rect 4738 805 4750 839
rect 4784 805 4796 839
rect 4738 771 4796 805
rect 4738 737 4750 771
rect 4784 737 4796 771
rect 4738 703 4796 737
rect 4738 669 4750 703
rect 4784 669 4796 703
rect 4738 654 4796 669
<< mvndiffc >>
rect 451 2122 485 2156
rect 451 1554 485 1588
rect 597 2122 631 2156
rect 597 1554 631 1588
rect 741 2128 775 2162
rect 741 1560 775 1594
rect 895 2128 929 2162
rect 1292 1667 1326 1701
rect 1450 1667 1484 1701
rect 1580 1667 1614 1701
rect 1738 1667 1772 1701
rect 1912 1667 1946 1701
rect 2070 1667 2104 1701
rect 2254 1667 2288 1701
rect 2412 1667 2446 1701
rect 2658 1667 2692 1701
rect 2816 1667 2850 1701
rect 3002 1667 3036 1701
rect 3160 1667 3194 1701
rect 3624 1677 3658 1711
rect 3782 1677 3816 1711
rect 3932 1677 3966 1711
rect 4090 1677 4124 1711
rect 4284 1679 4318 1713
rect 4442 1679 4476 1713
rect 4592 1679 4626 1713
rect 4750 1679 4784 1713
rect 5582 1678 5616 1712
rect 5740 1678 5774 1712
rect 5890 1678 5924 1712
rect 6048 1678 6082 1712
rect 6242 1680 6276 1714
rect 6400 1680 6434 1714
rect 6550 1680 6584 1714
rect 6708 1680 6742 1714
rect 895 1560 929 1594
rect 451 894 485 928
rect 451 326 485 360
rect 597 894 631 928
rect 597 326 631 360
rect 741 900 775 934
rect 741 332 775 366
rect 895 900 929 934
rect 1292 439 1326 473
rect 1450 439 1484 473
rect 1580 439 1614 473
rect 1738 439 1772 473
rect 1912 439 1946 473
rect 2070 439 2104 473
rect 2254 439 2288 473
rect 2412 439 2446 473
rect 2658 439 2692 473
rect 2816 439 2850 473
rect 3002 439 3036 473
rect 3160 439 3194 473
rect 3624 449 3658 483
rect 3782 449 3816 483
rect 3932 449 3966 483
rect 4090 449 4124 483
rect 4284 451 4318 485
rect 4442 451 4476 485
rect 4592 451 4626 485
rect 4750 451 4784 485
rect 895 332 929 366
<< mvpdiffc >>
rect 1292 2023 1326 2057
rect 1292 1955 1326 1989
rect 1292 1887 1326 1921
rect 1450 2023 1484 2057
rect 1450 1955 1484 1989
rect 1450 1887 1484 1921
rect 1580 2023 1614 2057
rect 1580 1955 1614 1989
rect 1580 1887 1614 1921
rect 1738 2023 1772 2057
rect 1738 1955 1772 1989
rect 1738 1887 1772 1921
rect 1912 2023 1946 2057
rect 1912 1955 1946 1989
rect 1912 1887 1946 1921
rect 2070 2023 2104 2057
rect 2070 1955 2104 1989
rect 2070 1887 2104 1921
rect 2254 2023 2288 2057
rect 2254 1955 2288 1989
rect 2254 1887 2288 1921
rect 2412 2023 2446 2057
rect 2412 1955 2446 1989
rect 2412 1887 2446 1921
rect 2658 2023 2692 2057
rect 2658 1955 2692 1989
rect 2658 1887 2692 1921
rect 2816 2023 2850 2057
rect 2816 1955 2850 1989
rect 2816 1887 2850 1921
rect 3002 2023 3036 2057
rect 3002 1955 3036 1989
rect 3002 1887 3036 1921
rect 3160 2023 3194 2057
rect 3160 1955 3194 1989
rect 3160 1887 3194 1921
rect 3624 2033 3658 2067
rect 3624 1965 3658 1999
rect 3624 1897 3658 1931
rect 3782 2033 3816 2067
rect 3782 1965 3816 1999
rect 3782 1897 3816 1931
rect 3932 2033 3966 2067
rect 3932 1965 3966 1999
rect 3932 1897 3966 1931
rect 4090 2033 4124 2067
rect 4090 1965 4124 1999
rect 4090 1897 4124 1931
rect 4284 2033 4318 2067
rect 4284 1965 4318 1999
rect 4284 1897 4318 1931
rect 4442 2033 4476 2067
rect 4442 1965 4476 1999
rect 4442 1897 4476 1931
rect 4592 2033 4626 2067
rect 4592 1965 4626 1999
rect 4592 1897 4626 1931
rect 4750 2033 4784 2067
rect 4750 1965 4784 1999
rect 4750 1897 4784 1931
rect 5582 2034 5616 2068
rect 5582 1966 5616 2000
rect 5582 1898 5616 1932
rect 5740 2034 5774 2068
rect 5740 1966 5774 2000
rect 5740 1898 5774 1932
rect 5890 2034 5924 2068
rect 5890 1966 5924 2000
rect 5890 1898 5924 1932
rect 6048 2034 6082 2068
rect 6048 1966 6082 2000
rect 6048 1898 6082 1932
rect 6242 2034 6276 2068
rect 6242 1966 6276 2000
rect 6242 1898 6276 1932
rect 6400 2034 6434 2068
rect 6400 1966 6434 2000
rect 6400 1898 6434 1932
rect 6550 2034 6584 2068
rect 6550 1966 6584 2000
rect 6550 1898 6584 1932
rect 6708 2034 6742 2068
rect 6708 1966 6742 2000
rect 6708 1898 6742 1932
rect 1292 795 1326 829
rect 1292 727 1326 761
rect 1292 659 1326 693
rect 1450 795 1484 829
rect 1450 727 1484 761
rect 1450 659 1484 693
rect 1580 795 1614 829
rect 1580 727 1614 761
rect 1580 659 1614 693
rect 1738 795 1772 829
rect 1738 727 1772 761
rect 1738 659 1772 693
rect 1912 795 1946 829
rect 1912 727 1946 761
rect 1912 659 1946 693
rect 2070 795 2104 829
rect 2070 727 2104 761
rect 2070 659 2104 693
rect 2254 795 2288 829
rect 2254 727 2288 761
rect 2254 659 2288 693
rect 2412 795 2446 829
rect 2412 727 2446 761
rect 2412 659 2446 693
rect 2658 795 2692 829
rect 2658 727 2692 761
rect 2658 659 2692 693
rect 2816 795 2850 829
rect 2816 727 2850 761
rect 2816 659 2850 693
rect 3002 795 3036 829
rect 3002 727 3036 761
rect 3002 659 3036 693
rect 3160 795 3194 829
rect 3160 727 3194 761
rect 3160 659 3194 693
rect 3624 805 3658 839
rect 3624 737 3658 771
rect 3624 669 3658 703
rect 3782 805 3816 839
rect 3782 737 3816 771
rect 3782 669 3816 703
rect 3932 805 3966 839
rect 3932 737 3966 771
rect 3932 669 3966 703
rect 4090 805 4124 839
rect 4090 737 4124 771
rect 4090 669 4124 703
rect 4284 805 4318 839
rect 4284 737 4318 771
rect 4284 669 4318 703
rect 4442 805 4476 839
rect 4442 737 4476 771
rect 4442 669 4476 703
rect 4592 805 4626 839
rect 4592 737 4626 771
rect 4592 669 4626 703
rect 4750 805 4784 839
rect 4750 737 4784 771
rect 4750 669 4784 703
<< psubdiff >>
rect 1206 1524 1841 1576
rect 1206 1490 1235 1524
rect 1269 1490 1303 1524
rect 1337 1490 1371 1524
rect 1405 1490 1439 1524
rect 1473 1490 1507 1524
rect 1541 1490 1575 1524
rect 1609 1490 1643 1524
rect 1677 1490 1711 1524
rect 1745 1490 1779 1524
rect 1813 1490 1841 1524
rect 1206 1448 1841 1490
rect 3586 1535 4126 1588
rect 3586 1501 3635 1535
rect 3669 1501 3703 1535
rect 3737 1501 3771 1535
rect 3805 1501 3839 1535
rect 3873 1501 3907 1535
rect 3941 1501 3975 1535
rect 4009 1501 4043 1535
rect 4077 1501 4126 1535
rect 3586 1448 4126 1501
rect 5544 1536 6084 1588
rect 5544 1502 5594 1536
rect 5628 1502 5662 1536
rect 5696 1502 5730 1536
rect 5764 1502 5798 1536
rect 5832 1502 5866 1536
rect 5900 1502 5934 1536
rect 5968 1502 6002 1536
rect 6036 1502 6084 1536
rect 5544 1448 6084 1502
rect 1206 296 1841 348
rect 1206 262 1235 296
rect 1269 262 1303 296
rect 1337 262 1371 296
rect 1405 262 1439 296
rect 1473 262 1507 296
rect 1541 262 1575 296
rect 1609 262 1643 296
rect 1677 262 1711 296
rect 1745 262 1779 296
rect 1813 262 1841 296
rect 1206 220 1841 262
rect 3586 307 4126 360
rect 3586 273 3635 307
rect 3669 273 3703 307
rect 3737 273 3771 307
rect 3805 273 3839 307
rect 3873 273 3907 307
rect 3941 273 3975 307
rect 4009 273 4043 307
rect 4077 273 4126 307
rect 3586 220 4126 273
<< mvnsubdiff >>
rect 1230 2226 1762 2278
rect 1230 2192 1277 2226
rect 1311 2192 1345 2226
rect 1379 2192 1413 2226
rect 1447 2192 1481 2226
rect 1515 2192 1549 2226
rect 1583 2192 1617 2226
rect 1651 2192 1685 2226
rect 1719 2192 1762 2226
rect 1230 2138 1762 2192
rect 3616 2225 4136 2268
rect 3616 2191 3655 2225
rect 3689 2191 3723 2225
rect 3757 2191 3791 2225
rect 3825 2191 3859 2225
rect 3893 2191 3927 2225
rect 3961 2191 3995 2225
rect 4029 2191 4063 2225
rect 4097 2191 4136 2225
rect 3616 2148 4136 2191
rect 5574 2224 6094 2268
rect 5574 2190 5614 2224
rect 5648 2190 5682 2224
rect 5716 2190 5750 2224
rect 5784 2190 5818 2224
rect 5852 2190 5886 2224
rect 5920 2190 5954 2224
rect 5988 2190 6022 2224
rect 6056 2190 6094 2224
rect 5574 2148 6094 2190
rect 1230 998 1762 1050
rect 1230 964 1277 998
rect 1311 964 1345 998
rect 1379 964 1413 998
rect 1447 964 1481 998
rect 1515 964 1549 998
rect 1583 964 1617 998
rect 1651 964 1685 998
rect 1719 964 1762 998
rect 1230 910 1762 964
rect 3616 997 4136 1040
rect 3616 963 3655 997
rect 3689 963 3723 997
rect 3757 963 3791 997
rect 3825 963 3859 997
rect 3893 963 3927 997
rect 3961 963 3995 997
rect 4029 963 4063 997
rect 4097 963 4136 997
rect 3616 920 4136 963
<< psubdiffcont >>
rect 1235 1490 1269 1524
rect 1303 1490 1337 1524
rect 1371 1490 1405 1524
rect 1439 1490 1473 1524
rect 1507 1490 1541 1524
rect 1575 1490 1609 1524
rect 1643 1490 1677 1524
rect 1711 1490 1745 1524
rect 1779 1490 1813 1524
rect 3635 1501 3669 1535
rect 3703 1501 3737 1535
rect 3771 1501 3805 1535
rect 3839 1501 3873 1535
rect 3907 1501 3941 1535
rect 3975 1501 4009 1535
rect 4043 1501 4077 1535
rect 5594 1502 5628 1536
rect 5662 1502 5696 1536
rect 5730 1502 5764 1536
rect 5798 1502 5832 1536
rect 5866 1502 5900 1536
rect 5934 1502 5968 1536
rect 6002 1502 6036 1536
rect 1235 262 1269 296
rect 1303 262 1337 296
rect 1371 262 1405 296
rect 1439 262 1473 296
rect 1507 262 1541 296
rect 1575 262 1609 296
rect 1643 262 1677 296
rect 1711 262 1745 296
rect 1779 262 1813 296
rect 3635 273 3669 307
rect 3703 273 3737 307
rect 3771 273 3805 307
rect 3839 273 3873 307
rect 3907 273 3941 307
rect 3975 273 4009 307
rect 4043 273 4077 307
<< mvnsubdiffcont >>
rect 1277 2192 1311 2226
rect 1345 2192 1379 2226
rect 1413 2192 1447 2226
rect 1481 2192 1515 2226
rect 1549 2192 1583 2226
rect 1617 2192 1651 2226
rect 1685 2192 1719 2226
rect 3655 2191 3689 2225
rect 3723 2191 3757 2225
rect 3791 2191 3825 2225
rect 3859 2191 3893 2225
rect 3927 2191 3961 2225
rect 3995 2191 4029 2225
rect 4063 2191 4097 2225
rect 5614 2190 5648 2224
rect 5682 2190 5716 2224
rect 5750 2190 5784 2224
rect 5818 2190 5852 2224
rect 5886 2190 5920 2224
rect 5954 2190 5988 2224
rect 6022 2190 6056 2224
rect 1277 964 1311 998
rect 1345 964 1379 998
rect 1413 964 1447 998
rect 1481 964 1515 998
rect 1549 964 1583 998
rect 1617 964 1651 998
rect 1685 964 1719 998
rect 3655 963 3689 997
rect 3723 963 3757 997
rect 3791 963 3825 997
rect 3859 963 3893 997
rect 3927 963 3961 997
rect 3995 963 4029 997
rect 4063 963 4097 997
<< poly >>
rect 1338 2072 1438 2098
rect 1626 2072 1726 2098
rect 1958 2072 2058 2098
rect 2300 2072 2400 2098
rect 2704 2072 2804 2098
rect 3048 2072 3148 2098
rect 3670 2082 3770 2108
rect 3978 2082 4078 2108
rect 4330 2082 4430 2108
rect 4638 2082 4738 2108
rect 5628 2082 5728 2108
rect 5936 2082 6036 2108
rect 6288 2082 6388 2108
rect 6596 2082 6696 2108
rect 1338 1844 1438 1872
rect 1121 1819 1438 1844
rect 1121 1785 1151 1819
rect 1185 1785 1438 1819
rect 1121 1761 1438 1785
rect 1338 1734 1438 1761
rect 1626 1819 1726 1872
rect 1626 1785 1655 1819
rect 1689 1785 1726 1819
rect 1626 1734 1726 1785
rect 1958 1829 2058 1872
rect 2300 1850 2400 1872
rect 2503 1850 2589 1851
rect 1958 1817 2207 1829
rect 1958 1783 2155 1817
rect 2189 1783 2207 1817
rect 1958 1771 2207 1783
rect 2300 1827 2594 1850
rect 2300 1793 2529 1827
rect 2563 1793 2594 1827
rect 1958 1734 2058 1771
rect 2300 1759 2594 1793
rect 2704 1815 2804 1872
rect 2704 1781 2739 1815
rect 2773 1781 2804 1815
rect 2300 1734 2400 1759
rect 2704 1734 2804 1781
rect 2901 1825 2955 1831
rect 3048 1825 3148 1872
rect 2901 1815 3148 1825
rect 2901 1781 2911 1815
rect 2945 1781 3148 1815
rect 3536 1841 3602 1849
rect 3670 1841 3770 1882
rect 3536 1839 3770 1841
rect 3536 1805 3552 1839
rect 3586 1805 3770 1839
rect 3536 1802 3770 1805
rect 3536 1795 3602 1802
rect 2901 1771 3148 1781
rect 2901 1765 2955 1771
rect 3048 1734 3148 1771
rect 3670 1744 3770 1802
rect 3850 1832 3916 1840
rect 3978 1832 4078 1882
rect 3850 1830 4078 1832
rect 3850 1796 3866 1830
rect 3900 1796 4078 1830
rect 3850 1793 4078 1796
rect 3850 1786 3916 1793
rect 3978 1744 4078 1793
rect 4172 1824 4238 1834
rect 4330 1824 4430 1882
rect 4172 1790 4188 1824
rect 4222 1790 4430 1824
rect 4509 1842 4563 1858
rect 4509 1808 4519 1842
rect 4553 1840 4563 1842
rect 4638 1840 4738 1882
rect 4553 1809 4738 1840
rect 4553 1808 4563 1809
rect 4509 1792 4563 1808
rect 4172 1789 4430 1790
rect 4172 1780 4238 1789
rect 4330 1746 4430 1789
rect 4638 1746 4738 1809
rect 5494 1842 5560 1850
rect 5628 1842 5728 1882
rect 5494 1840 5728 1842
rect 5494 1806 5510 1840
rect 5544 1806 5728 1840
rect 5494 1802 5728 1806
rect 5494 1796 5560 1802
rect 5628 1744 5728 1802
rect 5808 1832 5874 1840
rect 5936 1832 6036 1882
rect 5808 1830 6036 1832
rect 5808 1796 5824 1830
rect 5858 1796 6036 1830
rect 5808 1794 6036 1796
rect 5808 1786 5874 1794
rect 5936 1744 6036 1794
rect 6130 1824 6196 1834
rect 6288 1824 6388 1882
rect 6130 1790 6146 1824
rect 6180 1790 6388 1824
rect 6468 1842 6522 1858
rect 6468 1808 6478 1842
rect 6512 1840 6522 1842
rect 6596 1840 6696 1882
rect 6512 1810 6696 1840
rect 6512 1808 6522 1810
rect 6468 1792 6522 1808
rect 6130 1780 6196 1790
rect 6288 1746 6388 1790
rect 6596 1746 6696 1810
rect 1338 1608 1438 1634
rect 1626 1608 1726 1634
rect 1958 1608 2058 1634
rect 2300 1608 2400 1634
rect 2704 1608 2804 1634
rect 3048 1608 3148 1634
rect 3670 1618 3770 1644
rect 3978 1618 4078 1644
rect 4330 1620 4430 1646
rect 4638 1620 4738 1646
rect 5628 1618 5728 1644
rect 5936 1618 6036 1644
rect 6288 1620 6388 1646
rect 6596 1620 6696 1646
rect 1338 844 1438 870
rect 1626 844 1726 870
rect 1958 844 2058 870
rect 2300 844 2400 870
rect 2704 844 2804 870
rect 3048 844 3148 870
rect 3670 854 3770 880
rect 3978 854 4078 880
rect 4330 854 4430 880
rect 4638 854 4738 880
rect 1338 616 1438 644
rect 1121 591 1438 616
rect 1121 557 1151 591
rect 1185 557 1438 591
rect 1121 533 1438 557
rect 1338 506 1438 533
rect 1626 591 1726 644
rect 1626 557 1655 591
rect 1689 557 1726 591
rect 1626 506 1726 557
rect 1958 601 2058 644
rect 2300 622 2400 644
rect 2503 622 2589 623
rect 1958 589 2207 601
rect 1958 555 2155 589
rect 2189 555 2207 589
rect 1958 543 2207 555
rect 2300 599 2594 622
rect 2300 565 2529 599
rect 2563 565 2594 599
rect 1958 506 2058 543
rect 2300 531 2594 565
rect 2704 587 2804 644
rect 2704 553 2739 587
rect 2773 553 2804 587
rect 2300 506 2400 531
rect 2704 506 2804 553
rect 2901 597 2955 603
rect 3048 597 3148 644
rect 2901 587 3148 597
rect 2901 553 2911 587
rect 2945 553 3148 587
rect 3536 613 3602 621
rect 3670 613 3770 654
rect 3536 611 3770 613
rect 3536 577 3552 611
rect 3586 577 3770 611
rect 3536 574 3770 577
rect 3536 567 3602 574
rect 2901 543 3148 553
rect 2901 537 2955 543
rect 3048 506 3148 543
rect 3670 516 3770 574
rect 3850 604 3916 612
rect 3978 604 4078 654
rect 3850 602 4078 604
rect 3850 568 3866 602
rect 3900 568 4078 602
rect 3850 565 4078 568
rect 3850 558 3916 565
rect 3978 516 4078 565
rect 4172 596 4238 606
rect 4330 596 4430 654
rect 4172 562 4188 596
rect 4222 562 4430 596
rect 4509 614 4563 630
rect 4509 580 4519 614
rect 4553 612 4563 614
rect 4638 612 4738 654
rect 4553 581 4738 612
rect 4553 580 4563 581
rect 4509 564 4563 580
rect 4172 561 4430 562
rect 4172 552 4238 561
rect 4330 518 4430 561
rect 4638 518 4738 581
rect 1338 380 1438 406
rect 1626 380 1726 406
rect 1958 380 2058 406
rect 2300 380 2400 406
rect 2704 380 2804 406
rect 3048 380 3148 406
rect 3670 390 3770 416
rect 3978 390 4078 416
rect 4330 392 4430 418
rect 4638 392 4738 418
<< polycont >>
rect 1151 1785 1185 1819
rect 1655 1785 1689 1819
rect 2155 1783 2189 1817
rect 2529 1793 2563 1827
rect 2739 1781 2773 1815
rect 2911 1781 2945 1815
rect 3552 1805 3586 1839
rect 3866 1796 3900 1830
rect 4188 1790 4222 1824
rect 4519 1808 4553 1842
rect 5510 1806 5544 1840
rect 5824 1796 5858 1830
rect 6146 1790 6180 1824
rect 6478 1808 6512 1842
rect 1151 557 1185 591
rect 1655 557 1689 591
rect 2155 555 2189 589
rect 2529 565 2563 599
rect 2739 553 2773 587
rect 2911 553 2945 587
rect 3552 577 3586 611
rect 3866 568 3900 602
rect 4188 562 4222 596
rect 4519 580 4553 614
<< mvndiffres >>
rect 426 1645 510 2065
rect 572 1645 656 2065
rect 716 1651 800 2071
rect 870 1651 954 2071
rect 426 417 510 837
rect 572 417 656 837
rect 716 423 800 843
rect 870 423 954 843
<< locali >>
rect 1230 2226 1762 2278
rect 1230 2192 1265 2226
rect 1311 2192 1337 2226
rect 1379 2192 1409 2226
rect 1447 2192 1481 2226
rect 1515 2192 1549 2226
rect 1587 2192 1617 2226
rect 1659 2192 1685 2226
rect 1731 2192 1762 2226
rect 3606 2225 4146 2278
rect 422 2140 451 2156
rect 485 2140 514 2156
rect 422 2122 448 2140
rect 489 2122 514 2140
rect 568 2140 597 2156
rect 631 2140 660 2156
rect 568 2122 592 2140
rect 633 2122 660 2140
rect 712 2145 741 2162
rect 775 2145 804 2162
rect 712 2128 738 2145
rect 779 2128 804 2145
rect 866 2145 895 2162
rect 929 2145 958 2162
rect 866 2128 891 2145
rect 932 2128 958 2145
rect 1230 2138 1762 2192
rect 2509 2145 2955 2199
rect 438 2100 448 2122
rect 489 2100 498 2122
rect 438 2082 498 2100
rect 584 2100 592 2122
rect 633 2100 644 2122
rect 584 2082 644 2100
rect 728 2105 738 2128
rect 779 2105 788 2128
rect 728 2088 788 2105
rect 882 2105 891 2128
rect 932 2105 942 2128
rect 882 2088 942 2105
rect 1292 2057 1326 2076
rect 1292 1989 1326 1991
rect 1292 1953 1326 1955
rect 1292 1868 1326 1887
rect 1450 2057 1484 2076
rect 1450 1989 1484 1991
rect 1450 1953 1484 1955
rect 1450 1868 1484 1887
rect 1580 2057 1614 2076
rect 1580 1989 1614 1991
rect 1580 1953 1614 1955
rect 1580 1868 1614 1887
rect 1738 2057 1772 2076
rect 1738 1989 1772 1991
rect 1738 1953 1772 1955
rect 1738 1868 1772 1887
rect 1912 2057 1946 2076
rect 1912 1989 1946 1991
rect 1912 1953 1946 1955
rect 1912 1868 1946 1887
rect 2070 2057 2104 2076
rect 2070 1989 2104 1991
rect 2070 1953 2104 1955
rect 2070 1868 2104 1887
rect 2254 2057 2288 2076
rect 2254 1989 2288 1991
rect 2254 1953 2288 1955
rect 2254 1868 2288 1887
rect 2412 2057 2446 2076
rect 2509 1995 2563 2145
rect 2658 2057 2692 2076
rect 2412 1989 2446 1991
rect 2412 1953 2446 1955
rect 2412 1868 2446 1887
rect 2507 1973 2585 1995
rect 2507 1939 2529 1973
rect 2563 1939 2585 1973
rect 1137 1838 1200 1850
rect 1133 1819 1204 1838
rect 2507 1835 2585 1939
rect 2658 1989 2692 1991
rect 2658 1953 2692 1955
rect 2658 1868 2692 1887
rect 2816 2057 2850 2076
rect 2816 1989 2850 1991
rect 2816 1953 2850 1955
rect 2816 1868 2850 1887
rect 1655 1826 1689 1835
rect 2153 1829 2191 1835
rect 1133 1785 1151 1819
rect 1185 1785 1204 1819
rect 1133 1767 1204 1785
rect 1648 1819 1696 1826
rect 1648 1785 1655 1819
rect 1689 1785 1696 1819
rect 1648 1778 1696 1785
rect 2143 1817 2201 1829
rect 2143 1783 2155 1817
rect 2189 1783 2201 1817
rect 2497 1827 2595 1835
rect 2497 1793 2529 1827
rect 2563 1793 2595 1827
rect 2739 1822 2773 1831
rect 2497 1786 2595 1793
rect 2732 1815 2780 1822
rect 2901 1815 2955 2145
rect 3606 2191 3655 2225
rect 3713 2191 3723 2225
rect 3785 2191 3791 2225
rect 3857 2191 3859 2225
rect 3893 2191 3895 2225
rect 3961 2191 3967 2225
rect 4029 2191 4039 2225
rect 4097 2191 4146 2225
rect 3606 2138 4146 2191
rect 5564 2224 6104 2278
rect 5564 2190 5614 2224
rect 5672 2190 5682 2224
rect 5744 2190 5750 2224
rect 5816 2190 5818 2224
rect 5852 2190 5854 2224
rect 5920 2190 5926 2224
rect 5988 2190 5998 2224
rect 6056 2190 6104 2224
rect 5564 2138 6104 2190
rect 3002 2057 3036 2076
rect 3002 1989 3036 1991
rect 3002 1953 3036 1955
rect 3002 1868 3036 1887
rect 3160 2057 3194 2076
rect 3160 1989 3194 1991
rect 3160 1953 3194 1955
rect 3160 1868 3194 1887
rect 3624 2067 3658 2086
rect 3624 1999 3658 2001
rect 3624 1963 3658 1965
rect 3624 1878 3658 1897
rect 3782 2067 3816 2086
rect 3782 1999 3816 2001
rect 3782 1963 3816 1965
rect 3782 1878 3816 1897
rect 3932 2067 3966 2086
rect 3932 1999 3966 2001
rect 3932 1963 3966 1965
rect 3932 1878 3966 1897
rect 4090 2067 4124 2086
rect 4090 1999 4124 2001
rect 4090 1963 4124 1965
rect 4090 1878 4124 1897
rect 4284 2067 4318 2086
rect 4284 1999 4318 2001
rect 4284 1963 4318 1965
rect 4284 1878 4318 1897
rect 4442 2067 4476 2086
rect 4442 1999 4476 2001
rect 4442 1963 4476 1965
rect 4442 1878 4476 1897
rect 4592 2067 4626 2086
rect 4592 1999 4626 2001
rect 4592 1963 4626 1965
rect 4592 1878 4626 1897
rect 4750 2067 4784 2086
rect 4750 1999 4784 2001
rect 4750 1963 4784 1965
rect 4750 1878 4784 1897
rect 5582 2068 5616 2086
rect 5582 2000 5616 2002
rect 5582 1964 5616 1966
rect 5582 1878 5616 1898
rect 5740 2068 5774 2086
rect 5740 2000 5774 2002
rect 5740 1964 5774 1966
rect 5740 1878 5774 1898
rect 5890 2068 5924 2086
rect 5890 2000 5924 2002
rect 5890 1964 5924 1966
rect 5890 1878 5924 1898
rect 6048 2068 6082 2086
rect 6048 2000 6082 2002
rect 6048 1964 6082 1966
rect 6048 1878 6082 1898
rect 6242 2068 6276 2086
rect 6242 2000 6276 2002
rect 6242 1964 6276 1966
rect 6242 1878 6276 1898
rect 6400 2068 6434 2086
rect 6400 2000 6434 2002
rect 6400 1964 6434 1966
rect 6400 1878 6434 1898
rect 6550 2068 6584 2086
rect 6550 2000 6584 2002
rect 6550 1964 6584 1966
rect 6550 1878 6584 1898
rect 6708 2068 6742 2086
rect 6708 2000 6742 2002
rect 6708 1964 6742 1966
rect 6708 1878 6742 1898
rect 3552 1842 3586 1855
rect 3550 1839 3589 1842
rect 1655 1769 1689 1778
rect 2143 1771 2201 1783
rect 2507 1772 2585 1786
rect 2732 1781 2739 1815
rect 2773 1781 2780 1815
rect 2895 1781 2911 1815
rect 2945 1781 2961 1815
rect 3550 1805 3552 1839
rect 3586 1805 3589 1839
rect 3866 1833 3900 1846
rect 5510 1842 5544 1856
rect 3550 1803 3589 1805
rect 3864 1830 3903 1833
rect 3552 1789 3586 1803
rect 3864 1796 3866 1830
rect 3900 1796 3903 1830
rect 3864 1794 3903 1796
rect 4188 1825 4222 1840
rect 4188 1824 4223 1825
rect 2732 1774 2780 1781
rect 1137 1755 1200 1767
rect 2153 1765 2191 1771
rect 1292 1701 1326 1738
rect 438 1612 498 1628
rect 438 1588 447 1612
rect 488 1588 498 1612
rect 584 1612 644 1628
rect 584 1588 594 1612
rect 635 1588 644 1612
rect 728 1617 788 1634
rect 728 1594 738 1617
rect 779 1594 788 1617
rect 882 1618 942 1634
rect 1292 1630 1326 1667
rect 1450 1701 1484 1738
rect 1450 1630 1484 1667
rect 1580 1701 1614 1738
rect 1580 1630 1614 1667
rect 1738 1701 1772 1738
rect 1738 1630 1772 1667
rect 1912 1701 1946 1738
rect 1912 1630 1946 1667
rect 2070 1701 2104 1738
rect 2070 1630 2104 1667
rect 2234 1701 2302 1744
rect 2234 1667 2254 1701
rect 2288 1667 2302 1701
rect 882 1594 892 1618
rect 933 1594 942 1618
rect 422 1572 447 1588
rect 488 1572 514 1588
rect 422 1554 451 1572
rect 485 1554 514 1572
rect 568 1572 594 1588
rect 635 1572 660 1588
rect 568 1554 597 1572
rect 631 1554 660 1572
rect 712 1577 738 1594
rect 779 1577 804 1594
rect 712 1560 741 1577
rect 775 1560 804 1577
rect 866 1578 892 1594
rect 933 1578 958 1594
rect 866 1560 895 1578
rect 929 1560 958 1578
rect 1206 1524 1842 1588
rect 1206 1490 1235 1524
rect 1289 1490 1303 1524
rect 1361 1490 1371 1524
rect 1433 1490 1439 1524
rect 1505 1490 1507 1524
rect 1541 1490 1543 1524
rect 1609 1490 1615 1524
rect 1677 1490 1687 1524
rect 1745 1490 1759 1524
rect 1813 1490 1842 1524
rect 1206 1448 1842 1490
rect 2234 1499 2302 1667
rect 2412 1701 2446 1738
rect 2412 1630 2446 1667
rect 2234 1465 2251 1499
rect 2285 1465 2302 1499
rect 2234 1448 2302 1465
rect 2524 1403 2578 1772
rect 2739 1765 2773 1774
rect 2901 1771 2955 1781
rect 3866 1780 3900 1794
rect 4222 1790 4223 1824
rect 4503 1808 4519 1842
rect 4553 1808 4569 1842
rect 5508 1840 5548 1842
rect 5508 1806 5510 1840
rect 5544 1806 5548 1840
rect 5824 1834 5858 1846
rect 5508 1804 5548 1806
rect 5822 1830 5862 1834
rect 5510 1790 5544 1804
rect 5822 1796 5824 1830
rect 5858 1796 5862 1830
rect 5822 1794 5862 1796
rect 6146 1826 6180 1840
rect 6146 1824 6182 1826
rect 4188 1774 4222 1790
rect 5824 1780 5858 1794
rect 6180 1790 6182 1824
rect 6462 1808 6478 1842
rect 6512 1808 6528 1842
rect 6146 1774 6180 1790
rect 2658 1701 2692 1738
rect 2658 1630 2692 1667
rect 2816 1701 2850 1738
rect 2816 1630 2850 1667
rect 3002 1701 3036 1738
rect 3002 1630 3036 1667
rect 3160 1701 3194 1738
rect 3160 1630 3194 1667
rect 3624 1711 3658 1748
rect 3624 1640 3658 1677
rect 3782 1711 3816 1748
rect 3782 1640 3816 1677
rect 3932 1711 3966 1748
rect 3932 1640 3966 1677
rect 4090 1711 4124 1748
rect 4090 1640 4124 1677
rect 4284 1713 4318 1750
rect 4284 1642 4318 1679
rect 4442 1713 4476 1750
rect 4442 1642 4476 1679
rect 4592 1713 4626 1750
rect 4592 1642 4626 1679
rect 4750 1713 4784 1750
rect 4750 1642 4784 1679
rect 5582 1712 5616 1748
rect 5582 1640 5616 1678
rect 5740 1712 5774 1748
rect 5740 1640 5774 1678
rect 5890 1712 5924 1748
rect 5890 1640 5924 1678
rect 6048 1712 6082 1748
rect 6048 1640 6082 1678
rect 6242 1714 6276 1750
rect 6242 1642 6276 1680
rect 6400 1714 6434 1750
rect 6400 1642 6434 1680
rect 6550 1714 6584 1750
rect 6550 1642 6584 1680
rect 6708 1714 6742 1750
rect 6708 1642 6742 1680
rect 3586 1535 4126 1588
rect 3586 1501 3623 1535
rect 3669 1501 3695 1535
rect 3737 1501 3767 1535
rect 3805 1501 3839 1535
rect 3873 1501 3907 1535
rect 3945 1501 3975 1535
rect 4017 1501 4043 1535
rect 4089 1501 4126 1535
rect 3586 1448 4126 1501
rect 5544 1536 6084 1588
rect 5544 1502 5582 1536
rect 5628 1502 5654 1536
rect 5696 1502 5726 1536
rect 5764 1502 5798 1536
rect 5832 1502 5866 1536
rect 5904 1502 5934 1536
rect 5976 1502 6002 1536
rect 6048 1502 6084 1536
rect 5544 1448 6084 1502
rect 1230 998 1762 1050
rect 1230 964 1265 998
rect 1311 964 1337 998
rect 1379 964 1409 998
rect 1447 964 1481 998
rect 1515 964 1549 998
rect 1587 964 1617 998
rect 1659 964 1685 998
rect 1731 964 1762 998
rect 3606 997 4146 1050
rect 422 912 451 928
rect 485 912 514 928
rect 422 894 448 912
rect 489 894 514 912
rect 568 912 597 928
rect 631 912 660 928
rect 568 894 592 912
rect 633 894 660 912
rect 712 917 741 934
rect 775 917 804 934
rect 712 900 738 917
rect 779 900 804 917
rect 866 917 895 934
rect 929 917 958 934
rect 866 900 891 917
rect 932 900 958 917
rect 1230 910 1762 964
rect 2509 917 2955 971
rect 438 872 448 894
rect 489 872 498 894
rect 438 854 498 872
rect 584 872 592 894
rect 633 872 644 894
rect 584 854 644 872
rect 728 877 738 900
rect 779 877 788 900
rect 728 860 788 877
rect 882 877 891 900
rect 932 877 942 900
rect 882 860 942 877
rect 1292 829 1326 848
rect 1292 761 1326 763
rect 1292 725 1326 727
rect 1292 640 1326 659
rect 1450 829 1484 848
rect 1450 761 1484 763
rect 1450 725 1484 727
rect 1450 640 1484 659
rect 1580 829 1614 848
rect 1580 761 1614 763
rect 1580 725 1614 727
rect 1580 640 1614 659
rect 1738 829 1772 848
rect 1738 761 1772 763
rect 1738 725 1772 727
rect 1738 640 1772 659
rect 1912 829 1946 848
rect 1912 761 1946 763
rect 1912 725 1946 727
rect 1912 640 1946 659
rect 2070 829 2104 848
rect 2070 761 2104 763
rect 2070 725 2104 727
rect 2070 640 2104 659
rect 2254 829 2288 848
rect 2254 761 2288 763
rect 2254 725 2288 727
rect 2254 640 2288 659
rect 2412 829 2446 848
rect 2509 767 2563 917
rect 2658 829 2692 848
rect 2412 761 2446 763
rect 2412 725 2446 727
rect 2412 640 2446 659
rect 2507 745 2585 767
rect 2507 711 2529 745
rect 2563 711 2585 745
rect 1137 610 1200 622
rect 1133 591 1204 610
rect 2507 607 2585 711
rect 2658 761 2692 763
rect 2658 725 2692 727
rect 2658 640 2692 659
rect 2816 829 2850 848
rect 2816 761 2850 763
rect 2816 725 2850 727
rect 2816 640 2850 659
rect 1655 598 1689 607
rect 2153 601 2191 607
rect 1133 557 1151 591
rect 1185 557 1204 591
rect 1133 539 1204 557
rect 1648 591 1696 598
rect 1648 557 1655 591
rect 1689 557 1696 591
rect 1648 550 1696 557
rect 2143 589 2201 601
rect 2143 555 2155 589
rect 2189 555 2201 589
rect 2497 599 2595 607
rect 2497 565 2529 599
rect 2563 565 2595 599
rect 2739 594 2773 603
rect 2497 558 2595 565
rect 2732 587 2780 594
rect 2901 587 2955 917
rect 3606 963 3655 997
rect 3713 963 3723 997
rect 3785 963 3791 997
rect 3857 963 3859 997
rect 3893 963 3895 997
rect 3961 963 3967 997
rect 4029 963 4039 997
rect 4097 963 4146 997
rect 3606 910 4146 963
rect 3002 829 3036 848
rect 3002 761 3036 763
rect 3002 725 3036 727
rect 3002 640 3036 659
rect 3160 829 3194 848
rect 3160 761 3194 763
rect 3160 725 3194 727
rect 3160 640 3194 659
rect 3624 839 3658 858
rect 3624 771 3658 773
rect 3624 735 3658 737
rect 3624 650 3658 669
rect 3782 839 3816 858
rect 3782 771 3816 773
rect 3782 735 3816 737
rect 3782 650 3816 669
rect 3932 839 3966 858
rect 3932 771 3966 773
rect 3932 735 3966 737
rect 3932 650 3966 669
rect 4090 839 4124 858
rect 4090 771 4124 773
rect 4090 735 4124 737
rect 4090 650 4124 669
rect 4284 839 4318 858
rect 4284 771 4318 773
rect 4284 735 4318 737
rect 4284 650 4318 669
rect 4442 839 4476 858
rect 4442 771 4476 773
rect 4442 735 4476 737
rect 4442 650 4476 669
rect 4592 839 4626 858
rect 4592 771 4626 773
rect 4592 735 4626 737
rect 4592 650 4626 669
rect 4750 839 4784 858
rect 4750 771 4784 773
rect 4750 735 4784 737
rect 4750 650 4784 669
rect 3552 614 3586 627
rect 3550 611 3589 614
rect 1655 541 1689 550
rect 2143 543 2201 555
rect 2507 544 2585 558
rect 2732 553 2739 587
rect 2773 553 2780 587
rect 2895 553 2911 587
rect 2945 553 2961 587
rect 3550 577 3552 611
rect 3586 577 3589 611
rect 3866 605 3900 618
rect 3550 575 3589 577
rect 3864 602 3903 605
rect 3552 561 3586 575
rect 3864 568 3866 602
rect 3900 568 3903 602
rect 3864 566 3903 568
rect 4188 597 4222 612
rect 4188 596 4223 597
rect 2732 546 2780 553
rect 1137 527 1200 539
rect 2153 537 2191 543
rect 1292 473 1326 510
rect 438 384 498 400
rect 438 360 447 384
rect 488 360 498 384
rect 584 384 644 400
rect 584 360 594 384
rect 635 360 644 384
rect 728 389 788 406
rect 728 366 738 389
rect 779 366 788 389
rect 882 390 942 406
rect 1292 402 1326 439
rect 1450 473 1484 510
rect 1450 402 1484 439
rect 1580 473 1614 510
rect 1580 402 1614 439
rect 1738 473 1772 510
rect 1738 402 1772 439
rect 1912 473 1946 510
rect 1912 402 1946 439
rect 2070 473 2104 510
rect 2070 402 2104 439
rect 2234 473 2302 516
rect 2234 439 2254 473
rect 2288 439 2302 473
rect 882 366 892 390
rect 933 366 942 390
rect 422 344 447 360
rect 488 344 514 360
rect 422 326 451 344
rect 485 326 514 344
rect 568 344 594 360
rect 635 344 660 360
rect 568 326 597 344
rect 631 326 660 344
rect 712 349 738 366
rect 779 349 804 366
rect 712 332 741 349
rect 775 332 804 349
rect 866 350 892 366
rect 933 350 958 366
rect 866 332 895 350
rect 929 332 958 350
rect 1206 296 1842 360
rect 1206 262 1235 296
rect 1289 262 1303 296
rect 1361 262 1371 296
rect 1433 262 1439 296
rect 1505 262 1507 296
rect 1541 262 1543 296
rect 1609 262 1615 296
rect 1677 262 1687 296
rect 1745 262 1759 296
rect 1813 262 1842 296
rect 1206 220 1842 262
rect 2234 271 2302 439
rect 2412 473 2446 510
rect 2412 402 2446 439
rect 2234 237 2251 271
rect 2285 237 2302 271
rect 2234 220 2302 237
rect 2524 175 2578 544
rect 2739 537 2773 546
rect 2901 543 2955 553
rect 3866 552 3900 566
rect 4222 562 4223 596
rect 4503 580 4519 614
rect 4553 580 4569 614
rect 4188 546 4222 562
rect 2658 473 2692 510
rect 2658 402 2692 439
rect 2816 473 2850 510
rect 2816 402 2850 439
rect 3002 473 3036 510
rect 3002 402 3036 439
rect 3160 473 3194 510
rect 3160 402 3194 439
rect 3624 483 3658 520
rect 3624 412 3658 449
rect 3782 483 3816 520
rect 3782 412 3816 449
rect 3932 483 3966 520
rect 3932 412 3966 449
rect 4090 483 4124 520
rect 4090 412 4124 449
rect 4284 485 4318 522
rect 4284 414 4318 451
rect 4442 485 4476 522
rect 4442 414 4476 451
rect 4592 485 4626 522
rect 4592 414 4626 451
rect 4750 485 4784 522
rect 4750 414 4784 451
rect 3586 307 4126 360
rect 3586 273 3623 307
rect 3669 273 3695 307
rect 3737 273 3767 307
rect 3805 273 3839 307
rect 3873 273 3907 307
rect 3945 273 3975 307
rect 4017 273 4043 307
rect 4089 273 4126 307
rect 3586 220 4126 273
<< viali >>
rect 1265 2192 1277 2226
rect 1277 2192 1299 2226
rect 1337 2192 1345 2226
rect 1345 2192 1371 2226
rect 1409 2192 1413 2226
rect 1413 2192 1443 2226
rect 1481 2192 1515 2226
rect 1553 2192 1583 2226
rect 1583 2192 1587 2226
rect 1625 2192 1651 2226
rect 1651 2192 1659 2226
rect 1697 2192 1719 2226
rect 1719 2192 1731 2226
rect 448 2122 451 2140
rect 451 2122 485 2140
rect 485 2122 489 2140
rect 592 2122 597 2140
rect 597 2122 631 2140
rect 631 2122 633 2140
rect 738 2128 741 2145
rect 741 2128 775 2145
rect 775 2128 779 2145
rect 891 2128 895 2145
rect 895 2128 929 2145
rect 929 2128 932 2145
rect 448 2100 489 2122
rect 592 2100 633 2122
rect 738 2105 779 2128
rect 891 2105 932 2128
rect 1292 2023 1326 2025
rect 1292 1991 1326 2023
rect 1292 1921 1326 1953
rect 1292 1919 1326 1921
rect 1450 2023 1484 2025
rect 1450 1991 1484 2023
rect 1450 1921 1484 1953
rect 1450 1919 1484 1921
rect 1580 2023 1614 2025
rect 1580 1991 1614 2023
rect 1580 1921 1614 1953
rect 1580 1919 1614 1921
rect 1738 2023 1772 2025
rect 1738 1991 1772 2023
rect 1738 1921 1772 1953
rect 1738 1919 1772 1921
rect 1912 2023 1946 2025
rect 1912 1991 1946 2023
rect 1912 1921 1946 1953
rect 1912 1919 1946 1921
rect 2070 2023 2104 2025
rect 2070 1991 2104 2023
rect 2070 1921 2104 1953
rect 2070 1919 2104 1921
rect 2254 2023 2288 2025
rect 2254 1991 2288 2023
rect 2254 1921 2288 1953
rect 2254 1919 2288 1921
rect 2412 2023 2446 2025
rect 2412 1991 2446 2023
rect 2658 2023 2692 2025
rect 2412 1921 2446 1953
rect 2412 1919 2446 1921
rect 2529 1939 2563 1973
rect 2658 1991 2692 2023
rect 2658 1921 2692 1953
rect 2658 1919 2692 1921
rect 2816 2023 2850 2025
rect 2816 1991 2850 2023
rect 2816 1921 2850 1953
rect 2816 1919 2850 1921
rect 1151 1785 1185 1819
rect 1655 1785 1689 1819
rect 2155 1783 2189 1817
rect 3679 2191 3689 2225
rect 3689 2191 3713 2225
rect 3751 2191 3757 2225
rect 3757 2191 3785 2225
rect 3823 2191 3825 2225
rect 3825 2191 3857 2225
rect 3895 2191 3927 2225
rect 3927 2191 3929 2225
rect 3967 2191 3995 2225
rect 3995 2191 4001 2225
rect 4039 2191 4063 2225
rect 4063 2191 4073 2225
rect 5638 2190 5648 2224
rect 5648 2190 5672 2224
rect 5710 2190 5716 2224
rect 5716 2190 5744 2224
rect 5782 2190 5784 2224
rect 5784 2190 5816 2224
rect 5854 2190 5886 2224
rect 5886 2190 5888 2224
rect 5926 2190 5954 2224
rect 5954 2190 5960 2224
rect 5998 2190 6022 2224
rect 6022 2190 6032 2224
rect 3002 2023 3036 2025
rect 3002 1991 3036 2023
rect 3002 1921 3036 1953
rect 3002 1919 3036 1921
rect 3160 2023 3194 2025
rect 3160 1991 3194 2023
rect 3160 1921 3194 1953
rect 3160 1919 3194 1921
rect 3624 2033 3658 2035
rect 3624 2001 3658 2033
rect 3624 1931 3658 1963
rect 3624 1929 3658 1931
rect 3782 2033 3816 2035
rect 3782 2001 3816 2033
rect 3782 1931 3816 1963
rect 3782 1929 3816 1931
rect 3932 2033 3966 2035
rect 3932 2001 3966 2033
rect 3932 1931 3966 1963
rect 3932 1929 3966 1931
rect 4090 2033 4124 2035
rect 4090 2001 4124 2033
rect 4090 1931 4124 1963
rect 4090 1929 4124 1931
rect 4284 2033 4318 2035
rect 4284 2001 4318 2033
rect 4284 1931 4318 1963
rect 4284 1929 4318 1931
rect 4442 2033 4476 2035
rect 4442 2001 4476 2033
rect 4442 1931 4476 1963
rect 4442 1929 4476 1931
rect 4592 2033 4626 2035
rect 4592 2001 4626 2033
rect 4592 1931 4626 1963
rect 4592 1929 4626 1931
rect 4750 2033 4784 2035
rect 4750 2001 4784 2033
rect 4750 1931 4784 1963
rect 4750 1929 4784 1931
rect 5582 2034 5616 2036
rect 5582 2002 5616 2034
rect 5582 1932 5616 1964
rect 5582 1930 5616 1932
rect 5740 2034 5774 2036
rect 5740 2002 5774 2034
rect 5740 1932 5774 1964
rect 5740 1930 5774 1932
rect 5890 2034 5924 2036
rect 5890 2002 5924 2034
rect 5890 1932 5924 1964
rect 5890 1930 5924 1932
rect 6048 2034 6082 2036
rect 6048 2002 6082 2034
rect 6048 1932 6082 1964
rect 6048 1930 6082 1932
rect 6242 2034 6276 2036
rect 6242 2002 6276 2034
rect 6242 1932 6276 1964
rect 6242 1930 6276 1932
rect 6400 2034 6434 2036
rect 6400 2002 6434 2034
rect 6400 1932 6434 1964
rect 6400 1930 6434 1932
rect 6550 2034 6584 2036
rect 6550 2002 6584 2034
rect 6550 1932 6584 1964
rect 6550 1930 6584 1932
rect 6708 2034 6742 2036
rect 6708 2002 6742 2034
rect 6708 1932 6742 1964
rect 6708 1930 6742 1932
rect 2739 1781 2773 1815
rect 3552 1805 3586 1839
rect 3866 1796 3900 1830
rect 1292 1667 1326 1701
rect 447 1588 488 1612
rect 594 1588 635 1612
rect 738 1594 779 1617
rect 1450 1667 1484 1701
rect 1580 1667 1614 1701
rect 1738 1667 1772 1701
rect 1912 1667 1946 1701
rect 2070 1667 2104 1701
rect 2254 1667 2288 1701
rect 892 1594 933 1618
rect 447 1572 451 1588
rect 451 1572 485 1588
rect 485 1572 488 1588
rect 594 1572 597 1588
rect 597 1572 631 1588
rect 631 1572 635 1588
rect 738 1577 741 1594
rect 741 1577 775 1594
rect 775 1577 779 1594
rect 892 1578 895 1594
rect 895 1578 929 1594
rect 929 1578 933 1594
rect 1255 1490 1269 1524
rect 1269 1490 1289 1524
rect 1327 1490 1337 1524
rect 1337 1490 1361 1524
rect 1399 1490 1405 1524
rect 1405 1490 1433 1524
rect 1471 1490 1473 1524
rect 1473 1490 1505 1524
rect 1543 1490 1575 1524
rect 1575 1490 1577 1524
rect 1615 1490 1643 1524
rect 1643 1490 1649 1524
rect 1687 1490 1711 1524
rect 1711 1490 1721 1524
rect 1759 1490 1779 1524
rect 1779 1490 1793 1524
rect 2412 1667 2446 1701
rect 2251 1465 2285 1499
rect 4188 1790 4222 1824
rect 4519 1808 4553 1842
rect 5510 1806 5544 1840
rect 5824 1796 5858 1830
rect 6146 1790 6180 1824
rect 6478 1808 6512 1842
rect 2658 1667 2692 1701
rect 2816 1667 2850 1701
rect 3002 1667 3036 1701
rect 3160 1667 3194 1701
rect 3624 1677 3658 1711
rect 3782 1677 3816 1711
rect 3932 1677 3966 1711
rect 4090 1677 4124 1711
rect 4284 1679 4318 1713
rect 4442 1679 4476 1713
rect 4592 1679 4626 1713
rect 4750 1679 4784 1713
rect 5582 1678 5616 1712
rect 5740 1678 5774 1712
rect 5890 1678 5924 1712
rect 6048 1678 6082 1712
rect 6242 1680 6276 1714
rect 6400 1680 6434 1714
rect 6550 1680 6584 1714
rect 6708 1680 6742 1714
rect 3623 1501 3635 1535
rect 3635 1501 3657 1535
rect 3695 1501 3703 1535
rect 3703 1501 3729 1535
rect 3767 1501 3771 1535
rect 3771 1501 3801 1535
rect 3839 1501 3873 1535
rect 3911 1501 3941 1535
rect 3941 1501 3945 1535
rect 3983 1501 4009 1535
rect 4009 1501 4017 1535
rect 4055 1501 4077 1535
rect 4077 1501 4089 1535
rect 5582 1502 5594 1536
rect 5594 1502 5616 1536
rect 5654 1502 5662 1536
rect 5662 1502 5688 1536
rect 5726 1502 5730 1536
rect 5730 1502 5760 1536
rect 5798 1502 5832 1536
rect 5870 1502 5900 1536
rect 5900 1502 5904 1536
rect 5942 1502 5968 1536
rect 5968 1502 5976 1536
rect 6014 1502 6036 1536
rect 6036 1502 6048 1536
rect 2524 1349 2578 1403
rect 1265 964 1277 998
rect 1277 964 1299 998
rect 1337 964 1345 998
rect 1345 964 1371 998
rect 1409 964 1413 998
rect 1413 964 1443 998
rect 1481 964 1515 998
rect 1553 964 1583 998
rect 1583 964 1587 998
rect 1625 964 1651 998
rect 1651 964 1659 998
rect 1697 964 1719 998
rect 1719 964 1731 998
rect 448 894 451 912
rect 451 894 485 912
rect 485 894 489 912
rect 592 894 597 912
rect 597 894 631 912
rect 631 894 633 912
rect 738 900 741 917
rect 741 900 775 917
rect 775 900 779 917
rect 891 900 895 917
rect 895 900 929 917
rect 929 900 932 917
rect 448 872 489 894
rect 592 872 633 894
rect 738 877 779 900
rect 891 877 932 900
rect 1292 795 1326 797
rect 1292 763 1326 795
rect 1292 693 1326 725
rect 1292 691 1326 693
rect 1450 795 1484 797
rect 1450 763 1484 795
rect 1450 693 1484 725
rect 1450 691 1484 693
rect 1580 795 1614 797
rect 1580 763 1614 795
rect 1580 693 1614 725
rect 1580 691 1614 693
rect 1738 795 1772 797
rect 1738 763 1772 795
rect 1738 693 1772 725
rect 1738 691 1772 693
rect 1912 795 1946 797
rect 1912 763 1946 795
rect 1912 693 1946 725
rect 1912 691 1946 693
rect 2070 795 2104 797
rect 2070 763 2104 795
rect 2070 693 2104 725
rect 2070 691 2104 693
rect 2254 795 2288 797
rect 2254 763 2288 795
rect 2254 693 2288 725
rect 2254 691 2288 693
rect 2412 795 2446 797
rect 2412 763 2446 795
rect 2658 795 2692 797
rect 2412 693 2446 725
rect 2412 691 2446 693
rect 2529 711 2563 745
rect 2658 763 2692 795
rect 2658 693 2692 725
rect 2658 691 2692 693
rect 2816 795 2850 797
rect 2816 763 2850 795
rect 2816 693 2850 725
rect 2816 691 2850 693
rect 1151 557 1185 591
rect 1655 557 1689 591
rect 2155 555 2189 589
rect 3679 963 3689 997
rect 3689 963 3713 997
rect 3751 963 3757 997
rect 3757 963 3785 997
rect 3823 963 3825 997
rect 3825 963 3857 997
rect 3895 963 3927 997
rect 3927 963 3929 997
rect 3967 963 3995 997
rect 3995 963 4001 997
rect 4039 963 4063 997
rect 4063 963 4073 997
rect 3002 795 3036 797
rect 3002 763 3036 795
rect 3002 693 3036 725
rect 3002 691 3036 693
rect 3160 795 3194 797
rect 3160 763 3194 795
rect 3160 693 3194 725
rect 3160 691 3194 693
rect 3624 805 3658 807
rect 3624 773 3658 805
rect 3624 703 3658 735
rect 3624 701 3658 703
rect 3782 805 3816 807
rect 3782 773 3816 805
rect 3782 703 3816 735
rect 3782 701 3816 703
rect 3932 805 3966 807
rect 3932 773 3966 805
rect 3932 703 3966 735
rect 3932 701 3966 703
rect 4090 805 4124 807
rect 4090 773 4124 805
rect 4090 703 4124 735
rect 4090 701 4124 703
rect 4284 805 4318 807
rect 4284 773 4318 805
rect 4284 703 4318 735
rect 4284 701 4318 703
rect 4442 805 4476 807
rect 4442 773 4476 805
rect 4442 703 4476 735
rect 4442 701 4476 703
rect 4592 805 4626 807
rect 4592 773 4626 805
rect 4592 703 4626 735
rect 4592 701 4626 703
rect 4750 805 4784 807
rect 4750 773 4784 805
rect 4750 703 4784 735
rect 4750 701 4784 703
rect 2739 553 2773 587
rect 3552 577 3586 611
rect 3866 568 3900 602
rect 1292 439 1326 473
rect 447 360 488 384
rect 594 360 635 384
rect 738 366 779 389
rect 1450 439 1484 473
rect 1580 439 1614 473
rect 1738 439 1772 473
rect 1912 439 1946 473
rect 2070 439 2104 473
rect 2254 439 2288 473
rect 892 366 933 390
rect 447 344 451 360
rect 451 344 485 360
rect 485 344 488 360
rect 594 344 597 360
rect 597 344 631 360
rect 631 344 635 360
rect 738 349 741 366
rect 741 349 775 366
rect 775 349 779 366
rect 892 350 895 366
rect 895 350 929 366
rect 929 350 933 366
rect 1255 262 1269 296
rect 1269 262 1289 296
rect 1327 262 1337 296
rect 1337 262 1361 296
rect 1399 262 1405 296
rect 1405 262 1433 296
rect 1471 262 1473 296
rect 1473 262 1505 296
rect 1543 262 1575 296
rect 1575 262 1577 296
rect 1615 262 1643 296
rect 1643 262 1649 296
rect 1687 262 1711 296
rect 1711 262 1721 296
rect 1759 262 1779 296
rect 1779 262 1793 296
rect 2412 439 2446 473
rect 2251 237 2285 271
rect 4188 562 4222 596
rect 4519 580 4553 614
rect 2658 439 2692 473
rect 2816 439 2850 473
rect 3002 439 3036 473
rect 3160 439 3194 473
rect 3624 449 3658 483
rect 3782 449 3816 483
rect 3932 449 3966 483
rect 4090 449 4124 483
rect 4284 451 4318 485
rect 4442 451 4476 485
rect 4592 451 4626 485
rect 4750 451 4784 485
rect 3623 273 3635 307
rect 3635 273 3657 307
rect 3695 273 3703 307
rect 3703 273 3729 307
rect 3767 273 3771 307
rect 3771 273 3801 307
rect 3839 273 3873 307
rect 3911 273 3941 307
rect 3941 273 3945 307
rect 3983 273 4009 307
rect 4009 273 4017 307
rect 4055 273 4077 307
rect 4077 273 4089 307
rect 2524 121 2578 175
<< metal1 >>
rect 4911 2416 4963 2422
rect 3354 2369 4789 2408
rect 1230 2235 1762 2278
rect 1230 2226 1280 2235
rect 1332 2226 1344 2235
rect 1230 2192 1265 2226
rect 1332 2192 1337 2226
rect 1230 2183 1280 2192
rect 1332 2183 1344 2192
rect 1396 2183 1408 2235
rect 1460 2183 1472 2235
rect 1524 2183 1536 2235
rect 1588 2183 1600 2235
rect 1652 2226 1664 2235
rect 1716 2226 1762 2235
rect 1659 2192 1664 2226
rect 1731 2192 1762 2226
rect 3354 2211 3393 2369
rect 4620 2327 4626 2334
rect 4440 2288 4626 2327
rect 1652 2183 1664 2192
rect 1716 2183 1762 2192
rect 432 2164 504 2168
rect 432 2112 442 2164
rect 494 2112 504 2164
rect 578 2162 650 2168
rect 432 2100 448 2112
rect 489 2100 504 2112
rect 564 2160 650 2162
rect 564 2108 584 2160
rect 636 2108 650 2160
rect 564 2106 592 2108
rect 432 2070 504 2100
rect 578 2100 592 2106
rect 633 2100 650 2108
rect 578 2070 650 2100
rect 722 2145 794 2174
rect 722 2105 738 2145
rect 779 2105 794 2145
rect 722 2076 794 2105
rect 876 2145 948 2174
rect 876 2105 891 2145
rect 932 2105 948 2145
rect 1230 2138 1762 2183
rect 876 2076 948 2105
rect 446 2030 490 2070
rect 738 2010 782 2076
rect 260 2002 315 2008
rect 728 1958 734 2010
rect 786 1958 792 2010
rect 260 1717 315 1947
rect 738 1918 782 1958
rect 890 1918 934 2076
rect 1289 2072 1330 2138
rect 1575 2072 1617 2138
rect 1823 2135 2569 2180
rect 1286 2025 1332 2072
rect 1286 1991 1292 2025
rect 1326 1991 1332 2025
rect 1286 1953 1332 1991
rect 1286 1919 1292 1953
rect 1326 1919 1332 1953
rect 590 1874 782 1918
rect 254 1662 260 1717
rect 315 1662 321 1717
rect 590 1640 634 1874
rect 880 1866 886 1918
rect 938 1866 944 1918
rect 1286 1872 1332 1919
rect 1444 2025 1490 2072
rect 1444 1991 1450 2025
rect 1484 1991 1490 2025
rect 1444 1953 1490 1991
rect 1444 1919 1450 1953
rect 1484 1919 1490 1953
rect 1444 1872 1490 1919
rect 1574 2025 1620 2072
rect 1574 1991 1580 2025
rect 1614 1991 1620 2025
rect 1574 1953 1620 1991
rect 1574 1919 1580 1953
rect 1614 1919 1620 1953
rect 1574 1872 1620 1919
rect 1732 2069 1778 2072
rect 1823 2069 1868 2135
rect 1732 2025 1868 2069
rect 1732 1991 1738 2025
rect 1772 2024 1868 2025
rect 1906 2025 1952 2072
rect 1772 1991 1778 2024
rect 1732 1953 1778 1991
rect 1906 1991 1912 2025
rect 1946 1991 1952 2025
rect 1906 1956 1952 1991
rect 1880 1954 1952 1956
rect 1732 1919 1738 1953
rect 1772 1919 1778 1953
rect 1732 1872 1778 1919
rect 1810 1953 1952 1954
rect 1810 1929 1912 1953
rect 1810 1912 1817 1929
rect 1811 1877 1817 1912
rect 1869 1919 1912 1929
rect 1946 1919 1952 1953
rect 1869 1912 1952 1919
rect 1869 1877 1875 1912
rect 1906 1872 1952 1912
rect 2064 2028 2110 2072
rect 2248 2028 2294 2072
rect 2064 2025 2294 2028
rect 2064 1991 2070 2025
rect 2104 1991 2254 2025
rect 2288 1991 2294 2025
rect 2064 1953 2294 1991
rect 2064 1919 2070 1953
rect 2104 1919 2254 1953
rect 2288 1919 2294 1953
rect 2064 1902 2294 1919
rect 2064 1872 2110 1902
rect 2248 1872 2294 1902
rect 2406 2025 2452 2072
rect 2406 1991 2412 2025
rect 2446 1991 2452 2025
rect 2524 2001 2569 2135
rect 3000 2172 3393 2211
rect 3606 2234 4146 2278
rect 3606 2182 3658 2234
rect 3710 2225 3722 2234
rect 3774 2225 3786 2234
rect 3838 2225 3850 2234
rect 3902 2225 3914 2234
rect 3966 2225 3978 2234
rect 4030 2225 4042 2234
rect 3713 2191 3722 2225
rect 3785 2191 3786 2225
rect 3966 2191 3967 2225
rect 4030 2191 4039 2225
rect 3710 2182 3722 2191
rect 3774 2182 3786 2191
rect 3838 2182 3850 2191
rect 3902 2182 3914 2191
rect 3966 2182 3978 2191
rect 4030 2182 4042 2191
rect 4094 2182 4146 2234
rect 2656 2128 2698 2129
rect 2640 2120 2698 2128
rect 2640 2068 2651 2120
rect 2703 2068 2709 2120
rect 3000 2072 3039 2172
rect 3606 2138 4146 2182
rect 3623 2082 3669 2138
rect 3618 2081 3669 2082
rect 2640 2025 2698 2068
rect 2406 1953 2452 1991
rect 2406 1919 2412 1953
rect 2446 1919 2452 1953
rect 2406 1912 2452 1919
rect 2495 1973 2597 2001
rect 2495 1939 2529 1973
rect 2563 1939 2597 1973
rect 2406 1872 2456 1912
rect 2495 1911 2597 1939
rect 2640 1991 2658 2025
rect 2692 1991 2698 2025
rect 2640 1953 2698 1991
rect 2640 1919 2658 1953
rect 2692 1919 2698 1953
rect 890 1812 934 1866
rect 1127 1831 1210 1850
rect 734 1768 934 1812
rect 1030 1829 1210 1831
rect 1030 1777 1037 1829
rect 1089 1819 1210 1829
rect 1089 1785 1151 1819
rect 1185 1785 1210 1819
rect 1089 1777 1210 1785
rect 1030 1776 1210 1777
rect 734 1646 778 1768
rect 1127 1755 1210 1776
rect 1450 1838 1484 1872
rect 1450 1828 1702 1838
rect 1450 1776 1640 1828
rect 1692 1776 1702 1828
rect 1450 1766 1702 1776
rect 1450 1734 1490 1766
rect 1735 1734 1774 1872
rect 2067 1734 2106 1872
rect 2137 1835 2207 1841
rect 2137 1826 2213 1835
rect 2137 1774 2152 1826
rect 2204 1774 2213 1826
rect 2137 1765 2213 1774
rect 2137 1759 2207 1765
rect 2250 1734 2289 1872
rect 2412 1838 2456 1872
rect 2640 1872 2698 1919
rect 2810 2025 2856 2072
rect 2810 1991 2816 2025
rect 2850 2012 2856 2025
rect 2996 2025 3042 2072
rect 2996 2012 3002 2025
rect 2850 1991 3002 2012
rect 3036 1991 3042 2025
rect 3154 2025 3200 2072
rect 3154 2015 3160 2025
rect 3194 2015 3200 2025
rect 3618 2035 3664 2081
rect 2810 1953 3042 1991
rect 3144 1963 3150 2015
rect 3202 1963 3208 2015
rect 3618 2001 3624 2035
rect 3658 2001 3664 2035
rect 3618 1963 3664 2001
rect 2810 1919 2816 1953
rect 2850 1919 3002 1953
rect 3036 1919 3042 1953
rect 2810 1902 3042 1919
rect 2810 1872 2856 1902
rect 2996 1872 3042 1902
rect 3154 1953 3200 1963
rect 3154 1919 3160 1953
rect 3194 1919 3200 1953
rect 3154 1872 3200 1919
rect 3618 1929 3624 1963
rect 3658 1929 3664 1963
rect 3618 1882 3664 1929
rect 3776 2035 3822 2082
rect 3776 2001 3782 2035
rect 3816 2001 3822 2035
rect 3776 1963 3822 2001
rect 3776 1929 3782 1963
rect 3816 1929 3822 1963
rect 3776 1882 3822 1929
rect 3926 2035 3972 2138
rect 4440 2082 4479 2288
rect 4620 2282 4626 2288
rect 4678 2282 4684 2334
rect 4750 2082 4789 2369
rect 4963 2375 6897 2405
rect 4911 2358 4963 2364
rect 6744 2327 6750 2334
rect 6398 2288 6750 2327
rect 5564 2234 6104 2278
rect 5564 2182 5616 2234
rect 5668 2224 5680 2234
rect 5732 2224 5744 2234
rect 5796 2224 5808 2234
rect 5860 2224 5872 2234
rect 5924 2224 5936 2234
rect 5988 2224 6000 2234
rect 5672 2190 5680 2224
rect 5924 2190 5926 2224
rect 5988 2190 5998 2224
rect 5668 2182 5680 2190
rect 5732 2182 5744 2190
rect 5796 2182 5808 2190
rect 5860 2182 5872 2190
rect 5924 2182 5936 2190
rect 5988 2182 6000 2190
rect 6052 2182 6104 2234
rect 5564 2138 6104 2182
rect 5582 2082 5628 2138
rect 3926 2001 3932 2035
rect 3966 2001 3972 2035
rect 3926 1963 3972 2001
rect 3926 1929 3932 1963
rect 3966 1929 3972 1963
rect 3926 1882 3972 1929
rect 4084 2035 4130 2082
rect 4084 2001 4090 2035
rect 4124 2001 4130 2035
rect 4278 2035 4324 2082
rect 4278 2009 4284 2035
rect 4084 1963 4130 2001
rect 4084 1929 4090 1963
rect 4124 1929 4130 1963
rect 4167 2007 4284 2009
rect 4167 1955 4174 2007
rect 4226 2001 4284 2007
rect 4318 2001 4324 2035
rect 4226 1963 4324 2001
rect 4226 1955 4284 1963
rect 4167 1954 4284 1955
rect 4084 1882 4130 1929
rect 4278 1929 4284 1954
rect 4318 1929 4324 1963
rect 4278 1882 4324 1929
rect 4436 2035 4482 2082
rect 4436 2001 4442 2035
rect 4476 2002 4482 2035
rect 4586 2035 4632 2082
rect 4586 2002 4592 2035
rect 4476 2001 4592 2002
rect 4626 2001 4632 2035
rect 4436 1963 4632 2001
rect 4436 1929 4442 1963
rect 4476 1936 4592 1963
rect 4476 1929 4482 1936
rect 4436 1882 4482 1929
rect 4586 1929 4592 1936
rect 4626 1929 4632 1963
rect 4586 1882 4632 1929
rect 4744 2035 4790 2082
rect 4744 2001 4750 2035
rect 4784 2001 4790 2035
rect 5576 2036 5622 2082
rect 4909 2006 4939 2015
rect 4744 1963 4790 2001
rect 4744 1929 4750 1963
rect 4784 1929 4790 1963
rect 4892 1954 4898 2006
rect 4950 1954 4956 2006
rect 5576 2002 5582 2036
rect 5616 2002 5622 2036
rect 5576 1964 5622 2002
rect 4744 1882 4790 1929
rect 4908 1913 4939 1954
rect 5576 1930 5582 1964
rect 5616 1930 5622 1964
rect 2640 1838 2684 1872
rect 2412 1794 2538 1838
rect 1124 1714 1130 1718
rect 1020 1670 1130 1714
rect 1020 1646 1064 1670
rect 1124 1666 1130 1670
rect 1182 1666 1188 1718
rect 1286 1701 1332 1734
rect 1286 1667 1292 1701
rect 1326 1667 1332 1701
rect 1286 1663 1332 1667
rect 260 1618 316 1624
rect 432 1618 504 1640
rect 316 1612 504 1618
rect 316 1572 447 1612
rect 488 1572 504 1612
rect 316 1562 504 1572
rect 260 1556 316 1562
rect 432 1542 504 1562
rect 578 1612 650 1640
rect 578 1572 594 1612
rect 635 1572 650 1612
rect 578 1542 650 1572
rect 722 1617 794 1646
rect 722 1577 738 1617
rect 779 1577 794 1617
rect 722 1548 794 1577
rect 876 1618 1064 1646
rect 876 1578 892 1618
rect 933 1602 1064 1618
rect 1281 1634 1332 1663
rect 1444 1701 1490 1734
rect 1444 1667 1450 1701
rect 1484 1667 1490 1701
rect 1574 1701 1620 1734
rect 1574 1672 1580 1701
rect 1444 1634 1490 1667
rect 1572 1667 1580 1672
rect 1614 1672 1620 1701
rect 1732 1701 1778 1734
rect 1906 1718 1952 1734
rect 1614 1667 1622 1672
rect 933 1578 948 1602
rect 1281 1588 1331 1634
rect 1572 1588 1622 1667
rect 1732 1667 1738 1701
rect 1772 1667 1778 1701
rect 1732 1634 1778 1667
rect 1896 1666 1902 1718
rect 1954 1666 1960 1718
rect 2064 1701 2110 1734
rect 2064 1667 2070 1701
rect 2104 1667 2110 1701
rect 1906 1634 1952 1666
rect 2064 1634 2110 1667
rect 2248 1701 2294 1734
rect 2406 1716 2452 1734
rect 2248 1667 2254 1701
rect 2288 1667 2294 1701
rect 2248 1634 2294 1667
rect 2398 1664 2404 1716
rect 2456 1664 2462 1716
rect 2406 1634 2452 1664
rect 1906 1602 1950 1634
rect 2494 1602 2538 1794
rect 876 1548 948 1578
rect 1206 1533 1842 1588
rect 1906 1558 2538 1602
rect 2576 1794 2684 1838
rect 2714 1824 2786 1834
rect 2576 1596 2620 1794
rect 2714 1772 2724 1824
rect 2776 1772 2786 1824
rect 2714 1762 2786 1772
rect 2815 1734 2854 1872
rect 3000 1734 3039 1872
rect 3154 1828 3198 1872
rect 3150 1822 3202 1828
rect 3437 1797 3443 1849
rect 3495 1842 3501 1849
rect 3544 1842 3595 1854
rect 3495 1839 3595 1842
rect 3495 1805 3552 1839
rect 3586 1805 3595 1839
rect 3495 1803 3595 1805
rect 3495 1797 3501 1803
rect 3544 1791 3595 1803
rect 3779 1833 3818 1882
rect 3858 1840 3909 1845
rect 3852 1833 3858 1840
rect 3779 1794 3858 1833
rect 3150 1764 3202 1770
rect 3779 1744 3818 1794
rect 3852 1788 3858 1794
rect 3910 1788 3916 1840
rect 4088 1826 4127 1882
rect 4182 1826 4229 1837
rect 4088 1824 4229 1826
rect 4088 1791 4188 1824
rect 3858 1782 3909 1788
rect 4088 1744 4127 1791
rect 4182 1790 4188 1791
rect 4222 1790 4229 1824
rect 4182 1778 4229 1790
rect 2648 1728 2700 1734
rect 2648 1670 2658 1676
rect 2652 1667 2658 1670
rect 2692 1670 2700 1676
rect 2810 1701 2856 1734
rect 2692 1667 2698 1670
rect 2652 1634 2698 1667
rect 2810 1667 2816 1701
rect 2850 1667 2856 1701
rect 2810 1634 2856 1667
rect 2996 1701 3042 1734
rect 2996 1667 3002 1701
rect 3036 1667 3042 1701
rect 2996 1634 3042 1667
rect 3154 1701 3200 1734
rect 3154 1667 3160 1701
rect 3194 1667 3200 1701
rect 3154 1634 3200 1667
rect 3156 1596 3200 1634
rect 2576 1552 3200 1596
rect 3618 1711 3664 1744
rect 3618 1677 3624 1711
rect 3658 1677 3664 1711
rect 3618 1644 3664 1677
rect 3776 1711 3822 1744
rect 3776 1677 3782 1711
rect 3816 1677 3822 1711
rect 3926 1711 3972 1744
rect 3926 1682 3932 1711
rect 3776 1644 3822 1677
rect 3924 1677 3932 1682
rect 3966 1677 3972 1711
rect 3924 1644 3972 1677
rect 4084 1711 4130 1744
rect 4084 1677 4090 1711
rect 4124 1677 4130 1711
rect 4084 1644 4130 1677
rect 3618 1588 3662 1644
rect 3924 1588 3971 1644
rect 1206 1481 1242 1533
rect 1294 1481 1306 1533
rect 1358 1524 1370 1533
rect 1422 1524 1434 1533
rect 1486 1524 1498 1533
rect 1550 1524 1562 1533
rect 1614 1524 1626 1533
rect 1678 1524 1690 1533
rect 1361 1490 1370 1524
rect 1433 1490 1434 1524
rect 1614 1490 1615 1524
rect 1678 1490 1687 1524
rect 1358 1481 1370 1490
rect 1422 1481 1434 1490
rect 1486 1481 1498 1490
rect 1550 1481 1562 1490
rect 1614 1481 1626 1490
rect 1678 1481 1690 1490
rect 1742 1481 1754 1533
rect 1806 1481 1842 1533
rect 3586 1544 4126 1588
rect 3586 1535 3638 1544
rect 3690 1535 3702 1544
rect 1206 1448 1842 1481
rect 2228 1503 2308 1528
rect 2228 1499 3399 1503
rect 2228 1465 2251 1499
rect 2285 1465 3399 1499
rect 2228 1461 3399 1465
rect 2228 1436 2308 1461
rect 2518 1403 2584 1415
rect 154 1349 160 1403
rect 214 1349 2524 1403
rect 2578 1349 2584 1403
rect 2518 1337 2584 1349
rect 3357 1308 3399 1461
rect 3586 1501 3623 1535
rect 3690 1501 3695 1535
rect 3586 1492 3638 1501
rect 3690 1492 3702 1501
rect 3754 1492 3766 1544
rect 3818 1492 3830 1544
rect 3882 1492 3894 1544
rect 3946 1492 3958 1544
rect 4010 1535 4022 1544
rect 4074 1535 4126 1544
rect 4017 1501 4022 1535
rect 4089 1501 4126 1535
rect 4010 1492 4022 1501
rect 4074 1492 4126 1501
rect 3586 1448 4126 1492
rect 3441 1343 3447 1395
rect 3499 1388 3505 1395
rect 4188 1388 4227 1778
rect 4440 1746 4479 1882
rect 4510 1851 4562 1857
rect 4507 1802 4510 1848
rect 4562 1802 4565 1848
rect 4757 1806 4786 1882
rect 4510 1793 4562 1799
rect 4757 1778 4862 1806
rect 4278 1713 4324 1746
rect 4278 1679 4284 1713
rect 4318 1679 4324 1713
rect 4278 1646 4324 1679
rect 4436 1726 4482 1746
rect 4586 1726 4632 1746
rect 4744 1726 4790 1746
rect 4436 1713 4632 1726
rect 4436 1679 4442 1713
rect 4476 1679 4592 1713
rect 4626 1679 4632 1713
rect 4436 1660 4632 1679
rect 4738 1674 4744 1726
rect 4796 1674 4802 1726
rect 4436 1646 4482 1660
rect 4586 1646 4632 1660
rect 4744 1646 4790 1674
rect 4284 1496 4312 1646
rect 4440 1601 4479 1646
rect 4434 1595 4486 1601
rect 4434 1537 4486 1543
rect 4834 1496 4862 1778
rect 4908 1728 4938 1913
rect 5576 1882 5622 1930
rect 5734 2036 5780 2082
rect 5734 2002 5740 2036
rect 5774 2002 5780 2036
rect 5734 1964 5780 2002
rect 5734 1930 5740 1964
rect 5774 1930 5780 1964
rect 5734 1882 5780 1930
rect 5884 2036 5930 2138
rect 6398 2082 6438 2288
rect 6744 2282 6750 2288
rect 6802 2282 6808 2334
rect 6867 2322 6897 2375
rect 6867 2293 6898 2322
rect 5884 2002 5890 2036
rect 5924 2002 5930 2036
rect 5884 1964 5930 2002
rect 5884 1930 5890 1964
rect 5924 1930 5930 1964
rect 5884 1882 5930 1930
rect 6042 2036 6088 2082
rect 6042 2002 6048 2036
rect 6082 2002 6088 2036
rect 6236 2036 6282 2082
rect 6236 2010 6242 2036
rect 6042 1964 6088 2002
rect 6042 1930 6048 1964
rect 6082 1930 6088 1964
rect 6126 2008 6242 2010
rect 6126 1956 6132 2008
rect 6184 2002 6242 2008
rect 6276 2002 6282 2036
rect 6184 1964 6282 2002
rect 6184 1956 6242 1964
rect 6126 1954 6242 1956
rect 6042 1882 6088 1930
rect 6236 1930 6242 1954
rect 6276 1930 6282 1964
rect 6236 1882 6282 1930
rect 6394 2036 6440 2082
rect 6394 2002 6400 2036
rect 6434 2002 6440 2036
rect 6544 2036 6590 2082
rect 6544 2002 6550 2036
rect 6584 2002 6590 2036
rect 6394 1964 6590 2002
rect 6394 1930 6400 1964
rect 6434 1936 6550 1964
rect 6434 1930 6440 1936
rect 6394 1882 6440 1930
rect 6544 1930 6550 1936
rect 6584 1930 6590 1964
rect 6544 1882 6590 1930
rect 6702 2036 6748 2082
rect 6702 2002 6708 2036
rect 6742 2002 6748 2036
rect 6868 2006 6898 2293
rect 6702 1964 6748 2002
rect 6702 1930 6708 1964
rect 6742 1930 6748 1964
rect 6850 1954 6856 2006
rect 6908 1954 6914 2006
rect 6702 1882 6748 1930
rect 6866 1914 6898 1954
rect 4993 1797 4999 1849
rect 5051 1842 5057 1849
rect 5502 1842 5554 1854
rect 5051 1840 5554 1842
rect 5051 1806 5510 1840
rect 5544 1806 5554 1840
rect 5051 1803 5554 1806
rect 5051 1797 5057 1803
rect 5502 1792 5554 1803
rect 5738 1834 5776 1882
rect 5816 1840 5868 1846
rect 5810 1834 5816 1840
rect 5738 1794 5816 1834
rect 5738 1744 5776 1794
rect 5810 1788 5816 1794
rect 5868 1788 5874 1840
rect 6046 1826 6086 1882
rect 6140 1826 6188 1838
rect 6046 1824 6188 1826
rect 6046 1792 6146 1824
rect 5816 1782 5868 1788
rect 6046 1744 6086 1792
rect 6140 1790 6146 1792
rect 6180 1790 6188 1824
rect 6140 1778 6188 1790
rect 4891 1676 4897 1728
rect 4949 1676 4955 1728
rect 5576 1712 5622 1744
rect 5576 1678 5582 1712
rect 5616 1678 5622 1712
rect 4284 1468 4862 1496
rect 3499 1349 4227 1388
rect 3499 1343 3505 1349
rect 4903 1308 4945 1676
rect 5576 1644 5622 1678
rect 5734 1712 5780 1744
rect 5734 1678 5740 1712
rect 5774 1678 5780 1712
rect 5884 1712 5930 1744
rect 5884 1682 5890 1712
rect 5734 1644 5780 1678
rect 5882 1678 5890 1682
rect 5924 1678 5930 1712
rect 5576 1588 5620 1644
rect 5882 1588 5930 1678
rect 6042 1712 6088 1744
rect 6042 1678 6048 1712
rect 6082 1678 6088 1712
rect 6042 1644 6088 1678
rect 5544 1544 6084 1588
rect 5544 1536 5596 1544
rect 5648 1536 5660 1544
rect 5544 1502 5582 1536
rect 5648 1502 5654 1536
rect 5544 1492 5596 1502
rect 5648 1492 5660 1502
rect 5712 1492 5724 1544
rect 5776 1492 5788 1544
rect 5840 1492 5852 1544
rect 5904 1492 5916 1544
rect 5968 1536 5980 1544
rect 6032 1536 6084 1544
rect 5976 1502 5980 1536
rect 6048 1502 6084 1536
rect 5968 1492 5980 1502
rect 6032 1492 6084 1502
rect 5544 1448 6084 1492
rect 4993 1343 4999 1395
rect 5051 1388 5057 1395
rect 6146 1388 6186 1778
rect 6398 1746 6438 1882
rect 6468 1852 6520 1858
rect 6466 1802 6468 1848
rect 6520 1802 6524 1848
rect 6716 1806 6744 1882
rect 6468 1794 6520 1800
rect 6716 1778 6818 1806
rect 6236 1714 6282 1746
rect 6236 1680 6242 1714
rect 6276 1680 6282 1714
rect 6236 1646 6282 1680
rect 6394 1726 6440 1746
rect 6544 1726 6590 1746
rect 6702 1726 6748 1746
rect 6394 1714 6590 1726
rect 6394 1680 6400 1714
rect 6434 1680 6550 1714
rect 6584 1680 6590 1714
rect 6394 1660 6590 1680
rect 6696 1674 6702 1726
rect 6754 1674 6760 1726
rect 6394 1646 6440 1660
rect 6544 1646 6590 1660
rect 6702 1646 6748 1674
rect 6242 1496 6270 1646
rect 6398 1602 6438 1646
rect 6392 1596 6444 1602
rect 6392 1538 6444 1544
rect 6790 1496 6818 1778
rect 6866 1728 6896 1914
rect 6850 1676 6856 1728
rect 6908 1676 6914 1728
rect 6242 1468 6818 1496
rect 6790 1404 6818 1468
rect 5051 1350 6186 1388
rect 6228 1376 6818 1404
rect 5051 1349 5454 1350
rect 5051 1343 5057 1349
rect 3357 1266 4945 1308
rect 4917 1225 4969 1231
rect 3354 1141 4789 1180
rect 6228 1213 6256 1376
rect 6790 1374 6818 1376
rect 4969 1185 6256 1213
rect 4917 1167 4969 1173
rect 1230 1007 1762 1050
rect 1230 998 1280 1007
rect 1332 998 1344 1007
rect 1230 964 1265 998
rect 1332 964 1337 998
rect 1230 955 1280 964
rect 1332 955 1344 964
rect 1396 955 1408 1007
rect 1460 955 1472 1007
rect 1524 955 1536 1007
rect 1588 955 1600 1007
rect 1652 998 1664 1007
rect 1716 998 1762 1007
rect 1659 964 1664 998
rect 1731 964 1762 998
rect 3354 983 3393 1141
rect 4620 1099 4626 1106
rect 4440 1060 4626 1099
rect 1652 955 1664 964
rect 1716 955 1762 964
rect 432 936 504 940
rect 432 884 442 936
rect 494 884 504 936
rect 578 934 650 940
rect 432 872 448 884
rect 489 872 504 884
rect 564 932 650 934
rect 564 880 584 932
rect 636 880 650 932
rect 564 878 592 880
rect 432 842 504 872
rect 578 872 592 878
rect 633 872 650 880
rect 578 842 650 872
rect 722 917 794 946
rect 722 877 738 917
rect 779 877 794 917
rect 722 848 794 877
rect 876 917 948 946
rect 876 877 891 917
rect 932 877 948 917
rect 1230 910 1762 955
rect 876 848 948 877
rect 446 802 490 842
rect 738 782 782 848
rect 260 774 315 780
rect 728 730 734 782
rect 786 730 792 782
rect 260 489 315 719
rect 738 690 782 730
rect 890 690 934 848
rect 1289 844 1330 910
rect 1575 844 1617 910
rect 1823 907 2569 952
rect 1286 797 1332 844
rect 1286 763 1292 797
rect 1326 763 1332 797
rect 1286 725 1332 763
rect 1286 691 1292 725
rect 1326 691 1332 725
rect 590 646 782 690
rect 254 434 260 489
rect 315 434 321 489
rect 590 412 634 646
rect 880 638 886 690
rect 938 638 944 690
rect 1286 644 1332 691
rect 1444 797 1490 844
rect 1444 763 1450 797
rect 1484 763 1490 797
rect 1444 725 1490 763
rect 1444 691 1450 725
rect 1484 691 1490 725
rect 1444 644 1490 691
rect 1574 797 1620 844
rect 1574 763 1580 797
rect 1614 763 1620 797
rect 1574 725 1620 763
rect 1574 691 1580 725
rect 1614 691 1620 725
rect 1574 644 1620 691
rect 1732 841 1778 844
rect 1823 841 1868 907
rect 1732 797 1868 841
rect 1732 763 1738 797
rect 1772 796 1868 797
rect 1906 797 1952 844
rect 1772 763 1778 796
rect 1732 725 1778 763
rect 1906 763 1912 797
rect 1946 763 1952 797
rect 1906 728 1952 763
rect 1880 726 1952 728
rect 1732 691 1738 725
rect 1772 691 1778 725
rect 1732 644 1778 691
rect 1810 725 1952 726
rect 1810 701 1912 725
rect 1810 684 1817 701
rect 1811 649 1817 684
rect 1869 691 1912 701
rect 1946 691 1952 725
rect 1869 684 1952 691
rect 1869 649 1875 684
rect 1906 644 1952 684
rect 2064 800 2110 844
rect 2248 800 2294 844
rect 2064 797 2294 800
rect 2064 763 2070 797
rect 2104 763 2254 797
rect 2288 763 2294 797
rect 2064 725 2294 763
rect 2064 691 2070 725
rect 2104 691 2254 725
rect 2288 691 2294 725
rect 2064 674 2294 691
rect 2064 644 2110 674
rect 2248 644 2294 674
rect 2406 797 2452 844
rect 2406 763 2412 797
rect 2446 763 2452 797
rect 2524 773 2569 907
rect 3000 944 3393 983
rect 3606 1006 4146 1050
rect 3606 954 3658 1006
rect 3710 997 3722 1006
rect 3774 997 3786 1006
rect 3838 997 3850 1006
rect 3902 997 3914 1006
rect 3966 997 3978 1006
rect 4030 997 4042 1006
rect 3713 963 3722 997
rect 3785 963 3786 997
rect 3966 963 3967 997
rect 4030 963 4039 997
rect 3710 954 3722 963
rect 3774 954 3786 963
rect 3838 954 3850 963
rect 3902 954 3914 963
rect 3966 954 3978 963
rect 4030 954 4042 963
rect 4094 954 4146 1006
rect 2656 900 2698 901
rect 2640 892 2698 900
rect 2640 840 2651 892
rect 2703 840 2709 892
rect 3000 844 3039 944
rect 3606 910 4146 954
rect 3623 854 3669 910
rect 3618 853 3669 854
rect 2640 797 2698 840
rect 2406 725 2452 763
rect 2406 691 2412 725
rect 2446 691 2452 725
rect 2406 684 2452 691
rect 2495 745 2597 773
rect 2495 711 2529 745
rect 2563 711 2597 745
rect 2406 644 2456 684
rect 2495 683 2597 711
rect 2640 763 2658 797
rect 2692 763 2698 797
rect 2640 725 2698 763
rect 2640 691 2658 725
rect 2692 691 2698 725
rect 890 584 934 638
rect 1127 603 1210 622
rect 734 540 934 584
rect 1030 601 1210 603
rect 1030 549 1037 601
rect 1089 591 1210 601
rect 1089 557 1151 591
rect 1185 557 1210 591
rect 1089 549 1210 557
rect 1030 548 1210 549
rect 734 418 778 540
rect 1127 527 1210 548
rect 1450 610 1484 644
rect 1450 600 1702 610
rect 1450 548 1640 600
rect 1692 548 1702 600
rect 1450 538 1702 548
rect 1450 506 1490 538
rect 1735 506 1774 644
rect 2067 506 2106 644
rect 2137 607 2207 613
rect 2137 598 2213 607
rect 2137 546 2152 598
rect 2204 546 2213 598
rect 2137 537 2213 546
rect 2137 531 2207 537
rect 2250 506 2289 644
rect 2412 610 2456 644
rect 2640 644 2698 691
rect 2810 797 2856 844
rect 2810 763 2816 797
rect 2850 784 2856 797
rect 2996 797 3042 844
rect 2996 784 3002 797
rect 2850 763 3002 784
rect 3036 763 3042 797
rect 3154 797 3200 844
rect 3154 787 3160 797
rect 3194 787 3200 797
rect 3618 807 3664 853
rect 2810 725 3042 763
rect 3144 735 3150 787
rect 3202 735 3208 787
rect 3618 773 3624 807
rect 3658 773 3664 807
rect 3618 735 3664 773
rect 2810 691 2816 725
rect 2850 691 3002 725
rect 3036 691 3042 725
rect 2810 674 3042 691
rect 2810 644 2856 674
rect 2996 644 3042 674
rect 3154 725 3200 735
rect 3154 691 3160 725
rect 3194 691 3200 725
rect 3154 644 3200 691
rect 3618 701 3624 735
rect 3658 701 3664 735
rect 3618 654 3664 701
rect 3776 807 3822 854
rect 3776 773 3782 807
rect 3816 773 3822 807
rect 3776 735 3822 773
rect 3776 701 3782 735
rect 3816 701 3822 735
rect 3776 654 3822 701
rect 3926 807 3972 910
rect 4440 854 4479 1060
rect 4620 1054 4626 1060
rect 4678 1054 4684 1106
rect 4750 854 4789 1141
rect 3926 773 3932 807
rect 3966 773 3972 807
rect 3926 735 3972 773
rect 3926 701 3932 735
rect 3966 701 3972 735
rect 3926 654 3972 701
rect 4084 807 4130 854
rect 4084 773 4090 807
rect 4124 773 4130 807
rect 4278 807 4324 854
rect 4278 781 4284 807
rect 4084 735 4130 773
rect 4084 701 4090 735
rect 4124 701 4130 735
rect 4167 779 4284 781
rect 4167 727 4174 779
rect 4226 773 4284 779
rect 4318 773 4324 807
rect 4226 735 4324 773
rect 4226 727 4284 735
rect 4167 726 4284 727
rect 4084 654 4130 701
rect 4278 701 4284 726
rect 4318 701 4324 735
rect 4278 654 4324 701
rect 4436 807 4482 854
rect 4436 773 4442 807
rect 4476 774 4482 807
rect 4586 807 4632 854
rect 4586 774 4592 807
rect 4476 773 4592 774
rect 4626 773 4632 807
rect 4436 735 4632 773
rect 4436 701 4442 735
rect 4476 708 4592 735
rect 4476 701 4482 708
rect 4436 654 4482 701
rect 4586 701 4592 708
rect 4626 701 4632 735
rect 4586 654 4632 701
rect 4744 807 4790 854
rect 4744 773 4750 807
rect 4784 773 4790 807
rect 4909 778 4939 787
rect 4744 735 4790 773
rect 4744 701 4750 735
rect 4784 701 4790 735
rect 4892 726 4898 778
rect 4950 726 4956 778
rect 4744 654 4790 701
rect 4908 685 4939 726
rect 2640 610 2684 644
rect 2412 566 2538 610
rect 1124 486 1130 490
rect 1020 442 1130 486
rect 1020 418 1064 442
rect 1124 438 1130 442
rect 1182 438 1188 490
rect 1286 473 1332 506
rect 1286 439 1292 473
rect 1326 439 1332 473
rect 1286 435 1332 439
rect 260 390 316 396
rect 432 390 504 412
rect 316 384 504 390
rect 316 344 447 384
rect 488 344 504 384
rect 316 334 504 344
rect 260 328 316 334
rect 432 314 504 334
rect 578 384 650 412
rect 578 344 594 384
rect 635 344 650 384
rect 578 314 650 344
rect 722 389 794 418
rect 722 349 738 389
rect 779 349 794 389
rect 722 320 794 349
rect 876 390 1064 418
rect 876 350 892 390
rect 933 374 1064 390
rect 1281 406 1332 435
rect 1444 473 1490 506
rect 1444 439 1450 473
rect 1484 439 1490 473
rect 1574 473 1620 506
rect 1574 444 1580 473
rect 1444 406 1490 439
rect 1572 439 1580 444
rect 1614 444 1620 473
rect 1732 473 1778 506
rect 1906 490 1952 506
rect 1614 439 1622 444
rect 933 350 948 374
rect 1281 360 1331 406
rect 1572 360 1622 439
rect 1732 439 1738 473
rect 1772 439 1778 473
rect 1732 406 1778 439
rect 1896 438 1902 490
rect 1954 438 1960 490
rect 2064 473 2110 506
rect 2064 439 2070 473
rect 2104 439 2110 473
rect 1906 406 1952 438
rect 2064 406 2110 439
rect 2248 473 2294 506
rect 2406 488 2452 506
rect 2248 439 2254 473
rect 2288 439 2294 473
rect 2248 406 2294 439
rect 2398 436 2404 488
rect 2456 436 2462 488
rect 2406 406 2452 436
rect 1906 374 1950 406
rect 2494 374 2538 566
rect 876 320 948 350
rect 1206 305 1842 360
rect 1906 330 2538 374
rect 2576 566 2684 610
rect 2714 596 2786 606
rect 2576 368 2620 566
rect 2714 544 2724 596
rect 2776 544 2786 596
rect 2714 534 2786 544
rect 2815 506 2854 644
rect 3000 506 3039 644
rect 3154 600 3198 644
rect 3150 594 3202 600
rect 3437 569 3443 621
rect 3495 614 3501 621
rect 3544 614 3595 626
rect 3495 611 3595 614
rect 3495 577 3552 611
rect 3586 577 3595 611
rect 3495 575 3595 577
rect 3495 569 3501 575
rect 3544 563 3595 575
rect 3779 605 3818 654
rect 3858 612 3909 617
rect 3852 605 3858 612
rect 3779 566 3858 605
rect 3150 536 3202 542
rect 3779 516 3818 566
rect 3852 560 3858 566
rect 3910 560 3916 612
rect 4088 598 4127 654
rect 4182 598 4229 609
rect 4088 596 4229 598
rect 4088 563 4188 596
rect 3858 554 3909 560
rect 4088 516 4127 563
rect 4182 562 4188 563
rect 4222 562 4229 596
rect 4182 550 4229 562
rect 2648 500 2700 506
rect 2648 442 2658 448
rect 2652 439 2658 442
rect 2692 442 2700 448
rect 2810 473 2856 506
rect 2692 439 2698 442
rect 2652 406 2698 439
rect 2810 439 2816 473
rect 2850 439 2856 473
rect 2810 406 2856 439
rect 2996 473 3042 506
rect 2996 439 3002 473
rect 3036 439 3042 473
rect 2996 406 3042 439
rect 3154 473 3200 506
rect 3154 439 3160 473
rect 3194 439 3200 473
rect 3154 406 3200 439
rect 3156 368 3200 406
rect 2576 324 3200 368
rect 3618 483 3664 516
rect 3618 449 3624 483
rect 3658 449 3664 483
rect 3618 416 3664 449
rect 3776 483 3822 516
rect 3776 449 3782 483
rect 3816 449 3822 483
rect 3926 483 3972 516
rect 3926 454 3932 483
rect 3776 416 3822 449
rect 3924 449 3932 454
rect 3966 449 3972 483
rect 3924 416 3972 449
rect 4084 483 4130 516
rect 4084 449 4090 483
rect 4124 449 4130 483
rect 4084 416 4130 449
rect 3618 360 3662 416
rect 3924 360 3971 416
rect 1206 253 1242 305
rect 1294 253 1306 305
rect 1358 296 1370 305
rect 1422 296 1434 305
rect 1486 296 1498 305
rect 1550 296 1562 305
rect 1614 296 1626 305
rect 1678 296 1690 305
rect 1361 262 1370 296
rect 1433 262 1434 296
rect 1614 262 1615 296
rect 1678 262 1687 296
rect 1358 253 1370 262
rect 1422 253 1434 262
rect 1486 253 1498 262
rect 1550 253 1562 262
rect 1614 253 1626 262
rect 1678 253 1690 262
rect 1742 253 1754 305
rect 1806 253 1842 305
rect 3586 316 4126 360
rect 3586 307 3638 316
rect 3690 307 3702 316
rect 1206 220 1842 253
rect 2228 275 2308 300
rect 2228 271 3399 275
rect 2228 237 2251 271
rect 2285 237 3399 271
rect 2228 233 3399 237
rect 2228 208 2308 233
rect 2518 175 2584 187
rect 154 121 160 175
rect 214 121 2524 175
rect 2578 121 2584 175
rect 2518 109 2584 121
rect 3357 80 3399 233
rect 3586 273 3623 307
rect 3690 273 3695 307
rect 3586 264 3638 273
rect 3690 264 3702 273
rect 3754 264 3766 316
rect 3818 264 3830 316
rect 3882 264 3894 316
rect 3946 264 3958 316
rect 4010 307 4022 316
rect 4074 307 4126 316
rect 4017 273 4022 307
rect 4089 273 4126 307
rect 4010 264 4022 273
rect 4074 264 4126 273
rect 3586 220 4126 264
rect 3441 115 3447 167
rect 3499 160 3505 167
rect 4188 160 4227 550
rect 4440 518 4479 654
rect 4510 623 4562 629
rect 4507 574 4510 620
rect 4562 574 4565 620
rect 4757 578 4786 654
rect 4510 565 4562 571
rect 4757 550 4862 578
rect 4278 485 4324 518
rect 4278 451 4284 485
rect 4318 451 4324 485
rect 4278 418 4324 451
rect 4436 498 4482 518
rect 4586 498 4632 518
rect 4744 498 4790 518
rect 4436 485 4632 498
rect 4436 451 4442 485
rect 4476 451 4592 485
rect 4626 451 4632 485
rect 4436 432 4632 451
rect 4738 446 4744 498
rect 4796 446 4802 498
rect 4436 418 4482 432
rect 4586 418 4632 432
rect 4744 418 4790 446
rect 4284 268 4312 418
rect 4440 373 4479 418
rect 4434 367 4486 373
rect 4434 309 4486 315
rect 4834 268 4862 550
rect 4908 500 4938 685
rect 4891 448 4897 500
rect 4949 448 4955 500
rect 4284 240 4862 268
rect 3499 121 4227 160
rect 3499 115 3505 121
rect 4903 80 4945 448
rect 3357 38 4945 80
<< via1 >>
rect 1280 2226 1332 2235
rect 1344 2226 1396 2235
rect 1280 2192 1299 2226
rect 1299 2192 1332 2226
rect 1344 2192 1371 2226
rect 1371 2192 1396 2226
rect 1280 2183 1332 2192
rect 1344 2183 1396 2192
rect 1408 2226 1460 2235
rect 1408 2192 1409 2226
rect 1409 2192 1443 2226
rect 1443 2192 1460 2226
rect 1408 2183 1460 2192
rect 1472 2226 1524 2235
rect 1472 2192 1481 2226
rect 1481 2192 1515 2226
rect 1515 2192 1524 2226
rect 1472 2183 1524 2192
rect 1536 2226 1588 2235
rect 1536 2192 1553 2226
rect 1553 2192 1587 2226
rect 1587 2192 1588 2226
rect 1536 2183 1588 2192
rect 1600 2226 1652 2235
rect 1664 2226 1716 2235
rect 1600 2192 1625 2226
rect 1625 2192 1652 2226
rect 1664 2192 1697 2226
rect 1697 2192 1716 2226
rect 1600 2183 1652 2192
rect 1664 2183 1716 2192
rect 442 2140 494 2164
rect 442 2112 448 2140
rect 448 2112 489 2140
rect 489 2112 494 2140
rect 584 2140 636 2160
rect 584 2108 592 2140
rect 592 2108 633 2140
rect 633 2108 636 2140
rect 260 1947 315 2002
rect 734 1958 786 2010
rect 260 1662 315 1717
rect 886 1866 938 1918
rect 1817 1877 1869 1929
rect 3658 2225 3710 2234
rect 3722 2225 3774 2234
rect 3786 2225 3838 2234
rect 3850 2225 3902 2234
rect 3914 2225 3966 2234
rect 3978 2225 4030 2234
rect 4042 2225 4094 2234
rect 3658 2191 3679 2225
rect 3679 2191 3710 2225
rect 3722 2191 3751 2225
rect 3751 2191 3774 2225
rect 3786 2191 3823 2225
rect 3823 2191 3838 2225
rect 3850 2191 3857 2225
rect 3857 2191 3895 2225
rect 3895 2191 3902 2225
rect 3914 2191 3929 2225
rect 3929 2191 3966 2225
rect 3978 2191 4001 2225
rect 4001 2191 4030 2225
rect 4042 2191 4073 2225
rect 4073 2191 4094 2225
rect 3658 2182 3710 2191
rect 3722 2182 3774 2191
rect 3786 2182 3838 2191
rect 3850 2182 3902 2191
rect 3914 2182 3966 2191
rect 3978 2182 4030 2191
rect 4042 2182 4094 2191
rect 2651 2068 2703 2120
rect 1037 1777 1089 1829
rect 1640 1819 1692 1828
rect 1640 1785 1655 1819
rect 1655 1785 1689 1819
rect 1689 1785 1692 1819
rect 1640 1776 1692 1785
rect 2152 1817 2204 1826
rect 2152 1783 2155 1817
rect 2155 1783 2189 1817
rect 2189 1783 2204 1817
rect 2152 1774 2204 1783
rect 3150 1991 3160 2015
rect 3160 1991 3194 2015
rect 3194 1991 3202 2015
rect 3150 1963 3202 1991
rect 4626 2282 4678 2334
rect 4911 2364 4963 2416
rect 5616 2224 5668 2234
rect 5680 2224 5732 2234
rect 5744 2224 5796 2234
rect 5808 2224 5860 2234
rect 5872 2224 5924 2234
rect 5936 2224 5988 2234
rect 6000 2224 6052 2234
rect 5616 2190 5638 2224
rect 5638 2190 5668 2224
rect 5680 2190 5710 2224
rect 5710 2190 5732 2224
rect 5744 2190 5782 2224
rect 5782 2190 5796 2224
rect 5808 2190 5816 2224
rect 5816 2190 5854 2224
rect 5854 2190 5860 2224
rect 5872 2190 5888 2224
rect 5888 2190 5924 2224
rect 5936 2190 5960 2224
rect 5960 2190 5988 2224
rect 6000 2190 6032 2224
rect 6032 2190 6052 2224
rect 5616 2182 5668 2190
rect 5680 2182 5732 2190
rect 5744 2182 5796 2190
rect 5808 2182 5860 2190
rect 5872 2182 5924 2190
rect 5936 2182 5988 2190
rect 6000 2182 6052 2190
rect 4174 1955 4226 2007
rect 4898 1954 4950 2006
rect 1130 1666 1182 1718
rect 260 1562 316 1618
rect 1902 1701 1954 1718
rect 1902 1667 1912 1701
rect 1912 1667 1946 1701
rect 1946 1667 1954 1701
rect 1902 1666 1954 1667
rect 2404 1701 2456 1716
rect 2404 1667 2412 1701
rect 2412 1667 2446 1701
rect 2446 1667 2456 1701
rect 2404 1664 2456 1667
rect 2724 1815 2776 1824
rect 2724 1781 2739 1815
rect 2739 1781 2773 1815
rect 2773 1781 2776 1815
rect 2724 1772 2776 1781
rect 3150 1770 3202 1822
rect 3443 1797 3495 1849
rect 3858 1830 3910 1840
rect 3858 1796 3866 1830
rect 3866 1796 3900 1830
rect 3900 1796 3910 1830
rect 3858 1788 3910 1796
rect 2648 1701 2700 1728
rect 2648 1676 2658 1701
rect 2658 1676 2692 1701
rect 2692 1676 2700 1701
rect 1242 1524 1294 1533
rect 1242 1490 1255 1524
rect 1255 1490 1289 1524
rect 1289 1490 1294 1524
rect 1242 1481 1294 1490
rect 1306 1524 1358 1533
rect 1370 1524 1422 1533
rect 1434 1524 1486 1533
rect 1498 1524 1550 1533
rect 1562 1524 1614 1533
rect 1626 1524 1678 1533
rect 1690 1524 1742 1533
rect 1306 1490 1327 1524
rect 1327 1490 1358 1524
rect 1370 1490 1399 1524
rect 1399 1490 1422 1524
rect 1434 1490 1471 1524
rect 1471 1490 1486 1524
rect 1498 1490 1505 1524
rect 1505 1490 1543 1524
rect 1543 1490 1550 1524
rect 1562 1490 1577 1524
rect 1577 1490 1614 1524
rect 1626 1490 1649 1524
rect 1649 1490 1678 1524
rect 1690 1490 1721 1524
rect 1721 1490 1742 1524
rect 1306 1481 1358 1490
rect 1370 1481 1422 1490
rect 1434 1481 1486 1490
rect 1498 1481 1550 1490
rect 1562 1481 1614 1490
rect 1626 1481 1678 1490
rect 1690 1481 1742 1490
rect 1754 1524 1806 1533
rect 1754 1490 1759 1524
rect 1759 1490 1793 1524
rect 1793 1490 1806 1524
rect 1754 1481 1806 1490
rect 3638 1535 3690 1544
rect 3702 1535 3754 1544
rect 160 1349 214 1403
rect 3638 1501 3657 1535
rect 3657 1501 3690 1535
rect 3702 1501 3729 1535
rect 3729 1501 3754 1535
rect 3638 1492 3690 1501
rect 3702 1492 3754 1501
rect 3766 1535 3818 1544
rect 3766 1501 3767 1535
rect 3767 1501 3801 1535
rect 3801 1501 3818 1535
rect 3766 1492 3818 1501
rect 3830 1535 3882 1544
rect 3830 1501 3839 1535
rect 3839 1501 3873 1535
rect 3873 1501 3882 1535
rect 3830 1492 3882 1501
rect 3894 1535 3946 1544
rect 3894 1501 3911 1535
rect 3911 1501 3945 1535
rect 3945 1501 3946 1535
rect 3894 1492 3946 1501
rect 3958 1535 4010 1544
rect 4022 1535 4074 1544
rect 3958 1501 3983 1535
rect 3983 1501 4010 1535
rect 4022 1501 4055 1535
rect 4055 1501 4074 1535
rect 3958 1492 4010 1501
rect 4022 1492 4074 1501
rect 3447 1343 3499 1395
rect 4510 1842 4562 1851
rect 4510 1808 4519 1842
rect 4519 1808 4553 1842
rect 4553 1808 4562 1842
rect 4510 1799 4562 1808
rect 4744 1713 4796 1726
rect 4744 1679 4750 1713
rect 4750 1679 4784 1713
rect 4784 1679 4796 1713
rect 4744 1674 4796 1679
rect 4434 1543 4486 1595
rect 6750 2282 6802 2334
rect 6132 1956 6184 2008
rect 6856 1954 6908 2006
rect 4999 1797 5051 1849
rect 5816 1830 5868 1840
rect 5816 1796 5824 1830
rect 5824 1796 5858 1830
rect 5858 1796 5868 1830
rect 5816 1788 5868 1796
rect 4897 1676 4949 1728
rect 5596 1536 5648 1544
rect 5660 1536 5712 1544
rect 5596 1502 5616 1536
rect 5616 1502 5648 1536
rect 5660 1502 5688 1536
rect 5688 1502 5712 1536
rect 5596 1492 5648 1502
rect 5660 1492 5712 1502
rect 5724 1536 5776 1544
rect 5724 1502 5726 1536
rect 5726 1502 5760 1536
rect 5760 1502 5776 1536
rect 5724 1492 5776 1502
rect 5788 1536 5840 1544
rect 5788 1502 5798 1536
rect 5798 1502 5832 1536
rect 5832 1502 5840 1536
rect 5788 1492 5840 1502
rect 5852 1536 5904 1544
rect 5852 1502 5870 1536
rect 5870 1502 5904 1536
rect 5852 1492 5904 1502
rect 5916 1536 5968 1544
rect 5980 1536 6032 1544
rect 5916 1502 5942 1536
rect 5942 1502 5968 1536
rect 5980 1502 6014 1536
rect 6014 1502 6032 1536
rect 5916 1492 5968 1502
rect 5980 1492 6032 1502
rect 4999 1343 5051 1395
rect 6468 1842 6520 1852
rect 6468 1808 6478 1842
rect 6478 1808 6512 1842
rect 6512 1808 6520 1842
rect 6468 1800 6520 1808
rect 6702 1714 6754 1726
rect 6702 1680 6708 1714
rect 6708 1680 6742 1714
rect 6742 1680 6754 1714
rect 6702 1674 6754 1680
rect 6392 1544 6444 1596
rect 6856 1676 6908 1728
rect 4917 1173 4969 1225
rect 1280 998 1332 1007
rect 1344 998 1396 1007
rect 1280 964 1299 998
rect 1299 964 1332 998
rect 1344 964 1371 998
rect 1371 964 1396 998
rect 1280 955 1332 964
rect 1344 955 1396 964
rect 1408 998 1460 1007
rect 1408 964 1409 998
rect 1409 964 1443 998
rect 1443 964 1460 998
rect 1408 955 1460 964
rect 1472 998 1524 1007
rect 1472 964 1481 998
rect 1481 964 1515 998
rect 1515 964 1524 998
rect 1472 955 1524 964
rect 1536 998 1588 1007
rect 1536 964 1553 998
rect 1553 964 1587 998
rect 1587 964 1588 998
rect 1536 955 1588 964
rect 1600 998 1652 1007
rect 1664 998 1716 1007
rect 1600 964 1625 998
rect 1625 964 1652 998
rect 1664 964 1697 998
rect 1697 964 1716 998
rect 1600 955 1652 964
rect 1664 955 1716 964
rect 442 912 494 936
rect 442 884 448 912
rect 448 884 489 912
rect 489 884 494 912
rect 584 912 636 932
rect 584 880 592 912
rect 592 880 633 912
rect 633 880 636 912
rect 260 719 315 774
rect 734 730 786 782
rect 260 434 315 489
rect 886 638 938 690
rect 1817 649 1869 701
rect 3658 997 3710 1006
rect 3722 997 3774 1006
rect 3786 997 3838 1006
rect 3850 997 3902 1006
rect 3914 997 3966 1006
rect 3978 997 4030 1006
rect 4042 997 4094 1006
rect 3658 963 3679 997
rect 3679 963 3710 997
rect 3722 963 3751 997
rect 3751 963 3774 997
rect 3786 963 3823 997
rect 3823 963 3838 997
rect 3850 963 3857 997
rect 3857 963 3895 997
rect 3895 963 3902 997
rect 3914 963 3929 997
rect 3929 963 3966 997
rect 3978 963 4001 997
rect 4001 963 4030 997
rect 4042 963 4073 997
rect 4073 963 4094 997
rect 3658 954 3710 963
rect 3722 954 3774 963
rect 3786 954 3838 963
rect 3850 954 3902 963
rect 3914 954 3966 963
rect 3978 954 4030 963
rect 4042 954 4094 963
rect 2651 840 2703 892
rect 1037 549 1089 601
rect 1640 591 1692 600
rect 1640 557 1655 591
rect 1655 557 1689 591
rect 1689 557 1692 591
rect 1640 548 1692 557
rect 2152 589 2204 598
rect 2152 555 2155 589
rect 2155 555 2189 589
rect 2189 555 2204 589
rect 2152 546 2204 555
rect 3150 763 3160 787
rect 3160 763 3194 787
rect 3194 763 3202 787
rect 3150 735 3202 763
rect 4626 1054 4678 1106
rect 4174 727 4226 779
rect 4898 726 4950 778
rect 1130 438 1182 490
rect 260 334 316 390
rect 1902 473 1954 490
rect 1902 439 1912 473
rect 1912 439 1946 473
rect 1946 439 1954 473
rect 1902 438 1954 439
rect 2404 473 2456 488
rect 2404 439 2412 473
rect 2412 439 2446 473
rect 2446 439 2456 473
rect 2404 436 2456 439
rect 2724 587 2776 596
rect 2724 553 2739 587
rect 2739 553 2773 587
rect 2773 553 2776 587
rect 2724 544 2776 553
rect 3150 542 3202 594
rect 3443 569 3495 621
rect 3858 602 3910 612
rect 3858 568 3866 602
rect 3866 568 3900 602
rect 3900 568 3910 602
rect 3858 560 3910 568
rect 2648 473 2700 500
rect 2648 448 2658 473
rect 2658 448 2692 473
rect 2692 448 2700 473
rect 1242 296 1294 305
rect 1242 262 1255 296
rect 1255 262 1289 296
rect 1289 262 1294 296
rect 1242 253 1294 262
rect 1306 296 1358 305
rect 1370 296 1422 305
rect 1434 296 1486 305
rect 1498 296 1550 305
rect 1562 296 1614 305
rect 1626 296 1678 305
rect 1690 296 1742 305
rect 1306 262 1327 296
rect 1327 262 1358 296
rect 1370 262 1399 296
rect 1399 262 1422 296
rect 1434 262 1471 296
rect 1471 262 1486 296
rect 1498 262 1505 296
rect 1505 262 1543 296
rect 1543 262 1550 296
rect 1562 262 1577 296
rect 1577 262 1614 296
rect 1626 262 1649 296
rect 1649 262 1678 296
rect 1690 262 1721 296
rect 1721 262 1742 296
rect 1306 253 1358 262
rect 1370 253 1422 262
rect 1434 253 1486 262
rect 1498 253 1550 262
rect 1562 253 1614 262
rect 1626 253 1678 262
rect 1690 253 1742 262
rect 1754 296 1806 305
rect 1754 262 1759 296
rect 1759 262 1793 296
rect 1793 262 1806 296
rect 1754 253 1806 262
rect 3638 307 3690 316
rect 3702 307 3754 316
rect 160 121 214 175
rect 3638 273 3657 307
rect 3657 273 3690 307
rect 3702 273 3729 307
rect 3729 273 3754 307
rect 3638 264 3690 273
rect 3702 264 3754 273
rect 3766 307 3818 316
rect 3766 273 3767 307
rect 3767 273 3801 307
rect 3801 273 3818 307
rect 3766 264 3818 273
rect 3830 307 3882 316
rect 3830 273 3839 307
rect 3839 273 3873 307
rect 3873 273 3882 307
rect 3830 264 3882 273
rect 3894 307 3946 316
rect 3894 273 3911 307
rect 3911 273 3945 307
rect 3945 273 3946 307
rect 3894 264 3946 273
rect 3958 307 4010 316
rect 4022 307 4074 316
rect 3958 273 3983 307
rect 3983 273 4010 307
rect 4022 273 4055 307
rect 4055 273 4074 307
rect 3958 264 4010 273
rect 4022 264 4074 273
rect 3447 115 3499 167
rect 4510 614 4562 623
rect 4510 580 4519 614
rect 4519 580 4553 614
rect 4553 580 4562 614
rect 4510 571 4562 580
rect 4744 485 4796 498
rect 4744 451 4750 485
rect 4750 451 4784 485
rect 4784 451 4796 485
rect 4744 446 4796 451
rect 4434 315 4486 367
rect 4897 448 4949 500
<< metal2 >>
rect -76 2234 -8 2243
rect -76 1028 -8 2166
rect 156 1831 211 2456
rect 260 2002 315 2456
rect 1230 2237 1762 2278
rect 1230 2181 1270 2237
rect 1326 2235 1350 2237
rect 1406 2235 1430 2237
rect 1486 2235 1510 2237
rect 1566 2235 1590 2237
rect 1646 2235 1670 2237
rect 1332 2183 1344 2235
rect 1406 2183 1408 2235
rect 1588 2183 1590 2235
rect 1652 2183 1664 2235
rect 1326 2181 1350 2183
rect 1406 2181 1430 2183
rect 1486 2181 1510 2183
rect 1566 2181 1590 2183
rect 1646 2181 1670 2183
rect 1726 2181 1762 2237
rect 442 2164 494 2170
rect 582 2162 638 2168
rect 494 2160 858 2162
rect 494 2112 584 2160
rect 442 2108 584 2112
rect 636 2108 858 2160
rect 1230 2138 1762 2181
rect 2641 2120 2709 2128
rect 442 2106 1150 2108
rect 582 2100 638 2106
rect 802 2100 1150 2106
rect 2641 2100 2651 2120
rect 802 2068 2651 2100
rect 2703 2068 2709 2120
rect 802 2056 2709 2068
rect 802 2052 1150 2056
rect 734 2010 786 2016
rect 254 1947 260 2002
rect 315 1947 321 2002
rect 1278 2011 2733 2020
rect 3150 2015 3202 2021
rect 1278 2006 3150 2011
rect 786 1976 3150 2006
rect 786 1962 1322 1976
rect 2733 1967 3150 1976
rect 734 1952 786 1958
rect 3150 1957 3202 1963
rect 1812 1930 1872 1941
rect 886 1918 938 1924
rect 1812 1919 1814 1930
rect 938 1907 1124 1914
rect 1481 1907 1814 1919
rect 938 1885 1814 1907
rect 938 1873 1515 1885
rect 1812 1874 1814 1885
rect 1870 1919 1872 1930
rect 1870 1885 1873 1919
rect 1870 1874 1872 1885
rect 938 1870 1124 1873
rect 886 1860 938 1866
rect 1812 1863 1872 1874
rect 3446 1855 3487 2456
rect 4905 2364 4911 2416
rect 4963 2364 4969 2416
rect 5004 2368 5045 2456
rect 5164 2368 5205 2456
rect 5244 2368 5285 2456
rect 5324 2368 5365 2456
rect 5404 2368 5445 2456
rect 4626 2334 4678 2340
rect 4918 2328 4957 2364
rect 4678 2289 4957 2328
rect 3606 2236 4146 2278
rect 4626 2276 4678 2282
rect 3606 2180 3648 2236
rect 3704 2234 3728 2236
rect 3784 2234 3808 2236
rect 3864 2234 3888 2236
rect 3944 2234 3968 2236
rect 4024 2234 4048 2236
rect 3710 2182 3722 2234
rect 3784 2182 3786 2234
rect 3966 2182 3968 2234
rect 4030 2182 4042 2234
rect 3704 2180 3728 2182
rect 3784 2180 3808 2182
rect 3864 2180 3888 2182
rect 3944 2180 3968 2182
rect 4024 2180 4048 2182
rect 4104 2180 4146 2236
rect 3606 2138 4146 2180
rect 4173 2009 4228 2015
rect 4898 2009 4950 2012
rect 4173 2007 4966 2009
rect 4173 1955 4174 2007
rect 4226 2006 4966 2007
rect 4226 1955 4898 2006
rect 4173 1954 4898 1955
rect 4950 1954 4966 2006
rect 4173 1948 4228 1954
rect 4898 1948 4950 1954
rect 5004 1855 5046 2368
rect 3443 1849 3495 1855
rect 1036 1831 1091 1837
rect 156 1829 1091 1831
rect 156 1777 1037 1829
rect 1089 1777 1091 1829
rect 156 1776 1091 1777
rect 1036 1770 1091 1776
rect 1636 1832 1696 1838
rect 2149 1832 2207 1841
rect 1636 1829 2207 1832
rect 2720 1829 2780 1834
rect 1636 1828 2780 1829
rect 1636 1776 1640 1828
rect 1692 1826 2790 1828
rect 1692 1776 2152 1826
rect 1636 1774 2152 1776
rect 2204 1824 2790 1826
rect 2204 1774 2724 1824
rect 1636 1772 2724 1774
rect 2776 1772 2790 1824
rect 1636 1766 1696 1772
rect 2149 1771 2790 1772
rect 2149 1759 2207 1771
rect 2720 1768 2790 1771
rect 3144 1770 3150 1822
rect 3202 1770 3208 1822
rect 3858 1840 3910 1846
rect 3443 1791 3495 1797
rect 3857 1791 3858 1834
rect 2720 1762 2780 1768
rect 2650 1728 2698 1732
rect 260 1717 315 1723
rect 1130 1718 1182 1724
rect 315 1714 501 1717
rect 315 1670 1130 1714
rect 315 1662 501 1670
rect 1902 1718 1954 1724
rect 2404 1720 2456 1722
rect 1182 1670 1902 1714
rect 260 1656 315 1662
rect 1130 1660 1182 1666
rect 1902 1660 1954 1666
rect 2391 1718 2469 1720
rect 2391 1662 2402 1718
rect 2458 1662 2469 1718
rect 2642 1676 2648 1728
rect 2700 1724 2706 1728
rect 3152 1724 3196 1770
rect 3446 1752 3487 1791
rect 4504 1799 4510 1851
rect 4562 1799 4568 1851
rect 4999 1849 5051 1855
rect 3858 1782 3910 1788
rect 2700 1680 3196 1724
rect 3861 1735 3900 1782
rect 4519 1735 4553 1799
rect 4999 1791 5051 1797
rect 5004 1752 5046 1791
rect 5084 1752 5126 2368
rect 5164 1752 5206 2368
rect 5244 1752 5286 2368
rect 5324 1752 5366 2368
rect 5404 1752 5446 2368
rect 6750 2334 6802 2340
rect 6802 2289 7029 2328
rect 5564 2236 6104 2278
rect 6750 2276 6802 2282
rect 5564 2180 5606 2236
rect 5662 2234 5686 2236
rect 5742 2234 5766 2236
rect 5822 2234 5846 2236
rect 5902 2234 5926 2236
rect 5982 2234 6006 2236
rect 5668 2182 5680 2234
rect 5742 2182 5744 2234
rect 5924 2182 5926 2234
rect 5988 2182 6000 2234
rect 5662 2180 5686 2182
rect 5742 2180 5766 2182
rect 5822 2180 5846 2182
rect 5902 2180 5926 2182
rect 5982 2180 6006 2182
rect 6062 2180 6104 2236
rect 5564 2138 6104 2180
rect 6132 2010 6186 2016
rect 6856 2010 6908 2012
rect 6132 2008 6924 2010
rect 6184 2006 6924 2008
rect 6184 1956 6856 2006
rect 6132 1954 6856 1956
rect 6908 1954 6924 2006
rect 6132 1948 6186 1954
rect 6856 1948 6908 1954
rect 5816 1840 5868 1846
rect 6462 1800 6468 1852
rect 6520 1800 6526 1852
rect 5816 1782 5868 1788
rect 3861 1696 4555 1735
rect 4744 1726 4796 1732
rect 2700 1676 2706 1680
rect 2391 1660 2469 1662
rect 2404 1658 2456 1660
rect 2650 1636 2694 1676
rect 4897 1728 4949 1734
rect 4796 1686 4897 1715
rect -76 951 -8 960
rect 26 1558 94 1567
rect 26 322 94 1490
rect 156 1409 211 1598
rect 254 1562 260 1618
rect 316 1562 322 1618
rect 156 1403 214 1409
rect 156 1349 160 1403
rect 159 1228 214 1349
rect 260 1390 316 1562
rect 1206 1535 1842 1588
rect 1206 1533 1256 1535
rect 1312 1533 1336 1535
rect 1392 1533 1416 1535
rect 1472 1533 1496 1535
rect 1552 1533 1576 1535
rect 1632 1533 1656 1535
rect 1712 1533 1736 1535
rect 1792 1533 1842 1535
rect 1206 1481 1242 1533
rect 1486 1481 1496 1533
rect 1552 1481 1562 1533
rect 1806 1481 1842 1533
rect 1206 1479 1256 1481
rect 1312 1479 1336 1481
rect 1392 1479 1416 1481
rect 1472 1479 1496 1481
rect 1552 1479 1576 1481
rect 1632 1479 1656 1481
rect 1712 1479 1736 1481
rect 1792 1479 1842 1481
rect 1206 1448 1842 1479
rect 3446 1401 3487 1672
rect 4744 1668 4796 1674
rect 4897 1670 4949 1676
rect 5084 1672 5125 1752
rect 5164 1672 5205 1752
rect 5244 1672 5285 1752
rect 5324 1672 5365 1752
rect 5404 1672 5445 1752
rect 5820 1736 5858 1782
rect 6478 1736 6512 1800
rect 5820 1696 6514 1736
rect 6702 1726 6754 1732
rect 6856 1728 6908 1734
rect 6754 1686 6856 1716
rect 3586 1546 4126 1588
rect 3586 1490 3628 1546
rect 3684 1544 3708 1546
rect 3764 1544 3788 1546
rect 3844 1544 3868 1546
rect 3924 1544 3948 1546
rect 4004 1544 4028 1546
rect 3690 1492 3702 1544
rect 3764 1492 3766 1544
rect 3946 1492 3948 1544
rect 4010 1492 4022 1544
rect 3684 1490 3708 1492
rect 3764 1490 3788 1492
rect 3844 1490 3868 1492
rect 3924 1490 3948 1492
rect 4004 1490 4028 1492
rect 4084 1490 4126 1546
rect 4428 1543 4434 1595
rect 4486 1543 4492 1595
rect 3586 1448 4126 1490
rect 3446 1395 3499 1401
rect 156 603 211 1228
rect 260 774 315 1390
rect 3446 1343 3447 1395
rect 4441 1379 4480 1543
rect 5004 1401 5046 1672
rect 4999 1395 5051 1401
rect 3446 1337 3499 1343
rect 4999 1337 5051 1343
rect 1230 1009 1762 1050
rect 1230 953 1270 1009
rect 1326 1007 1350 1009
rect 1406 1007 1430 1009
rect 1486 1007 1510 1009
rect 1566 1007 1590 1009
rect 1646 1007 1670 1009
rect 1332 955 1344 1007
rect 1406 955 1408 1007
rect 1588 955 1590 1007
rect 1652 955 1664 1007
rect 1326 953 1350 955
rect 1406 953 1430 955
rect 1486 953 1510 955
rect 1566 953 1590 955
rect 1646 953 1670 955
rect 1726 953 1762 1009
rect 442 936 494 942
rect 582 934 638 940
rect 494 932 858 934
rect 494 884 584 932
rect 442 880 584 884
rect 636 880 858 932
rect 1230 910 1762 953
rect 2641 892 2709 900
rect 442 878 1150 880
rect 582 872 638 878
rect 802 872 1150 878
rect 2641 872 2651 892
rect 802 840 2651 872
rect 2703 840 2709 892
rect 802 828 2709 840
rect 802 824 1150 828
rect 734 782 786 788
rect 254 719 260 774
rect 315 719 321 774
rect 1278 783 2733 792
rect 3150 787 3202 793
rect 1278 778 3150 783
rect 786 748 3150 778
rect 786 734 1322 748
rect 2733 739 3150 748
rect 734 724 786 730
rect 3150 729 3202 735
rect 1812 702 1872 713
rect 886 690 938 696
rect 1812 691 1814 702
rect 938 679 1124 686
rect 1481 679 1814 691
rect 938 657 1814 679
rect 938 645 1515 657
rect 1812 646 1814 657
rect 1870 691 1872 702
rect 1870 657 1873 691
rect 1870 646 1872 657
rect 938 642 1124 645
rect 886 632 938 638
rect 1812 635 1872 646
rect 3446 627 3487 1337
rect 4911 1173 4917 1225
rect 4969 1173 4975 1225
rect 4626 1106 4678 1112
rect 4929 1100 4957 1173
rect 5004 1142 5046 1337
rect 5084 1142 5126 1672
rect 5164 1142 5206 1672
rect 5244 1142 5286 1672
rect 5324 1142 5366 1672
rect 5404 1142 5446 1672
rect 6702 1668 6754 1674
rect 6856 1670 6908 1676
rect 5544 1546 6084 1588
rect 5544 1490 5586 1546
rect 5642 1544 5666 1546
rect 5722 1544 5746 1546
rect 5802 1544 5826 1546
rect 5882 1544 5906 1546
rect 5962 1544 5986 1546
rect 5648 1492 5660 1544
rect 5722 1492 5724 1544
rect 5904 1492 5906 1544
rect 5968 1492 5980 1544
rect 5642 1490 5666 1492
rect 5722 1490 5746 1492
rect 5802 1490 5826 1492
rect 5882 1490 5906 1492
rect 5962 1490 5986 1492
rect 6042 1490 6084 1546
rect 6386 1544 6392 1596
rect 6444 1544 6450 1596
rect 5544 1448 6084 1490
rect 6400 1380 6438 1544
rect 4678 1061 4957 1100
rect 3606 1008 4146 1050
rect 4626 1048 4678 1054
rect 3606 952 3648 1008
rect 3704 1006 3728 1008
rect 3784 1006 3808 1008
rect 3864 1006 3888 1008
rect 3944 1006 3968 1008
rect 4024 1006 4048 1008
rect 3710 954 3722 1006
rect 3784 954 3786 1006
rect 3966 954 3968 1006
rect 4030 954 4042 1006
rect 3704 952 3728 954
rect 3784 952 3808 954
rect 3864 952 3888 954
rect 3944 952 3968 954
rect 4024 952 4048 954
rect 4104 952 4146 1008
rect 3606 910 4146 952
rect 4173 781 4228 787
rect 4898 781 4950 784
rect 4173 779 4966 781
rect 4173 727 4174 779
rect 4226 778 4966 779
rect 4226 727 4898 778
rect 4173 726 4898 727
rect 4950 726 4966 778
rect 4173 720 4228 726
rect 4898 720 4950 726
rect 3443 621 3495 627
rect 1036 603 1091 609
rect 156 601 1091 603
rect 156 549 1037 601
rect 1089 549 1091 601
rect 156 548 1091 549
rect 1036 542 1091 548
rect 1636 604 1696 610
rect 2149 604 2207 613
rect 1636 601 2207 604
rect 2720 601 2780 606
rect 1636 600 2780 601
rect 1636 548 1640 600
rect 1692 598 2790 600
rect 1692 548 2152 598
rect 1636 546 2152 548
rect 2204 596 2790 598
rect 2204 546 2724 596
rect 1636 544 2724 546
rect 2776 544 2790 596
rect 1636 538 1696 544
rect 2149 543 2790 544
rect 2149 531 2207 543
rect 2720 540 2790 543
rect 3144 542 3150 594
rect 3202 542 3208 594
rect 3858 612 3910 618
rect 3443 563 3495 569
rect 3857 563 3858 606
rect 2720 534 2780 540
rect 2650 500 2698 504
rect 260 489 315 495
rect 1130 490 1182 496
rect 315 486 501 489
rect 315 442 1130 486
rect 315 434 501 442
rect 1902 490 1954 496
rect 2404 492 2456 494
rect 1182 442 1902 486
rect 260 428 315 434
rect 1130 432 1182 438
rect 1902 432 1954 438
rect 2391 490 2469 492
rect 2391 434 2402 490
rect 2458 434 2469 490
rect 2642 448 2648 500
rect 2700 496 2706 500
rect 3152 496 3196 542
rect 3446 524 3487 563
rect 4504 571 4510 623
rect 4562 571 4568 623
rect 3858 554 3910 560
rect 2700 452 3196 496
rect 3861 507 3900 554
rect 4519 507 4553 571
rect 3861 468 4555 507
rect 4744 498 4796 504
rect 2700 448 2706 452
rect 2391 432 2469 434
rect 2404 430 2456 432
rect 2650 408 2694 448
rect 4897 500 4949 506
rect 4796 458 4897 487
rect 26 245 94 254
rect 156 181 211 370
rect 254 334 260 390
rect 316 334 322 390
rect 156 175 214 181
rect 156 121 160 175
rect 159 0 214 121
rect 260 162 316 334
rect 1206 307 1842 360
rect 1206 305 1256 307
rect 1312 305 1336 307
rect 1392 305 1416 307
rect 1472 305 1496 307
rect 1552 305 1576 307
rect 1632 305 1656 307
rect 1712 305 1736 307
rect 1792 305 1842 307
rect 1206 253 1242 305
rect 1486 253 1496 305
rect 1552 253 1562 305
rect 1806 253 1842 305
rect 1206 251 1256 253
rect 1312 251 1336 253
rect 1392 251 1416 253
rect 1472 251 1496 253
rect 1552 251 1576 253
rect 1632 251 1656 253
rect 1712 251 1736 253
rect 1792 251 1842 253
rect 1206 220 1842 251
rect 3446 173 3487 444
rect 4744 440 4796 446
rect 4897 442 4949 448
rect 3586 318 4126 360
rect 3586 262 3628 318
rect 3684 316 3708 318
rect 3764 316 3788 318
rect 3844 316 3868 318
rect 3924 316 3948 318
rect 4004 316 4028 318
rect 3690 264 3702 316
rect 3764 264 3766 316
rect 3946 264 3948 316
rect 4010 264 4022 316
rect 3684 262 3708 264
rect 3764 262 3788 264
rect 3844 262 3868 264
rect 3924 262 3948 264
rect 4004 262 4028 264
rect 4084 262 4126 318
rect 4428 315 4434 367
rect 4486 315 4492 367
rect 3586 220 4126 262
rect 3446 167 3499 173
rect 260 0 315 162
rect 3446 115 3447 167
rect 4441 151 4480 315
rect 3446 109 3499 115
rect 3446 0 3487 109
<< via2 >>
rect -76 2166 -8 2234
rect 1270 2235 1326 2237
rect 1350 2235 1406 2237
rect 1430 2235 1486 2237
rect 1510 2235 1566 2237
rect 1590 2235 1646 2237
rect 1670 2235 1726 2237
rect 1270 2183 1280 2235
rect 1280 2183 1326 2235
rect 1350 2183 1396 2235
rect 1396 2183 1406 2235
rect 1430 2183 1460 2235
rect 1460 2183 1472 2235
rect 1472 2183 1486 2235
rect 1510 2183 1524 2235
rect 1524 2183 1536 2235
rect 1536 2183 1566 2235
rect 1590 2183 1600 2235
rect 1600 2183 1646 2235
rect 1670 2183 1716 2235
rect 1716 2183 1726 2235
rect 1270 2181 1326 2183
rect 1350 2181 1406 2183
rect 1430 2181 1486 2183
rect 1510 2181 1566 2183
rect 1590 2181 1646 2183
rect 1670 2181 1726 2183
rect 1814 1929 1870 1930
rect 1814 1877 1817 1929
rect 1817 1877 1869 1929
rect 1869 1877 1870 1929
rect 1814 1874 1870 1877
rect 3648 2234 3704 2236
rect 3728 2234 3784 2236
rect 3808 2234 3864 2236
rect 3888 2234 3944 2236
rect 3968 2234 4024 2236
rect 4048 2234 4104 2236
rect 3648 2182 3658 2234
rect 3658 2182 3704 2234
rect 3728 2182 3774 2234
rect 3774 2182 3784 2234
rect 3808 2182 3838 2234
rect 3838 2182 3850 2234
rect 3850 2182 3864 2234
rect 3888 2182 3902 2234
rect 3902 2182 3914 2234
rect 3914 2182 3944 2234
rect 3968 2182 3978 2234
rect 3978 2182 4024 2234
rect 4048 2182 4094 2234
rect 4094 2182 4104 2234
rect 3648 2180 3704 2182
rect 3728 2180 3784 2182
rect 3808 2180 3864 2182
rect 3888 2180 3944 2182
rect 3968 2180 4024 2182
rect 4048 2180 4104 2182
rect 2402 1716 2458 1718
rect 2402 1664 2404 1716
rect 2404 1664 2456 1716
rect 2456 1664 2458 1716
rect 2402 1662 2458 1664
rect 5606 2234 5662 2236
rect 5686 2234 5742 2236
rect 5766 2234 5822 2236
rect 5846 2234 5902 2236
rect 5926 2234 5982 2236
rect 6006 2234 6062 2236
rect 5606 2182 5616 2234
rect 5616 2182 5662 2234
rect 5686 2182 5732 2234
rect 5732 2182 5742 2234
rect 5766 2182 5796 2234
rect 5796 2182 5808 2234
rect 5808 2182 5822 2234
rect 5846 2182 5860 2234
rect 5860 2182 5872 2234
rect 5872 2182 5902 2234
rect 5926 2182 5936 2234
rect 5936 2182 5982 2234
rect 6006 2182 6052 2234
rect 6052 2182 6062 2234
rect 5606 2180 5662 2182
rect 5686 2180 5742 2182
rect 5766 2180 5822 2182
rect 5846 2180 5902 2182
rect 5926 2180 5982 2182
rect 6006 2180 6062 2182
rect -76 960 -8 1028
rect 26 1490 94 1558
rect 1256 1533 1312 1535
rect 1336 1533 1392 1535
rect 1416 1533 1472 1535
rect 1496 1533 1552 1535
rect 1576 1533 1632 1535
rect 1656 1533 1712 1535
rect 1736 1533 1792 1535
rect 1256 1481 1294 1533
rect 1294 1481 1306 1533
rect 1306 1481 1312 1533
rect 1336 1481 1358 1533
rect 1358 1481 1370 1533
rect 1370 1481 1392 1533
rect 1416 1481 1422 1533
rect 1422 1481 1434 1533
rect 1434 1481 1472 1533
rect 1496 1481 1498 1533
rect 1498 1481 1550 1533
rect 1550 1481 1552 1533
rect 1576 1481 1614 1533
rect 1614 1481 1626 1533
rect 1626 1481 1632 1533
rect 1656 1481 1678 1533
rect 1678 1481 1690 1533
rect 1690 1481 1712 1533
rect 1736 1481 1742 1533
rect 1742 1481 1754 1533
rect 1754 1481 1792 1533
rect 1256 1479 1312 1481
rect 1336 1479 1392 1481
rect 1416 1479 1472 1481
rect 1496 1479 1552 1481
rect 1576 1479 1632 1481
rect 1656 1479 1712 1481
rect 1736 1479 1792 1481
rect 3628 1544 3684 1546
rect 3708 1544 3764 1546
rect 3788 1544 3844 1546
rect 3868 1544 3924 1546
rect 3948 1544 4004 1546
rect 4028 1544 4084 1546
rect 3628 1492 3638 1544
rect 3638 1492 3684 1544
rect 3708 1492 3754 1544
rect 3754 1492 3764 1544
rect 3788 1492 3818 1544
rect 3818 1492 3830 1544
rect 3830 1492 3844 1544
rect 3868 1492 3882 1544
rect 3882 1492 3894 1544
rect 3894 1492 3924 1544
rect 3948 1492 3958 1544
rect 3958 1492 4004 1544
rect 4028 1492 4074 1544
rect 4074 1492 4084 1544
rect 3628 1490 3684 1492
rect 3708 1490 3764 1492
rect 3788 1490 3844 1492
rect 3868 1490 3924 1492
rect 3948 1490 4004 1492
rect 4028 1490 4084 1492
rect 1270 1007 1326 1009
rect 1350 1007 1406 1009
rect 1430 1007 1486 1009
rect 1510 1007 1566 1009
rect 1590 1007 1646 1009
rect 1670 1007 1726 1009
rect 1270 955 1280 1007
rect 1280 955 1326 1007
rect 1350 955 1396 1007
rect 1396 955 1406 1007
rect 1430 955 1460 1007
rect 1460 955 1472 1007
rect 1472 955 1486 1007
rect 1510 955 1524 1007
rect 1524 955 1536 1007
rect 1536 955 1566 1007
rect 1590 955 1600 1007
rect 1600 955 1646 1007
rect 1670 955 1716 1007
rect 1716 955 1726 1007
rect 1270 953 1326 955
rect 1350 953 1406 955
rect 1430 953 1486 955
rect 1510 953 1566 955
rect 1590 953 1646 955
rect 1670 953 1726 955
rect 1814 701 1870 702
rect 1814 649 1817 701
rect 1817 649 1869 701
rect 1869 649 1870 701
rect 1814 646 1870 649
rect 5586 1544 5642 1546
rect 5666 1544 5722 1546
rect 5746 1544 5802 1546
rect 5826 1544 5882 1546
rect 5906 1544 5962 1546
rect 5986 1544 6042 1546
rect 5586 1492 5596 1544
rect 5596 1492 5642 1544
rect 5666 1492 5712 1544
rect 5712 1492 5722 1544
rect 5746 1492 5776 1544
rect 5776 1492 5788 1544
rect 5788 1492 5802 1544
rect 5826 1492 5840 1544
rect 5840 1492 5852 1544
rect 5852 1492 5882 1544
rect 5906 1492 5916 1544
rect 5916 1492 5962 1544
rect 5986 1492 6032 1544
rect 6032 1492 6042 1544
rect 5586 1490 5642 1492
rect 5666 1490 5722 1492
rect 5746 1490 5802 1492
rect 5826 1490 5882 1492
rect 5906 1490 5962 1492
rect 5986 1490 6042 1492
rect 3648 1006 3704 1008
rect 3728 1006 3784 1008
rect 3808 1006 3864 1008
rect 3888 1006 3944 1008
rect 3968 1006 4024 1008
rect 4048 1006 4104 1008
rect 3648 954 3658 1006
rect 3658 954 3704 1006
rect 3728 954 3774 1006
rect 3774 954 3784 1006
rect 3808 954 3838 1006
rect 3838 954 3850 1006
rect 3850 954 3864 1006
rect 3888 954 3902 1006
rect 3902 954 3914 1006
rect 3914 954 3944 1006
rect 3968 954 3978 1006
rect 3978 954 4024 1006
rect 4048 954 4094 1006
rect 4094 954 4104 1006
rect 3648 952 3704 954
rect 3728 952 3784 954
rect 3808 952 3864 954
rect 3888 952 3944 954
rect 3968 952 4024 954
rect 4048 952 4104 954
rect 2402 488 2458 490
rect 2402 436 2404 488
rect 2404 436 2456 488
rect 2456 436 2458 488
rect 2402 434 2458 436
rect 26 254 94 322
rect 1256 305 1312 307
rect 1336 305 1392 307
rect 1416 305 1472 307
rect 1496 305 1552 307
rect 1576 305 1632 307
rect 1656 305 1712 307
rect 1736 305 1792 307
rect 1256 253 1294 305
rect 1294 253 1306 305
rect 1306 253 1312 305
rect 1336 253 1358 305
rect 1358 253 1370 305
rect 1370 253 1392 305
rect 1416 253 1422 305
rect 1422 253 1434 305
rect 1434 253 1472 305
rect 1496 253 1498 305
rect 1498 253 1550 305
rect 1550 253 1552 305
rect 1576 253 1614 305
rect 1614 253 1626 305
rect 1626 253 1632 305
rect 1656 253 1678 305
rect 1678 253 1690 305
rect 1690 253 1712 305
rect 1736 253 1742 305
rect 1742 253 1754 305
rect 1754 253 1792 305
rect 1256 251 1312 253
rect 1336 251 1392 253
rect 1416 251 1472 253
rect 1496 251 1552 253
rect 1576 251 1632 253
rect 1656 251 1712 253
rect 1736 251 1792 253
rect 3628 316 3684 318
rect 3708 316 3764 318
rect 3788 316 3844 318
rect 3868 316 3924 318
rect 3948 316 4004 318
rect 4028 316 4084 318
rect 3628 264 3638 316
rect 3638 264 3684 316
rect 3708 264 3754 316
rect 3754 264 3764 316
rect 3788 264 3818 316
rect 3818 264 3830 316
rect 3830 264 3844 316
rect 3868 264 3882 316
rect 3882 264 3894 316
rect 3894 264 3924 316
rect 3948 264 3958 316
rect 3958 264 4004 316
rect 4028 264 4074 316
rect 4074 264 4084 316
rect 3628 262 3684 264
rect 3708 262 3764 264
rect 3788 262 3844 264
rect 3868 262 3924 264
rect 3948 262 4004 264
rect 4028 262 4084 264
<< metal3 >>
rect -120 2237 7606 2278
rect -120 2234 1270 2237
rect -120 2166 -76 2234
rect -8 2181 1270 2234
rect 1326 2181 1350 2237
rect 1406 2181 1430 2237
rect 1486 2181 1510 2237
rect 1566 2181 1590 2237
rect 1646 2181 1670 2237
rect 1726 2236 7606 2237
rect 1726 2181 3648 2236
rect -8 2180 3648 2181
rect 3704 2180 3728 2236
rect 3784 2180 3808 2236
rect 3864 2180 3888 2236
rect 3944 2180 3968 2236
rect 4024 2180 4048 2236
rect 4104 2180 5606 2236
rect 5662 2180 5686 2236
rect 5742 2180 5766 2236
rect 5822 2180 5846 2236
rect 5902 2180 5926 2236
rect 5982 2180 6006 2236
rect 6062 2180 7606 2236
rect -8 2166 7606 2180
rect -120 2138 7606 2166
rect 1807 1930 1877 1937
rect 1807 1874 1814 1930
rect 1870 1874 1877 1930
rect 1807 1867 1877 1874
rect 1812 1720 1872 1867
rect 2395 1720 2465 1725
rect 1812 1718 2465 1720
rect 1812 1662 2402 1718
rect 2458 1662 2465 1718
rect 1812 1660 2465 1662
rect 2395 1655 2465 1660
rect -120 1558 7606 1588
rect -120 1490 26 1558
rect 94 1546 7606 1558
rect 94 1535 3628 1546
rect 94 1490 1256 1535
rect -120 1479 1256 1490
rect 1312 1479 1336 1535
rect 1392 1479 1416 1535
rect 1472 1479 1496 1535
rect 1552 1479 1576 1535
rect 1632 1479 1656 1535
rect 1712 1479 1736 1535
rect 1792 1490 3628 1535
rect 3684 1490 3708 1546
rect 3764 1490 3788 1546
rect 3844 1490 3868 1546
rect 3924 1490 3948 1546
rect 4004 1490 4028 1546
rect 4084 1490 5586 1546
rect 5642 1490 5666 1546
rect 5722 1490 5746 1546
rect 5802 1490 5826 1546
rect 5882 1490 5906 1546
rect 5962 1490 5986 1546
rect 6042 1490 7606 1546
rect 1792 1479 7606 1490
rect -120 1448 7606 1479
rect -120 1028 7606 1050
rect -120 960 -76 1028
rect -8 1009 7606 1028
rect -8 960 1270 1009
rect -120 953 1270 960
rect 1326 953 1350 1009
rect 1406 953 1430 1009
rect 1486 953 1510 1009
rect 1566 953 1590 1009
rect 1646 953 1670 1009
rect 1726 1008 7606 1009
rect 1726 953 3648 1008
rect -120 952 3648 953
rect 3704 952 3728 1008
rect 3784 952 3808 1008
rect 3864 952 3888 1008
rect 3944 952 3968 1008
rect 4024 952 4048 1008
rect 4104 952 7606 1008
rect -120 910 7606 952
rect 1807 702 1877 709
rect 1807 646 1814 702
rect 1870 646 1877 702
rect 1807 639 1877 646
rect 1812 492 1872 639
rect 2395 492 2465 497
rect 1812 490 2465 492
rect 1812 434 2402 490
rect 2458 434 2465 490
rect 1812 432 2465 434
rect 2395 427 2465 432
rect -120 322 7606 360
rect -120 254 26 322
rect 94 318 7606 322
rect 94 307 3628 318
rect 94 254 1256 307
rect -120 251 1256 254
rect 1312 251 1336 307
rect 1392 251 1416 307
rect 1472 251 1496 307
rect 1552 251 1576 307
rect 1632 251 1656 307
rect 1712 251 1736 307
rect 1792 262 3628 307
rect 3684 262 3708 318
rect 3764 262 3788 318
rect 3844 262 3868 318
rect 3924 262 3948 318
rect 4004 262 4028 318
rect 4084 262 7606 318
rect 1792 251 7606 262
rect -120 220 7606 251
<< labels >>
rlabel metal3 -100 2234 -100 2234 7 VCC
port 1 w
rlabel metal3 -92 1522 -92 1522 7 VSS
port 2 w
rlabel metal2 184 2430 184 2430 7 D0
port 3 w
rlabel metal2 288 2432 288 2432 7 VREFL
port 4 w
rlabel metal2 186 20 186 20 7 D0_BUF
port 5 w
rlabel metal2 282 12 282 12 7 VREFH
port 6 w
rlabel metal2 3468 2450 3468 2450 7 D1
port 7 w
rlabel metal2 3468 12 3468 12 7 D1_BUF
port 8 w
rlabel metal2 5023 2436 5023 2436 7 D2
port 9 w
rlabel metal2 5023 1290 5023 1290 7 D2_BUF
port 10 w
rlabel metal2 7021 2310 7021 2310 7 VOUT
port 11 w
flabel metal1 5444 1804 5464 1842 7 FreeSans 600 0 0 0 switch_n_3v3_1.DX
flabel metal1 5416 1350 5444 1388 7 FreeSans 600 0 0 0 switch_n_3v3_1.DX_BUF
flabel metal3 6934 2138 6964 2278 3 FreeSans 600 0 0 0 switch_n_3v3_1.VCC
flabel metal3 6934 1448 6964 1588 3 FreeSans 600 0 0 0 switch_n_3v3_1.VSS
flabel metal3 4954 1448 4984 1588 7 FreeSans 600 0 0 0 switch_n_3v3_1.VSS
flabel metal3 4954 2138 4984 2278 7 FreeSans 600 0 0 0 switch_n_3v3_1.VCC
flabel metal2 5024 2354 5024 2354 1 FreeSans 400 0 0 0 switch_n_3v3_1.D2
flabel metal2 5104 2358 5104 2358 1 FreeSans 400 0 0 0 switch_n_3v3_1.D3
flabel metal2 5186 2358 5186 2358 1 FreeSans 400 0 0 0 switch_n_3v3_1.D4
flabel metal2 5266 2360 5266 2360 1 FreeSans 400 0 0 0 switch_n_3v3_1.D5
flabel metal2 5344 2360 5344 2360 1 FreeSans 400 0 0 0 switch_n_3v3_1.D6
flabel metal2 5424 2358 5424 2358 1 FreeSans 400 0 0 0 switch_n_3v3_1.D7
flabel metal1 6398 2302 6438 2326 3 FreeSans 600 0 0 0 switch_n_3v3_1.VOUT
flabel metal2 6400 1380 6438 1404 7 FreeSans 600 0 0 0 switch_n_3v3_1.VOUT
flabel metal1 5754 1778 5754 1778 7 FreeSans 600 0 0 0 switch_n_3v3_1.DX_
flabel metal1 6790 1374 6818 1398 3 FreeSans 600 0 0 0 switch_n_3v3_1.VREFH
flabel metal1 6868 2298 6898 2318 3 FreeSans 600 0 0 0 switch_n_3v3_1.VREFL
rlabel metal3 30 991 30 991 7 2_bit_dac_0[0].VCC
rlabel metal3 48 286 48 286 7 2_bit_dac_0[0].VSS
rlabel metal2 177 1186 177 1186 7 2_bit_dac_0[0].D0
rlabel metal2 288 1186 288 1186 7 2_bit_dac_0[0].VREFL
rlabel metal2 183 36 183 36 7 2_bit_dac_0[0].D0_BUF
rlabel metal2 291 19 291 19 7 2_bit_dac_0[0].VREFH
rlabel metal2 4938 1077 4938 1077 7 2_bit_dac_0[0].VOUT
rlabel metal2 3468 18 3468 18 7 2_bit_dac_0[0].D1_BUF
rlabel metal2 3466 1204 3466 1204 7 2_bit_dac_0[0].D1
flabel metal1 3374 966 3374 966 3 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.VOUTH
flabel metal1 3360 252 3360 252 3 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.VOUTL
flabel metal2 1136 662 1136 662 7 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.R_L
flabel metal1 2544 930 2544 930 3 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.DX_BUF
flabel metal2 1148 756 1148 756 7 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.R_H
flabel metal2 506 578 506 578 7 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.DX
flabel metal2 496 464 496 464 7 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.VREFL
flabel metal2 516 902 516 902 5 FreeSans 400 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.VREFH
flabel metal3 380 220 410 360 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.VSS
flabel metal3 380 910 410 1050 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch2n_3v3_0.VCC
flabel metal1 3486 575 3506 614 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.DX
flabel metal1 3457 121 3485 160 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_BUF
flabel metal3 4976 910 5006 1050 3 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal3 4976 220 5006 360 3 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal1 4440 1074 4479 1099 3 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal2 4441 151 4480 175 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.VOUT
flabel metal1 3796 550 3796 550 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_
flabel metal3 3314 220 3344 360 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.VSS
flabel metal3 3314 910 3344 1050 7 FreeSans 600 0 0 0 2_bit_dac_0[0].switch_n_3v3_v2_0.VCC
flabel metal1 4770 1107 4770 1107 1 FreeSans 480 0 0 40 2_bit_dac_0[0].switch_n_3v3_v2_0.VREFH
flabel metal1 4923 141 4923 141 5 FreeSans 480 0 0 -40 2_bit_dac_0[0].switch_n_3v3_v2_0.VREFL
rlabel metal3 30 2219 30 2219 7 2_bit_dac_0[1].VCC
rlabel metal3 48 1514 48 1514 7 2_bit_dac_0[1].VSS
rlabel metal2 177 2414 177 2414 7 2_bit_dac_0[1].D0
rlabel metal2 288 2414 288 2414 7 2_bit_dac_0[1].VREFL
rlabel metal2 183 1264 183 1264 7 2_bit_dac_0[1].D0_BUF
rlabel metal2 291 1247 291 1247 7 2_bit_dac_0[1].VREFH
rlabel metal2 4938 2305 4938 2305 7 2_bit_dac_0[1].VOUT
rlabel metal2 3468 1246 3468 1246 7 2_bit_dac_0[1].D1_BUF
rlabel metal2 3466 2432 3466 2432 7 2_bit_dac_0[1].D1
flabel metal1 3374 2194 3374 2194 3 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.VOUTH
flabel metal1 3360 1480 3360 1480 3 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.VOUTL
flabel metal2 1136 1890 1136 1890 7 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.R_L
flabel metal1 2544 2158 2544 2158 3 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.DX_BUF
flabel metal2 1148 1984 1148 1984 7 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.R_H
flabel metal2 506 1806 506 1806 7 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.DX
flabel metal2 496 1692 496 1692 7 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.VREFL
flabel metal2 516 2130 516 2130 5 FreeSans 400 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.VREFH
flabel metal3 380 1448 410 1588 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.VSS
flabel metal3 380 2138 410 2278 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch2n_3v3_0.VCC
flabel metal1 3486 1803 3506 1842 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.DX
flabel metal1 3457 1349 3485 1388 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_BUF
flabel metal3 4976 2138 5006 2278 3 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal3 4976 1448 5006 1588 3 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal1 4440 2302 4479 2327 3 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal2 4441 1379 4480 1403 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.VOUT
flabel metal1 3796 1778 3796 1778 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_
flabel metal3 3314 1448 3344 1588 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.VSS
flabel metal3 3314 2138 3344 2278 7 FreeSans 600 0 0 0 2_bit_dac_0[1].switch_n_3v3_v2_0.VCC
flabel metal1 4770 2335 4770 2335 1 FreeSans 480 0 0 40 2_bit_dac_0[1].switch_n_3v3_v2_0.VREFH
flabel metal1 4923 1369 4923 1369 5 FreeSans 480 0 0 -40 2_bit_dac_0[1].switch_n_3v3_v2_0.VREFL
<< end >>
