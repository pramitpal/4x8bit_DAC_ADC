magic
tech sky130A
magscale 1 2
timestamp 1687027365
<< nwell >>
rect -1580 1620 -900 2020
rect -1580 837 -1260 840
rect -1580 660 -1259 837
rect -1580 470 -900 660
<< nmos >>
rect -1122 736 -1082 820
<< pmos >>
rect -1393 675 -1353 775
<< mvnmos >>
rect -1365 1248 -1265 1448
rect -1207 1248 -1107 1448
<< mvpmos >>
rect -1450 1688 -1350 1788
rect -1171 1686 -1071 1786
<< ndiff >>
rect -1180 808 -1122 820
rect -1180 748 -1168 808
rect -1134 748 -1122 808
rect -1180 736 -1122 748
rect -1082 808 -1024 820
rect -1082 748 -1070 808
rect -1036 748 -1024 808
rect -1082 736 -1024 748
<< pdiff >>
rect -1451 763 -1393 775
rect -1451 687 -1439 763
rect -1405 687 -1393 763
rect -1451 675 -1393 687
rect -1353 763 -1295 775
rect -1353 687 -1341 763
rect -1307 687 -1295 763
rect -1353 675 -1295 687
<< mvndiff >>
rect -1423 1436 -1365 1448
rect -1423 1260 -1411 1436
rect -1377 1260 -1365 1436
rect -1423 1248 -1365 1260
rect -1265 1436 -1207 1448
rect -1265 1260 -1253 1436
rect -1219 1260 -1207 1436
rect -1265 1248 -1207 1260
rect -1107 1436 -1049 1448
rect -1107 1260 -1095 1436
rect -1061 1260 -1049 1436
rect -1107 1248 -1049 1260
<< mvpdiff >>
rect -1508 1776 -1450 1788
rect -1508 1700 -1496 1776
rect -1462 1700 -1450 1776
rect -1508 1688 -1450 1700
rect -1350 1776 -1292 1788
rect -1350 1700 -1338 1776
rect -1304 1700 -1292 1776
rect -1350 1688 -1292 1700
rect -1229 1774 -1171 1786
rect -1229 1698 -1217 1774
rect -1183 1698 -1171 1774
rect -1229 1686 -1171 1698
rect -1071 1774 -1013 1786
rect -1071 1698 -1059 1774
rect -1025 1698 -1013 1774
rect -1071 1686 -1013 1698
<< ndiffc >>
rect -1168 748 -1134 808
rect -1070 748 -1036 808
<< pdiffc >>
rect -1439 687 -1405 763
rect -1341 687 -1307 763
<< mvndiffc >>
rect -1411 1260 -1377 1436
rect -1253 1260 -1219 1436
rect -1095 1260 -1061 1436
<< mvpdiffc >>
rect -1496 1700 -1462 1776
rect -1338 1700 -1304 1776
rect -1217 1698 -1183 1774
rect -1059 1698 -1025 1774
<< psubdiff >>
rect -1420 1060 -1040 1080
rect -1420 1000 -1390 1060
rect -1070 1000 -1040 1060
rect -1420 980 -1040 1000
<< nsubdiff >>
rect -1420 600 -1040 620
rect -1420 540 -1390 600
rect -1070 540 -1040 600
rect -1420 520 -1040 540
<< mvnsubdiff >>
rect -1400 1930 -1020 1950
rect -1400 1870 -1370 1930
rect -1050 1870 -1020 1930
rect -1400 1850 -1020 1870
<< psubdiffcont >>
rect -1390 1000 -1070 1060
<< nsubdiffcont >>
rect -1390 540 -1070 600
<< mvnsubdiffcont >>
rect -1370 1870 -1050 1930
<< poly >>
rect -1450 1788 -1350 1814
rect -1171 1786 -1071 1812
rect -1450 1662 -1350 1688
rect -1417 1616 -1382 1662
rect -1171 1660 -1071 1686
rect -1138 1616 -1101 1660
rect -1432 1606 -1366 1616
rect -1432 1572 -1416 1606
rect -1382 1572 -1366 1606
rect -1432 1562 -1366 1572
rect -1152 1606 -1086 1616
rect -1152 1572 -1136 1606
rect -1102 1572 -1086 1606
rect -1152 1562 -1086 1572
rect -1365 1448 -1265 1474
rect -1207 1448 -1107 1474
rect -1365 1222 -1265 1248
rect -1207 1222 -1107 1248
rect -1330 1177 -1290 1222
rect -1170 1177 -1130 1222
rect -1343 1167 -1277 1177
rect -1343 1133 -1327 1167
rect -1293 1133 -1277 1167
rect -1343 1123 -1277 1133
rect -1183 1167 -1117 1177
rect -1183 1133 -1167 1167
rect -1133 1133 -1117 1167
rect -1183 1123 -1117 1133
rect -1406 907 -1340 917
rect -1406 873 -1390 907
rect -1356 873 -1340 907
rect -1406 863 -1340 873
rect -1135 907 -1069 917
rect -1135 873 -1119 907
rect -1085 873 -1069 907
rect -1135 863 -1069 873
rect -1393 775 -1353 863
rect -1122 820 -1082 863
rect -1122 710 -1082 736
rect -1393 649 -1353 675
<< polycont >>
rect -1416 1572 -1382 1606
rect -1136 1572 -1102 1606
rect -1327 1133 -1293 1167
rect -1167 1133 -1133 1167
rect -1390 873 -1356 907
rect -1119 873 -1085 907
<< locali >>
rect -1400 1930 -1020 1950
rect -1400 1870 -1370 1930
rect -1050 1870 -1020 1930
rect -1400 1850 -1020 1870
rect -1496 1776 -1462 1792
rect -1496 1684 -1462 1700
rect -1338 1776 -1304 1792
rect -1217 1774 -1183 1790
rect -1304 1700 -1301 1738
rect -1416 1607 -1382 1622
rect -1338 1608 -1301 1700
rect -1217 1682 -1183 1698
rect -1059 1774 -1025 1790
rect -1059 1682 -1025 1698
rect -1136 1608 -1102 1622
rect -1338 1606 -1100 1608
rect -1338 1572 -1136 1606
rect -1102 1572 -1100 1606
rect -1416 1556 -1382 1572
rect -1338 1571 -1100 1572
rect -1338 1527 -1301 1571
rect -1136 1556 -1102 1571
rect -1411 1436 -1377 1452
rect -1411 1244 -1377 1260
rect -1253 1436 -1219 1452
rect -1253 1244 -1219 1260
rect -1095 1436 -1061 1452
rect -1095 1244 -1061 1260
rect -1327 1170 -1293 1183
rect -1167 1170 -1133 1183
rect -1460 1167 -1290 1170
rect -1460 1133 -1327 1167
rect -1293 1133 -1290 1167
rect -1460 1130 -1290 1133
rect -1500 910 -1460 1130
rect -1327 1117 -1293 1130
rect -1167 1117 -1133 1130
rect -1420 1060 -1040 1080
rect -1420 1000 -1390 1060
rect -1070 1000 -1040 1060
rect -1420 980 -1040 1000
rect -1390 910 -1356 923
rect -1119 910 -1085 923
rect -1500 907 -1082 910
rect -1500 873 -1390 907
rect -1356 873 -1119 907
rect -1085 873 -1082 907
rect -1500 870 -1082 873
rect -1390 857 -1356 870
rect -1119 857 -1085 870
rect -1168 808 -1134 824
rect -1439 763 -1405 779
rect -1439 671 -1405 687
rect -1341 763 -1307 779
rect -1168 732 -1134 748
rect -1070 808 -1036 824
rect -1070 732 -1036 748
rect -1341 671 -1307 687
rect -1420 600 -1040 620
rect -1420 540 -1390 600
rect -1070 540 -1040 600
rect -1420 520 -1040 540
<< viali >>
rect -1370 1870 -1050 1930
rect -1496 1700 -1462 1776
rect -1338 1700 -1304 1776
rect -1217 1698 -1183 1774
rect -1059 1698 -1025 1774
rect -1416 1606 -1381 1607
rect -1416 1572 -1382 1606
rect -1382 1572 -1381 1606
rect -1338 1490 -1301 1527
rect -1411 1260 -1377 1436
rect -1253 1260 -1219 1436
rect -1095 1260 -1061 1436
rect -1500 1130 -1460 1170
rect -1170 1167 -1130 1170
rect -1170 1133 -1167 1167
rect -1167 1133 -1133 1167
rect -1133 1133 -1130 1167
rect -1170 1130 -1130 1133
rect -1390 1000 -1070 1060
rect -1439 687 -1405 763
rect -1341 687 -1307 763
rect -1168 748 -1134 808
rect -1070 748 -1036 808
rect -1390 540 -1070 600
<< metal1 >>
rect -1400 1930 -1020 1950
rect -1400 1906 -1370 1930
rect -1508 1870 -1370 1906
rect -1050 1870 -1020 1930
rect -1508 1854 -1020 1870
rect -1508 1776 -1456 1854
rect -1400 1850 -1020 1854
rect -1502 1700 -1496 1776
rect -1462 1700 -1456 1776
rect -1502 1688 -1456 1700
rect -1344 1776 -1298 1788
rect -1344 1700 -1338 1776
rect -1304 1700 -1298 1776
rect -1226 1775 -1174 1850
rect -1344 1688 -1298 1700
rect -1223 1774 -1177 1775
rect -1223 1698 -1217 1774
rect -1183 1698 -1177 1774
rect -1223 1686 -1177 1698
rect -1065 1774 -1019 1786
rect -1065 1698 -1059 1774
rect -1025 1698 -1019 1774
rect -1065 1686 -1019 1698
rect -1422 1607 -1375 1619
rect -1058 1607 -1023 1686
rect -1422 1572 -1416 1607
rect -1381 1572 -1023 1607
rect -1422 1560 -1375 1572
rect -1344 1527 -1295 1539
rect -1415 1490 -1338 1527
rect -1301 1490 -1295 1527
rect -1415 1448 -1378 1490
rect -1344 1478 -1295 1490
rect -1097 1448 -1062 1572
rect -1417 1436 -1371 1448
rect -1417 1260 -1411 1436
rect -1377 1260 -1371 1436
rect -1417 1248 -1371 1260
rect -1259 1436 -1213 1448
rect -1259 1260 -1253 1436
rect -1219 1267 -1213 1436
rect -1101 1436 -1055 1448
rect -1219 1260 -1212 1267
rect -1259 1248 -1212 1260
rect -1101 1260 -1095 1436
rect -1061 1289 -1055 1436
rect -1024 1289 -1018 1298
rect -1061 1260 -1018 1289
rect -1101 1254 -1018 1260
rect -1101 1248 -1055 1254
rect -1506 1176 -1454 1182
rect -1512 1124 -1506 1176
rect -1454 1124 -1448 1176
rect -1506 1118 -1454 1124
rect -1251 1080 -1212 1248
rect -1024 1246 -1018 1254
rect -966 1246 -960 1298
rect -1176 1170 -1124 1182
rect -1016 1176 -964 1182
rect -1176 1130 -1170 1170
rect -1130 1130 -1016 1170
rect -1176 1118 -1124 1130
rect -1016 1118 -964 1124
rect -1420 1060 -1030 1080
rect -1420 1000 -1390 1060
rect -1070 1000 -1030 1060
rect -1420 980 -1030 1000
rect -1262 894 -1256 946
rect -1204 894 -1198 946
rect -1445 763 -1399 775
rect -1445 687 -1439 763
rect -1405 687 -1399 763
rect -1445 675 -1399 687
rect -1347 770 -1301 775
rect -1250 770 -1210 894
rect -1070 820 -1030 980
rect -1174 808 -1128 820
rect -1174 770 -1168 808
rect -1347 763 -1168 770
rect -1347 687 -1341 763
rect -1307 748 -1168 763
rect -1134 748 -1128 808
rect -1307 736 -1128 748
rect -1076 808 -1030 820
rect -1076 748 -1070 808
rect -1036 748 -1030 808
rect -1076 736 -1030 748
rect -1307 720 -1130 736
rect -1307 687 -1301 720
rect -1347 675 -1301 687
rect -1440 620 -1400 675
rect -1440 600 -1040 620
rect -1440 540 -1390 600
rect -1070 540 -1040 600
rect -1440 520 -1040 540
<< via1 >>
rect -1370 1870 -1050 1930
rect -1506 1170 -1454 1176
rect -1506 1130 -1500 1170
rect -1500 1130 -1460 1170
rect -1460 1130 -1454 1170
rect -1506 1124 -1454 1130
rect -1018 1246 -966 1298
rect -1016 1124 -964 1176
rect -1390 1000 -1070 1060
rect -1256 894 -1204 946
rect -1390 540 -1070 600
<< metal2 >>
rect -1400 1930 -1020 1950
rect -1400 1870 -1370 1930
rect -1050 1870 -1020 1930
rect -1400 1850 -1020 1870
rect -1018 1298 -966 1304
rect -966 1255 -918 1290
rect -1018 1240 -966 1246
rect -1500 1182 -1460 1240
rect -1506 1176 -1454 1182
rect -1520 1130 -1506 1170
rect -1022 1124 -1016 1176
rect -964 1170 -958 1176
rect -964 1130 -956 1170
rect -964 1124 -958 1130
rect -1506 1118 -1454 1124
rect -1420 1060 -1040 1080
rect -1420 1000 -1390 1060
rect -1070 1000 -1040 1060
rect -1420 980 -1040 1000
rect -1256 946 -1204 952
rect -1010 940 -970 1124
rect -1204 900 -970 940
rect -1256 888 -1204 894
rect -1420 600 -1040 620
rect -1420 540 -1390 600
rect -1070 540 -1040 600
rect -1420 520 -1040 540
<< via2 >>
rect -1370 1870 -1050 1930
rect -1390 1000 -1070 1060
rect -1390 540 -1070 600
<< metal3 >>
rect -1580 1930 -900 1950
rect -1580 1870 -1370 1930
rect -1050 1870 -900 1930
rect -1580 1850 -900 1870
rect -1580 1060 -900 1080
rect -1580 1000 -1390 1060
rect -1070 1000 -900 1060
rect -1580 980 -900 1000
rect -1580 600 -900 620
rect -1580 540 -1390 600
rect -1070 540 -900 600
rect -1580 520 -900 540
<< labels >>
flabel metal3 s -1540 570 -1540 570 0 FreeSans 640 0 0 0 VCCD
flabel metal3 s -1540 1030 -1540 1030 0 FreeSans 640 0 0 0 VSSD
flabel metal3 s -1550 1910 -1550 1910 0 FreeSans 640 0 0 0 VDDA
flabel metal2 s -1480 1220 -1480 1220 0 FreeSans 640 0 0 0 VIN
flabel metal2 s -936 1270 -936 1270 0 FreeSans 640 0 0 0 VOUT
<< end >>
