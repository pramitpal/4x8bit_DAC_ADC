magic
tech sky130A
magscale 1 2
timestamp 1685807414
<< nwell >>
rect -6800 8 -6134 214
rect -6800 -64 -4672 8
rect -6752 -326 -4672 -64
rect -5248 -330 -4934 -326
<< pwell >>
rect -7272 62 -6982 68
rect -7562 -610 -6982 62
rect -6708 -524 -4730 -372
rect -6708 -530 -6095 -524
rect -7562 -616 -7280 -610
rect -6782 -710 -6095 -530
<< mvnmos >>
rect -6624 -498 -6524 -398
rect -6336 -498 -6236 -398
rect -6004 -498 -5904 -398
rect -5662 -498 -5562 -398
rect -5258 -498 -5158 -398
rect -4914 -498 -4814 -398
<< mvpmos >>
rect -6624 -260 -6524 -60
rect -6336 -260 -6236 -60
rect -6004 -260 -5904 -60
rect -5662 -260 -5562 -60
rect -5258 -260 -5158 -60
rect -4914 -260 -4814 -60
<< mvndiff >>
rect -7536 24 -7452 36
rect -7536 -10 -7511 24
rect -7477 -10 -7452 24
rect -7536 -67 -7452 -10
rect -7536 -544 -7452 -487
rect -7536 -578 -7511 -544
rect -7477 -578 -7452 -544
rect -7536 -590 -7452 -578
rect -7390 24 -7306 36
rect -7390 -10 -7365 24
rect -7331 -10 -7306 24
rect -7390 -67 -7306 -10
rect -7390 -544 -7306 -487
rect -7390 -578 -7365 -544
rect -7331 -578 -7306 -544
rect -7390 -590 -7306 -578
rect -7246 30 -7162 42
rect -7246 -4 -7221 30
rect -7187 -4 -7162 30
rect -7246 -61 -7162 -4
rect -7246 -538 -7162 -481
rect -7246 -572 -7221 -538
rect -7187 -572 -7162 -538
rect -7246 -584 -7162 -572
rect -7092 30 -7008 42
rect -7092 -4 -7067 30
rect -7033 -4 -7008 30
rect -7092 -61 -7008 -4
rect -7092 -538 -7008 -481
rect -6682 -431 -6624 -398
rect -6682 -465 -6670 -431
rect -6636 -465 -6624 -431
rect -6682 -498 -6624 -465
rect -6524 -431 -6466 -398
rect -6524 -465 -6512 -431
rect -6478 -465 -6466 -431
rect -6524 -498 -6466 -465
rect -6394 -431 -6336 -398
rect -6394 -465 -6382 -431
rect -6348 -465 -6336 -431
rect -6394 -498 -6336 -465
rect -6236 -431 -6178 -398
rect -6236 -465 -6224 -431
rect -6190 -465 -6178 -431
rect -6236 -498 -6178 -465
rect -6062 -431 -6004 -398
rect -6062 -465 -6050 -431
rect -6016 -465 -6004 -431
rect -6062 -498 -6004 -465
rect -5904 -431 -5846 -398
rect -5904 -465 -5892 -431
rect -5858 -465 -5846 -431
rect -5904 -498 -5846 -465
rect -5720 -431 -5662 -398
rect -5720 -465 -5708 -431
rect -5674 -465 -5662 -431
rect -5720 -498 -5662 -465
rect -5562 -431 -5504 -398
rect -5562 -465 -5550 -431
rect -5516 -465 -5504 -431
rect -5562 -498 -5504 -465
rect -5316 -431 -5258 -398
rect -5316 -465 -5304 -431
rect -5270 -465 -5258 -431
rect -5316 -498 -5258 -465
rect -5158 -431 -5100 -398
rect -5158 -465 -5146 -431
rect -5112 -465 -5100 -431
rect -5158 -498 -5100 -465
rect -4972 -431 -4914 -398
rect -4972 -465 -4960 -431
rect -4926 -465 -4914 -431
rect -4972 -498 -4914 -465
rect -4814 -431 -4756 -398
rect -4814 -465 -4802 -431
rect -4768 -465 -4756 -431
rect -4814 -498 -4756 -465
rect -7092 -572 -7067 -538
rect -7033 -572 -7008 -538
rect -7092 -584 -7008 -572
<< mvpdiff >>
rect -6682 -75 -6624 -60
rect -6682 -109 -6670 -75
rect -6636 -109 -6624 -75
rect -6682 -143 -6624 -109
rect -6682 -177 -6670 -143
rect -6636 -177 -6624 -143
rect -6682 -211 -6624 -177
rect -6682 -245 -6670 -211
rect -6636 -245 -6624 -211
rect -6682 -260 -6624 -245
rect -6524 -75 -6466 -60
rect -6524 -109 -6512 -75
rect -6478 -109 -6466 -75
rect -6524 -143 -6466 -109
rect -6524 -177 -6512 -143
rect -6478 -177 -6466 -143
rect -6524 -211 -6466 -177
rect -6524 -245 -6512 -211
rect -6478 -245 -6466 -211
rect -6524 -260 -6466 -245
rect -6394 -75 -6336 -60
rect -6394 -109 -6382 -75
rect -6348 -109 -6336 -75
rect -6394 -143 -6336 -109
rect -6394 -177 -6382 -143
rect -6348 -177 -6336 -143
rect -6394 -211 -6336 -177
rect -6394 -245 -6382 -211
rect -6348 -245 -6336 -211
rect -6394 -260 -6336 -245
rect -6236 -75 -6178 -60
rect -6236 -109 -6224 -75
rect -6190 -109 -6178 -75
rect -6236 -143 -6178 -109
rect -6236 -177 -6224 -143
rect -6190 -177 -6178 -143
rect -6236 -211 -6178 -177
rect -6236 -245 -6224 -211
rect -6190 -245 -6178 -211
rect -6236 -260 -6178 -245
rect -6062 -75 -6004 -60
rect -6062 -109 -6050 -75
rect -6016 -109 -6004 -75
rect -6062 -143 -6004 -109
rect -6062 -177 -6050 -143
rect -6016 -177 -6004 -143
rect -6062 -211 -6004 -177
rect -6062 -245 -6050 -211
rect -6016 -245 -6004 -211
rect -6062 -260 -6004 -245
rect -5904 -75 -5846 -60
rect -5904 -109 -5892 -75
rect -5858 -109 -5846 -75
rect -5904 -143 -5846 -109
rect -5904 -177 -5892 -143
rect -5858 -177 -5846 -143
rect -5904 -211 -5846 -177
rect -5904 -245 -5892 -211
rect -5858 -245 -5846 -211
rect -5904 -260 -5846 -245
rect -5720 -75 -5662 -60
rect -5720 -109 -5708 -75
rect -5674 -109 -5662 -75
rect -5720 -143 -5662 -109
rect -5720 -177 -5708 -143
rect -5674 -177 -5662 -143
rect -5720 -211 -5662 -177
rect -5720 -245 -5708 -211
rect -5674 -245 -5662 -211
rect -5720 -260 -5662 -245
rect -5562 -75 -5504 -60
rect -5562 -109 -5550 -75
rect -5516 -109 -5504 -75
rect -5562 -143 -5504 -109
rect -5562 -177 -5550 -143
rect -5516 -177 -5504 -143
rect -5562 -211 -5504 -177
rect -5562 -245 -5550 -211
rect -5516 -245 -5504 -211
rect -5562 -260 -5504 -245
rect -5316 -75 -5258 -60
rect -5316 -109 -5304 -75
rect -5270 -109 -5258 -75
rect -5316 -143 -5258 -109
rect -5316 -177 -5304 -143
rect -5270 -177 -5258 -143
rect -5316 -211 -5258 -177
rect -5316 -245 -5304 -211
rect -5270 -245 -5258 -211
rect -5316 -260 -5258 -245
rect -5158 -75 -5100 -60
rect -5158 -109 -5146 -75
rect -5112 -109 -5100 -75
rect -5158 -143 -5100 -109
rect -5158 -177 -5146 -143
rect -5112 -177 -5100 -143
rect -5158 -211 -5100 -177
rect -5158 -245 -5146 -211
rect -5112 -245 -5100 -211
rect -5158 -260 -5100 -245
rect -4972 -75 -4914 -60
rect -4972 -109 -4960 -75
rect -4926 -109 -4914 -75
rect -4972 -143 -4914 -109
rect -4972 -177 -4960 -143
rect -4926 -177 -4914 -143
rect -4972 -211 -4914 -177
rect -4972 -245 -4960 -211
rect -4926 -245 -4914 -211
rect -4972 -260 -4914 -245
rect -4814 -75 -4756 -60
rect -4814 -109 -4802 -75
rect -4768 -109 -4756 -75
rect -4814 -143 -4756 -109
rect -4814 -177 -4802 -143
rect -4768 -177 -4756 -143
rect -4814 -211 -4756 -177
rect -4814 -245 -4802 -211
rect -4768 -245 -4756 -211
rect -4814 -260 -4756 -245
<< mvndiffc >>
rect -7511 -10 -7477 24
rect -7511 -578 -7477 -544
rect -7365 -10 -7331 24
rect -7365 -578 -7331 -544
rect -7221 -4 -7187 30
rect -7221 -572 -7187 -538
rect -7067 -4 -7033 30
rect -6670 -465 -6636 -431
rect -6512 -465 -6478 -431
rect -6382 -465 -6348 -431
rect -6224 -465 -6190 -431
rect -6050 -465 -6016 -431
rect -5892 -465 -5858 -431
rect -5708 -465 -5674 -431
rect -5550 -465 -5516 -431
rect -5304 -465 -5270 -431
rect -5146 -465 -5112 -431
rect -4960 -465 -4926 -431
rect -4802 -465 -4768 -431
rect -7067 -572 -7033 -538
<< mvpdiffc >>
rect -6670 -109 -6636 -75
rect -6670 -177 -6636 -143
rect -6670 -245 -6636 -211
rect -6512 -109 -6478 -75
rect -6512 -177 -6478 -143
rect -6512 -245 -6478 -211
rect -6382 -109 -6348 -75
rect -6382 -177 -6348 -143
rect -6382 -245 -6348 -211
rect -6224 -109 -6190 -75
rect -6224 -177 -6190 -143
rect -6224 -245 -6190 -211
rect -6050 -109 -6016 -75
rect -6050 -177 -6016 -143
rect -6050 -245 -6016 -211
rect -5892 -109 -5858 -75
rect -5892 -177 -5858 -143
rect -5892 -245 -5858 -211
rect -5708 -109 -5674 -75
rect -5708 -177 -5674 -143
rect -5708 -245 -5674 -211
rect -5550 -109 -5516 -75
rect -5550 -177 -5516 -143
rect -5550 -245 -5516 -211
rect -5304 -109 -5270 -75
rect -5304 -177 -5270 -143
rect -5304 -245 -5270 -211
rect -5146 -109 -5112 -75
rect -5146 -177 -5112 -143
rect -5146 -245 -5112 -211
rect -4960 -109 -4926 -75
rect -4960 -177 -4926 -143
rect -4960 -245 -4926 -211
rect -4802 -109 -4768 -75
rect -4802 -177 -4768 -143
rect -4802 -245 -4768 -211
<< psubdiff >>
rect -6756 -608 -6121 -556
rect -6756 -642 -6727 -608
rect -6693 -642 -6659 -608
rect -6625 -642 -6591 -608
rect -6557 -642 -6523 -608
rect -6489 -642 -6455 -608
rect -6421 -642 -6387 -608
rect -6353 -642 -6319 -608
rect -6285 -642 -6251 -608
rect -6217 -642 -6183 -608
rect -6149 -642 -6121 -608
rect -6756 -684 -6121 -642
<< mvnsubdiff >>
rect -6732 94 -6200 146
rect -6732 60 -6685 94
rect -6651 60 -6617 94
rect -6583 60 -6549 94
rect -6515 60 -6481 94
rect -6447 60 -6413 94
rect -6379 60 -6345 94
rect -6311 60 -6277 94
rect -6243 60 -6200 94
rect -6732 6 -6200 60
<< psubdiffcont >>
rect -6727 -642 -6693 -608
rect -6659 -642 -6625 -608
rect -6591 -642 -6557 -608
rect -6523 -642 -6489 -608
rect -6455 -642 -6421 -608
rect -6387 -642 -6353 -608
rect -6319 -642 -6285 -608
rect -6251 -642 -6217 -608
rect -6183 -642 -6149 -608
<< mvnsubdiffcont >>
rect -6685 60 -6651 94
rect -6617 60 -6583 94
rect -6549 60 -6515 94
rect -6481 60 -6447 94
rect -6413 60 -6379 94
rect -6345 60 -6311 94
rect -6277 60 -6243 94
<< poly >>
rect -6624 -60 -6524 -34
rect -6336 -60 -6236 -34
rect -6004 -60 -5904 -34
rect -5662 -60 -5562 -34
rect -5258 -60 -5158 -34
rect -4914 -60 -4814 -34
rect -6624 -288 -6524 -260
rect -6841 -313 -6524 -288
rect -6841 -347 -6811 -313
rect -6777 -347 -6524 -313
rect -6841 -371 -6524 -347
rect -6624 -398 -6524 -371
rect -6336 -313 -6236 -260
rect -6336 -347 -6307 -313
rect -6273 -347 -6236 -313
rect -6336 -398 -6236 -347
rect -6004 -303 -5904 -260
rect -5662 -282 -5562 -260
rect -5459 -282 -5373 -281
rect -6004 -315 -5755 -303
rect -6004 -349 -5807 -315
rect -5773 -349 -5755 -315
rect -6004 -361 -5755 -349
rect -5662 -305 -5368 -282
rect -5662 -339 -5433 -305
rect -5399 -339 -5368 -305
rect -6004 -398 -5904 -361
rect -5662 -373 -5368 -339
rect -5258 -317 -5158 -260
rect -5258 -351 -5223 -317
rect -5189 -351 -5158 -317
rect -5662 -398 -5562 -373
rect -5258 -398 -5158 -351
rect -5061 -307 -5007 -301
rect -4914 -307 -4814 -260
rect -5061 -317 -4814 -307
rect -5061 -351 -5051 -317
rect -5017 -351 -4814 -317
rect -5061 -361 -4814 -351
rect -5061 -367 -5007 -361
rect -4914 -398 -4814 -361
rect -6624 -524 -6524 -498
rect -6336 -524 -6236 -498
rect -6004 -524 -5904 -498
rect -5662 -524 -5562 -498
rect -5258 -524 -5158 -498
rect -4914 -524 -4814 -498
<< polycont >>
rect -6811 -347 -6777 -313
rect -6307 -347 -6273 -313
rect -5807 -349 -5773 -315
rect -5433 -339 -5399 -305
rect -5223 -351 -5189 -317
rect -5051 -351 -5017 -317
<< mvndiffres >>
rect -7536 -487 -7452 -67
rect -7390 -487 -7306 -67
rect -7246 -481 -7162 -61
rect -7092 -481 -7008 -61
<< locali >>
rect -6732 94 -6200 146
rect -6732 60 -6697 94
rect -6651 60 -6625 94
rect -6583 60 -6553 94
rect -6515 60 -6481 94
rect -6447 60 -6413 94
rect -6375 60 -6345 94
rect -6303 60 -6277 94
rect -6231 60 -6200 94
rect -7540 -10 -7511 24
rect -7477 -10 -7448 24
rect -7394 -10 -7365 24
rect -7331 -10 -7302 24
rect -7250 -4 -7221 30
rect -7187 -4 -7158 30
rect -7096 -4 -7067 30
rect -7033 -4 -7004 30
rect -6732 6 -6200 60
rect -5453 13 -5007 67
rect -7524 -30 -7511 -10
rect -7477 -30 -7464 -10
rect -7524 -50 -7464 -30
rect -7378 -30 -7365 -10
rect -7331 -30 -7318 -10
rect -7378 -50 -7318 -30
rect -7234 -24 -7221 -4
rect -7187 -24 -7174 -4
rect -7234 -44 -7174 -24
rect -7080 -24 -7067 -4
rect -7033 -24 -7020 -4
rect -7080 -44 -7020 -24
rect -6670 -75 -6636 -56
rect -6670 -143 -6636 -141
rect -6670 -179 -6636 -177
rect -6670 -264 -6636 -245
rect -6512 -75 -6478 -56
rect -6512 -143 -6478 -141
rect -6512 -179 -6478 -177
rect -6512 -264 -6478 -245
rect -6382 -75 -6348 -56
rect -6382 -143 -6348 -141
rect -6382 -179 -6348 -177
rect -6382 -264 -6348 -245
rect -6224 -75 -6190 -56
rect -6224 -143 -6190 -141
rect -6224 -179 -6190 -177
rect -6224 -264 -6190 -245
rect -6050 -75 -6016 -56
rect -6050 -143 -6016 -141
rect -6050 -179 -6016 -177
rect -6050 -264 -6016 -245
rect -5892 -75 -5858 -56
rect -5892 -143 -5858 -141
rect -5892 -179 -5858 -177
rect -5892 -264 -5858 -245
rect -5708 -75 -5674 -56
rect -5708 -143 -5674 -141
rect -5708 -179 -5674 -177
rect -5708 -264 -5674 -245
rect -5550 -75 -5516 -56
rect -5453 -137 -5399 13
rect -5304 -75 -5270 -56
rect -5550 -143 -5516 -141
rect -5550 -179 -5516 -177
rect -5550 -264 -5516 -245
rect -5455 -159 -5377 -137
rect -5455 -193 -5433 -159
rect -5399 -193 -5377 -159
rect -6825 -294 -6762 -282
rect -6829 -313 -6758 -294
rect -5455 -297 -5377 -193
rect -5304 -143 -5270 -141
rect -5304 -179 -5270 -177
rect -5304 -264 -5270 -245
rect -5146 -75 -5112 -56
rect -5146 -143 -5112 -141
rect -5146 -179 -5112 -177
rect -5146 -264 -5112 -245
rect -6307 -306 -6273 -297
rect -5809 -303 -5771 -297
rect -6829 -347 -6811 -313
rect -6777 -347 -6758 -313
rect -6829 -365 -6758 -347
rect -6314 -313 -6266 -306
rect -6314 -347 -6307 -313
rect -6273 -347 -6266 -313
rect -6314 -354 -6266 -347
rect -5819 -315 -5761 -303
rect -5819 -349 -5807 -315
rect -5773 -349 -5761 -315
rect -5465 -305 -5367 -297
rect -5465 -339 -5433 -305
rect -5399 -339 -5367 -305
rect -5223 -310 -5189 -301
rect -5465 -346 -5367 -339
rect -5230 -317 -5182 -310
rect -5061 -317 -5007 13
rect -4960 -75 -4926 -56
rect -4960 -143 -4926 -141
rect -4960 -179 -4926 -177
rect -4960 -264 -4926 -245
rect -4802 -75 -4768 -56
rect -4802 -143 -4768 -141
rect -4802 -179 -4768 -177
rect -4802 -264 -4768 -245
rect -6307 -363 -6273 -354
rect -5819 -361 -5761 -349
rect -5455 -360 -5377 -346
rect -5230 -351 -5223 -317
rect -5189 -351 -5182 -317
rect -5067 -351 -5051 -317
rect -5017 -351 -5001 -317
rect -5230 -358 -5182 -351
rect -6825 -377 -6762 -365
rect -5809 -367 -5771 -361
rect -5223 -367 -5189 -358
rect -5061 -361 -5007 -351
rect -6670 -431 -6636 -394
rect -7524 -524 -7464 -504
rect -7524 -544 -7511 -524
rect -7477 -544 -7464 -524
rect -7378 -524 -7318 -504
rect -7378 -544 -7365 -524
rect -7331 -544 -7318 -524
rect -7234 -518 -7174 -498
rect -7234 -538 -7221 -518
rect -7187 -538 -7174 -518
rect -7080 -518 -7020 -498
rect -6670 -502 -6636 -465
rect -6512 -431 -6478 -394
rect -6512 -502 -6478 -465
rect -6382 -431 -6348 -394
rect -6382 -502 -6348 -465
rect -6224 -431 -6190 -394
rect -6224 -502 -6190 -465
rect -6050 -431 -6016 -394
rect -6050 -502 -6016 -465
rect -5892 -431 -5858 -394
rect -5892 -502 -5858 -465
rect -5728 -431 -5660 -388
rect -5728 -465 -5708 -431
rect -5674 -465 -5660 -431
rect -7080 -538 -7067 -518
rect -7033 -538 -7020 -518
rect -7540 -578 -7511 -544
rect -7477 -578 -7448 -544
rect -7394 -578 -7365 -544
rect -7331 -578 -7302 -544
rect -7250 -572 -7221 -538
rect -7187 -572 -7158 -538
rect -7096 -572 -7067 -538
rect -7033 -572 -7004 -538
rect -6756 -608 -6120 -544
rect -6756 -642 -6727 -608
rect -6673 -642 -6659 -608
rect -6601 -642 -6591 -608
rect -6529 -642 -6523 -608
rect -6457 -642 -6455 -608
rect -6421 -642 -6419 -608
rect -6353 -642 -6347 -608
rect -6285 -642 -6275 -608
rect -6217 -642 -6203 -608
rect -6149 -642 -6120 -608
rect -6756 -684 -6120 -642
rect -5728 -633 -5660 -465
rect -5550 -431 -5516 -394
rect -5550 -502 -5516 -465
rect -5304 -431 -5270 -394
rect -5304 -502 -5270 -465
rect -5146 -431 -5112 -394
rect -5146 -502 -5112 -465
rect -4960 -431 -4926 -394
rect -4960 -502 -4926 -465
rect -4802 -431 -4768 -394
rect -4802 -502 -4768 -465
rect -5728 -667 -5711 -633
rect -5677 -667 -5660 -633
rect -5728 -684 -5660 -667
<< viali >>
rect -6697 60 -6685 94
rect -6685 60 -6663 94
rect -6625 60 -6617 94
rect -6617 60 -6591 94
rect -6553 60 -6549 94
rect -6549 60 -6519 94
rect -6481 60 -6447 94
rect -6409 60 -6379 94
rect -6379 60 -6375 94
rect -6337 60 -6311 94
rect -6311 60 -6303 94
rect -6265 60 -6243 94
rect -6243 60 -6231 94
rect -7511 -10 -7477 4
rect -7365 -10 -7331 4
rect -7221 -4 -7187 10
rect -7067 -4 -7033 10
rect -7511 -30 -7477 -10
rect -7365 -30 -7331 -10
rect -7221 -24 -7187 -4
rect -7067 -24 -7033 -4
rect -6670 -109 -6636 -107
rect -6670 -141 -6636 -109
rect -6670 -211 -6636 -179
rect -6670 -213 -6636 -211
rect -6512 -109 -6478 -107
rect -6512 -141 -6478 -109
rect -6512 -211 -6478 -179
rect -6512 -213 -6478 -211
rect -6382 -109 -6348 -107
rect -6382 -141 -6348 -109
rect -6382 -211 -6348 -179
rect -6382 -213 -6348 -211
rect -6224 -109 -6190 -107
rect -6224 -141 -6190 -109
rect -6224 -211 -6190 -179
rect -6224 -213 -6190 -211
rect -6050 -109 -6016 -107
rect -6050 -141 -6016 -109
rect -6050 -211 -6016 -179
rect -6050 -213 -6016 -211
rect -5892 -109 -5858 -107
rect -5892 -141 -5858 -109
rect -5892 -211 -5858 -179
rect -5892 -213 -5858 -211
rect -5708 -109 -5674 -107
rect -5708 -141 -5674 -109
rect -5708 -211 -5674 -179
rect -5708 -213 -5674 -211
rect -5550 -109 -5516 -107
rect -5550 -141 -5516 -109
rect -5304 -109 -5270 -107
rect -5550 -211 -5516 -179
rect -5550 -213 -5516 -211
rect -5433 -193 -5399 -159
rect -5304 -141 -5270 -109
rect -5304 -211 -5270 -179
rect -5304 -213 -5270 -211
rect -5146 -109 -5112 -107
rect -5146 -141 -5112 -109
rect -5146 -211 -5112 -179
rect -5146 -213 -5112 -211
rect -6811 -347 -6777 -313
rect -6307 -347 -6273 -313
rect -5807 -349 -5773 -315
rect -4960 -109 -4926 -107
rect -4960 -141 -4926 -109
rect -4960 -211 -4926 -179
rect -4960 -213 -4926 -211
rect -4802 -109 -4768 -107
rect -4802 -141 -4768 -109
rect -4802 -211 -4768 -179
rect -4802 -213 -4768 -211
rect -5223 -351 -5189 -317
rect -6670 -465 -6636 -431
rect -7511 -544 -7477 -524
rect -7365 -544 -7331 -524
rect -7221 -538 -7187 -518
rect -6512 -465 -6478 -431
rect -6382 -465 -6348 -431
rect -6224 -465 -6190 -431
rect -6050 -465 -6016 -431
rect -5892 -465 -5858 -431
rect -5708 -465 -5674 -431
rect -7067 -538 -7033 -518
rect -7511 -558 -7477 -544
rect -7365 -558 -7331 -544
rect -7221 -552 -7187 -538
rect -7067 -552 -7033 -538
rect -6707 -642 -6693 -608
rect -6693 -642 -6673 -608
rect -6635 -642 -6625 -608
rect -6625 -642 -6601 -608
rect -6563 -642 -6557 -608
rect -6557 -642 -6529 -608
rect -6491 -642 -6489 -608
rect -6489 -642 -6457 -608
rect -6419 -642 -6387 -608
rect -6387 -642 -6385 -608
rect -6347 -642 -6319 -608
rect -6319 -642 -6313 -608
rect -6275 -642 -6251 -608
rect -6251 -642 -6241 -608
rect -6203 -642 -6183 -608
rect -6183 -642 -6169 -608
rect -5550 -465 -5516 -431
rect -5304 -465 -5270 -431
rect -5146 -465 -5112 -431
rect -4960 -465 -4926 -431
rect -4802 -465 -4768 -431
rect -5711 -667 -5677 -633
<< metal1 >>
rect -6732 103 -6200 146
rect -6732 94 -6682 103
rect -6630 94 -6618 103
rect -6732 60 -6697 94
rect -6630 60 -6625 94
rect -6732 51 -6682 60
rect -6630 51 -6618 60
rect -6566 51 -6554 103
rect -6502 51 -6490 103
rect -6438 51 -6426 103
rect -6374 51 -6362 103
rect -6310 94 -6298 103
rect -6246 94 -6200 103
rect -6303 60 -6298 94
rect -6231 60 -6200 94
rect -6310 51 -6298 60
rect -6246 51 -6200 60
rect -7530 32 -7458 36
rect -7530 -20 -7520 32
rect -7468 -20 -7458 32
rect -7384 30 -7312 36
rect -7530 -30 -7511 -20
rect -7477 -30 -7458 -20
rect -7398 28 -7312 30
rect -7398 -24 -7378 28
rect -7326 -24 -7312 28
rect -7398 -26 -7365 -24
rect -7530 -62 -7458 -30
rect -7384 -30 -7365 -26
rect -7331 -30 -7312 -24
rect -7384 -62 -7312 -30
rect -7240 10 -7168 42
rect -7240 -24 -7221 10
rect -7187 -24 -7168 10
rect -7240 -56 -7168 -24
rect -7086 10 -7014 42
rect -7086 -24 -7067 10
rect -7033 -24 -7014 10
rect -6732 6 -6200 51
rect -7086 -56 -7014 -24
rect -7516 -102 -7472 -62
rect -7224 -122 -7180 -56
rect -7234 -174 -7228 -122
rect -7176 -174 -7170 -122
rect -7224 -214 -7180 -174
rect -7072 -214 -7028 -56
rect -6673 -60 -6632 6
rect -6387 -60 -6345 6
rect -6139 3 -5393 48
rect -6676 -107 -6630 -60
rect -6676 -141 -6670 -107
rect -6636 -141 -6630 -107
rect -6676 -179 -6630 -141
rect -6676 -213 -6670 -179
rect -6636 -213 -6630 -179
rect -7372 -258 -7180 -214
rect -7372 -492 -7328 -258
rect -7082 -266 -7076 -214
rect -7024 -266 -7018 -214
rect -6676 -260 -6630 -213
rect -6518 -107 -6472 -60
rect -6518 -141 -6512 -107
rect -6478 -141 -6472 -107
rect -6518 -179 -6472 -141
rect -6518 -213 -6512 -179
rect -6478 -213 -6472 -179
rect -6518 -260 -6472 -213
rect -6388 -107 -6342 -60
rect -6388 -141 -6382 -107
rect -6348 -141 -6342 -107
rect -6388 -179 -6342 -141
rect -6388 -213 -6382 -179
rect -6348 -213 -6342 -179
rect -6388 -260 -6342 -213
rect -6230 -63 -6184 -60
rect -6139 -63 -6094 3
rect -6230 -107 -6094 -63
rect -6230 -141 -6224 -107
rect -6190 -108 -6094 -107
rect -6056 -107 -6010 -60
rect -6190 -141 -6184 -108
rect -6230 -179 -6184 -141
rect -6056 -141 -6050 -107
rect -6016 -141 -6010 -107
rect -6056 -176 -6010 -141
rect -6082 -178 -6010 -176
rect -6230 -213 -6224 -179
rect -6190 -213 -6184 -179
rect -6230 -260 -6184 -213
rect -6152 -179 -6010 -178
rect -6152 -203 -6050 -179
rect -6152 -220 -6145 -203
rect -6151 -255 -6145 -220
rect -6093 -213 -6050 -203
rect -6016 -213 -6010 -179
rect -6093 -220 -6010 -213
rect -6093 -255 -6087 -220
rect -6056 -260 -6010 -220
rect -5898 -104 -5852 -60
rect -5714 -104 -5668 -60
rect -5898 -107 -5668 -104
rect -5898 -141 -5892 -107
rect -5858 -141 -5708 -107
rect -5674 -141 -5668 -107
rect -5898 -179 -5668 -141
rect -5898 -213 -5892 -179
rect -5858 -213 -5708 -179
rect -5674 -213 -5668 -179
rect -5898 -230 -5668 -213
rect -5898 -260 -5852 -230
rect -5714 -260 -5668 -230
rect -5556 -107 -5510 -60
rect -5556 -141 -5550 -107
rect -5516 -141 -5510 -107
rect -5438 -131 -5393 3
rect -4962 40 -4569 79
rect -5306 -4 -5264 -3
rect -5322 -12 -5264 -4
rect -5322 -64 -5311 -12
rect -5259 -64 -5253 -12
rect -4962 -60 -4923 40
rect -5322 -107 -5264 -64
rect -5556 -179 -5510 -141
rect -5556 -213 -5550 -179
rect -5516 -213 -5510 -179
rect -5556 -220 -5510 -213
rect -5467 -159 -5365 -131
rect -5467 -193 -5433 -159
rect -5399 -193 -5365 -159
rect -5556 -260 -5506 -220
rect -5467 -221 -5365 -193
rect -5322 -141 -5304 -107
rect -5270 -141 -5264 -107
rect -5322 -179 -5264 -141
rect -5322 -213 -5304 -179
rect -5270 -213 -5264 -179
rect -7072 -320 -7028 -266
rect -6835 -301 -6752 -282
rect -7228 -364 -7028 -320
rect -6932 -303 -6752 -301
rect -6932 -355 -6925 -303
rect -6873 -313 -6752 -303
rect -6873 -347 -6811 -313
rect -6777 -347 -6752 -313
rect -6873 -355 -6752 -347
rect -6932 -356 -6752 -355
rect -7228 -486 -7184 -364
rect -6835 -377 -6752 -356
rect -6512 -294 -6478 -260
rect -6512 -304 -6260 -294
rect -6512 -356 -6322 -304
rect -6270 -356 -6260 -304
rect -6512 -366 -6260 -356
rect -6512 -398 -6472 -366
rect -6227 -398 -6188 -260
rect -5895 -398 -5856 -260
rect -5825 -297 -5755 -291
rect -5825 -306 -5749 -297
rect -5825 -358 -5810 -306
rect -5758 -358 -5749 -306
rect -5825 -367 -5749 -358
rect -5825 -373 -5755 -367
rect -5712 -398 -5673 -260
rect -5550 -294 -5506 -260
rect -5322 -260 -5264 -213
rect -5152 -107 -5106 -60
rect -5152 -141 -5146 -107
rect -5112 -120 -5106 -107
rect -4966 -107 -4920 -60
rect -4966 -120 -4960 -107
rect -5112 -141 -4960 -120
rect -4926 -141 -4920 -107
rect -4808 -107 -4762 -60
rect -4808 -117 -4802 -107
rect -4768 -117 -4762 -107
rect -5152 -179 -4920 -141
rect -4818 -169 -4812 -117
rect -4760 -169 -4754 -117
rect -5152 -213 -5146 -179
rect -5112 -213 -4960 -179
rect -4926 -213 -4920 -179
rect -5152 -230 -4920 -213
rect -5152 -260 -5106 -230
rect -4966 -260 -4920 -230
rect -4808 -179 -4762 -169
rect -4808 -213 -4802 -179
rect -4768 -213 -4762 -179
rect -4808 -260 -4762 -213
rect -5322 -294 -5278 -260
rect -5550 -338 -5424 -294
rect -6838 -418 -6832 -414
rect -6942 -462 -6832 -418
rect -6942 -486 -6898 -462
rect -6838 -466 -6832 -462
rect -6780 -466 -6774 -414
rect -6676 -431 -6630 -398
rect -6676 -465 -6670 -431
rect -6636 -465 -6630 -431
rect -6676 -469 -6630 -465
rect -7530 -524 -7458 -492
rect -7530 -558 -7511 -524
rect -7477 -558 -7458 -524
rect -7530 -590 -7458 -558
rect -7384 -524 -7312 -492
rect -7384 -558 -7365 -524
rect -7331 -558 -7312 -524
rect -7384 -590 -7312 -558
rect -7240 -518 -7168 -486
rect -7240 -552 -7221 -518
rect -7187 -552 -7168 -518
rect -7240 -584 -7168 -552
rect -7086 -518 -6898 -486
rect -7086 -552 -7067 -518
rect -7033 -530 -6898 -518
rect -6681 -498 -6630 -469
rect -6518 -431 -6472 -398
rect -6518 -465 -6512 -431
rect -6478 -465 -6472 -431
rect -6388 -431 -6342 -398
rect -6388 -460 -6382 -431
rect -6518 -498 -6472 -465
rect -6390 -465 -6382 -460
rect -6348 -460 -6342 -431
rect -6230 -431 -6184 -398
rect -6056 -414 -6010 -398
rect -6348 -465 -6340 -460
rect -7033 -552 -7014 -530
rect -6681 -544 -6631 -498
rect -6390 -544 -6340 -465
rect -6230 -465 -6224 -431
rect -6190 -465 -6184 -431
rect -6230 -498 -6184 -465
rect -6066 -466 -6060 -414
rect -6008 -466 -6002 -414
rect -5898 -431 -5852 -398
rect -5898 -465 -5892 -431
rect -5858 -465 -5852 -431
rect -6056 -498 -6010 -466
rect -5898 -498 -5852 -465
rect -5714 -431 -5668 -398
rect -5556 -416 -5510 -398
rect -5714 -465 -5708 -431
rect -5674 -465 -5668 -431
rect -5714 -498 -5668 -465
rect -5564 -468 -5558 -416
rect -5506 -468 -5500 -416
rect -5556 -498 -5510 -468
rect -6056 -530 -6012 -498
rect -5468 -530 -5424 -338
rect -7086 -584 -7014 -552
rect -6756 -599 -6120 -544
rect -6056 -574 -5424 -530
rect -5386 -338 -5278 -294
rect -5248 -308 -5176 -298
rect -5386 -536 -5342 -338
rect -5248 -360 -5238 -308
rect -5186 -360 -5176 -308
rect -5248 -370 -5176 -360
rect -5147 -398 -5108 -260
rect -4962 -398 -4923 -260
rect -4808 -304 -4764 -260
rect -4812 -310 -4760 -304
rect -4812 -368 -4760 -362
rect -5314 -404 -5262 -398
rect -5314 -462 -5304 -456
rect -5310 -465 -5304 -462
rect -5270 -462 -5262 -456
rect -5152 -431 -5106 -398
rect -5270 -465 -5264 -462
rect -5310 -498 -5264 -465
rect -5152 -465 -5146 -431
rect -5112 -465 -5106 -431
rect -5152 -498 -5106 -465
rect -4966 -431 -4920 -398
rect -4966 -465 -4960 -431
rect -4926 -465 -4920 -431
rect -4966 -498 -4920 -465
rect -4808 -431 -4762 -398
rect -4808 -465 -4802 -431
rect -4768 -465 -4762 -431
rect -4808 -498 -4762 -465
rect -4806 -536 -4762 -498
rect -5386 -580 -4762 -536
rect -6756 -651 -6720 -599
rect -6668 -651 -6656 -599
rect -6604 -608 -6592 -599
rect -6540 -608 -6528 -599
rect -6476 -608 -6464 -599
rect -6412 -608 -6400 -599
rect -6348 -608 -6336 -599
rect -6284 -608 -6272 -599
rect -6601 -642 -6592 -608
rect -6529 -642 -6528 -608
rect -6348 -642 -6347 -608
rect -6284 -642 -6275 -608
rect -6604 -651 -6592 -642
rect -6540 -651 -6528 -642
rect -6476 -651 -6464 -642
rect -6412 -651 -6400 -642
rect -6348 -651 -6336 -642
rect -6284 -651 -6272 -642
rect -6220 -651 -6208 -599
rect -6156 -651 -6120 -599
rect -6756 -684 -6120 -651
rect -5734 -629 -5654 -604
rect -5734 -633 -4563 -629
rect -5734 -667 -5711 -633
rect -5677 -667 -4563 -633
rect -5734 -671 -4563 -667
rect -5734 -696 -5654 -671
<< via1 >>
rect -6682 94 -6630 103
rect -6618 94 -6566 103
rect -6682 60 -6663 94
rect -6663 60 -6630 94
rect -6618 60 -6591 94
rect -6591 60 -6566 94
rect -6682 51 -6630 60
rect -6618 51 -6566 60
rect -6554 94 -6502 103
rect -6554 60 -6553 94
rect -6553 60 -6519 94
rect -6519 60 -6502 94
rect -6554 51 -6502 60
rect -6490 94 -6438 103
rect -6490 60 -6481 94
rect -6481 60 -6447 94
rect -6447 60 -6438 94
rect -6490 51 -6438 60
rect -6426 94 -6374 103
rect -6426 60 -6409 94
rect -6409 60 -6375 94
rect -6375 60 -6374 94
rect -6426 51 -6374 60
rect -6362 94 -6310 103
rect -6298 94 -6246 103
rect -6362 60 -6337 94
rect -6337 60 -6310 94
rect -6298 60 -6265 94
rect -6265 60 -6246 94
rect -6362 51 -6310 60
rect -6298 51 -6246 60
rect -7520 4 -7468 32
rect -7520 -20 -7511 4
rect -7511 -20 -7477 4
rect -7477 -20 -7468 4
rect -7378 4 -7326 28
rect -7378 -24 -7365 4
rect -7365 -24 -7331 4
rect -7331 -24 -7326 4
rect -7228 -174 -7176 -122
rect -7076 -266 -7024 -214
rect -6145 -255 -6093 -203
rect -5311 -64 -5259 -12
rect -6925 -355 -6873 -303
rect -6322 -313 -6270 -304
rect -6322 -347 -6307 -313
rect -6307 -347 -6273 -313
rect -6273 -347 -6270 -313
rect -6322 -356 -6270 -347
rect -5810 -315 -5758 -306
rect -5810 -349 -5807 -315
rect -5807 -349 -5773 -315
rect -5773 -349 -5758 -315
rect -5810 -358 -5758 -349
rect -4812 -141 -4802 -117
rect -4802 -141 -4768 -117
rect -4768 -141 -4760 -117
rect -4812 -169 -4760 -141
rect -6832 -466 -6780 -414
rect -6060 -431 -6008 -414
rect -6060 -465 -6050 -431
rect -6050 -465 -6016 -431
rect -6016 -465 -6008 -431
rect -6060 -466 -6008 -465
rect -5558 -431 -5506 -416
rect -5558 -465 -5550 -431
rect -5550 -465 -5516 -431
rect -5516 -465 -5506 -431
rect -5558 -468 -5506 -465
rect -5238 -317 -5186 -308
rect -5238 -351 -5223 -317
rect -5223 -351 -5189 -317
rect -5189 -351 -5186 -317
rect -5238 -360 -5186 -351
rect -4812 -362 -4760 -310
rect -5314 -431 -5262 -404
rect -5314 -456 -5304 -431
rect -5304 -456 -5270 -431
rect -5270 -456 -5262 -431
rect -6720 -608 -6668 -599
rect -6720 -642 -6707 -608
rect -6707 -642 -6673 -608
rect -6673 -642 -6668 -608
rect -6720 -651 -6668 -642
rect -6656 -608 -6604 -599
rect -6592 -608 -6540 -599
rect -6528 -608 -6476 -599
rect -6464 -608 -6412 -599
rect -6400 -608 -6348 -599
rect -6336 -608 -6284 -599
rect -6272 -608 -6220 -599
rect -6656 -642 -6635 -608
rect -6635 -642 -6604 -608
rect -6592 -642 -6563 -608
rect -6563 -642 -6540 -608
rect -6528 -642 -6491 -608
rect -6491 -642 -6476 -608
rect -6464 -642 -6457 -608
rect -6457 -642 -6419 -608
rect -6419 -642 -6412 -608
rect -6400 -642 -6385 -608
rect -6385 -642 -6348 -608
rect -6336 -642 -6313 -608
rect -6313 -642 -6284 -608
rect -6272 -642 -6241 -608
rect -6241 -642 -6220 -608
rect -6656 -651 -6604 -642
rect -6592 -651 -6540 -642
rect -6528 -651 -6476 -642
rect -6464 -651 -6412 -642
rect -6400 -651 -6348 -642
rect -6336 -651 -6284 -642
rect -6272 -651 -6220 -642
rect -6208 -608 -6156 -599
rect -6208 -642 -6203 -608
rect -6203 -642 -6169 -608
rect -6169 -642 -6156 -608
rect -6208 -651 -6156 -642
<< metal2 >>
rect -6732 105 -6200 146
rect -6732 49 -6692 105
rect -6636 103 -6612 105
rect -6556 103 -6532 105
rect -6476 103 -6452 105
rect -6396 103 -6372 105
rect -6316 103 -6292 105
rect -6630 51 -6618 103
rect -6556 51 -6554 103
rect -6374 51 -6372 103
rect -6310 51 -6298 103
rect -6636 49 -6612 51
rect -6556 49 -6532 51
rect -6476 49 -6452 51
rect -6396 49 -6372 51
rect -6316 49 -6292 51
rect -6236 49 -6200 105
rect -7520 32 -7468 38
rect -7380 30 -7324 36
rect -7468 28 -7104 30
rect -7468 -20 -7378 28
rect -7520 -24 -7378 -20
rect -7326 -24 -7104 28
rect -6732 6 -6200 49
rect -5321 -12 -5253 -4
rect -7520 -26 -6812 -24
rect -7380 -32 -7324 -26
rect -7160 -32 -6812 -26
rect -5321 -32 -5311 -12
rect -7160 -64 -5311 -32
rect -5259 -64 -5253 -12
rect -7160 -76 -5253 -64
rect -7160 -80 -6812 -76
rect -7228 -122 -7176 -116
rect -6684 -121 -5229 -112
rect -4812 -117 -4760 -111
rect -6684 -126 -4812 -121
rect -7176 -156 -4812 -126
rect -7176 -170 -6640 -156
rect -5229 -165 -4812 -156
rect -7228 -180 -7176 -174
rect -4812 -175 -4760 -169
rect -6150 -202 -6090 -191
rect -7076 -214 -7024 -208
rect -6150 -213 -6148 -202
rect -7024 -225 -6838 -218
rect -6481 -225 -6148 -213
rect -7024 -247 -6148 -225
rect -7024 -259 -6447 -247
rect -6150 -258 -6148 -247
rect -6092 -213 -6090 -202
rect -6092 -247 -6089 -213
rect -6092 -258 -6090 -247
rect -7024 -262 -6838 -259
rect -7076 -272 -7024 -266
rect -6150 -269 -6090 -258
rect -6926 -301 -6871 -295
rect -7491 -303 -6871 -301
rect -7491 -355 -6925 -303
rect -6873 -355 -6871 -303
rect -7491 -356 -6871 -355
rect -6926 -362 -6871 -356
rect -6326 -300 -6266 -294
rect -5813 -300 -5755 -291
rect -6326 -303 -5755 -300
rect -5242 -303 -5182 -298
rect -6326 -304 -5182 -303
rect -6326 -356 -6322 -304
rect -6270 -306 -5172 -304
rect -6270 -356 -5810 -306
rect -6326 -358 -5810 -356
rect -5758 -308 -5172 -306
rect -5758 -358 -5238 -308
rect -6326 -360 -5238 -358
rect -5186 -360 -5172 -308
rect -6326 -366 -6266 -360
rect -5813 -361 -5172 -360
rect -5813 -373 -5755 -361
rect -5242 -364 -5172 -361
rect -4818 -362 -4812 -310
rect -4760 -362 -4754 -310
rect -5242 -370 -5182 -364
rect -5312 -404 -5264 -400
rect -6832 -414 -6780 -408
rect -7490 -462 -6832 -418
rect -6060 -414 -6008 -408
rect -5558 -412 -5506 -410
rect -6780 -462 -6060 -418
rect -6832 -472 -6780 -466
rect -6060 -472 -6008 -466
rect -5571 -414 -5493 -412
rect -5571 -470 -5560 -414
rect -5504 -470 -5493 -414
rect -5320 -456 -5314 -404
rect -5262 -408 -5256 -404
rect -4810 -408 -4766 -362
rect -5262 -452 -4766 -408
rect -5262 -456 -5256 -452
rect -5571 -472 -5493 -470
rect -5558 -474 -5506 -472
rect -5312 -496 -5268 -456
rect -6756 -597 -6120 -544
rect -6756 -599 -6706 -597
rect -6650 -599 -6626 -597
rect -6570 -599 -6546 -597
rect -6490 -599 -6466 -597
rect -6410 -599 -6386 -597
rect -6330 -599 -6306 -597
rect -6250 -599 -6226 -597
rect -6170 -599 -6120 -597
rect -6756 -651 -6720 -599
rect -6476 -651 -6466 -599
rect -6410 -651 -6400 -599
rect -6156 -651 -6120 -599
rect -6756 -653 -6706 -651
rect -6650 -653 -6626 -651
rect -6570 -653 -6546 -651
rect -6490 -653 -6466 -651
rect -6410 -653 -6386 -651
rect -6330 -653 -6306 -651
rect -6250 -653 -6226 -651
rect -6170 -653 -6120 -651
rect -6756 -684 -6120 -653
<< via2 >>
rect -6692 103 -6636 105
rect -6612 103 -6556 105
rect -6532 103 -6476 105
rect -6452 103 -6396 105
rect -6372 103 -6316 105
rect -6292 103 -6236 105
rect -6692 51 -6682 103
rect -6682 51 -6636 103
rect -6612 51 -6566 103
rect -6566 51 -6556 103
rect -6532 51 -6502 103
rect -6502 51 -6490 103
rect -6490 51 -6476 103
rect -6452 51 -6438 103
rect -6438 51 -6426 103
rect -6426 51 -6396 103
rect -6372 51 -6362 103
rect -6362 51 -6316 103
rect -6292 51 -6246 103
rect -6246 51 -6236 103
rect -6692 49 -6636 51
rect -6612 49 -6556 51
rect -6532 49 -6476 51
rect -6452 49 -6396 51
rect -6372 49 -6316 51
rect -6292 49 -6236 51
rect -6148 -203 -6092 -202
rect -6148 -255 -6145 -203
rect -6145 -255 -6093 -203
rect -6093 -255 -6092 -203
rect -6148 -258 -6092 -255
rect -5560 -416 -5504 -414
rect -5560 -468 -5558 -416
rect -5558 -468 -5506 -416
rect -5506 -468 -5504 -416
rect -5560 -470 -5504 -468
rect -6706 -599 -6650 -597
rect -6626 -599 -6570 -597
rect -6546 -599 -6490 -597
rect -6466 -599 -6410 -597
rect -6386 -599 -6330 -597
rect -6306 -599 -6250 -597
rect -6226 -599 -6170 -597
rect -6706 -651 -6668 -599
rect -6668 -651 -6656 -599
rect -6656 -651 -6650 -599
rect -6626 -651 -6604 -599
rect -6604 -651 -6592 -599
rect -6592 -651 -6570 -599
rect -6546 -651 -6540 -599
rect -6540 -651 -6528 -599
rect -6528 -651 -6490 -599
rect -6466 -651 -6464 -599
rect -6464 -651 -6412 -599
rect -6412 -651 -6410 -599
rect -6386 -651 -6348 -599
rect -6348 -651 -6336 -599
rect -6336 -651 -6330 -599
rect -6306 -651 -6284 -599
rect -6284 -651 -6272 -599
rect -6272 -651 -6250 -599
rect -6226 -651 -6220 -599
rect -6220 -651 -6208 -599
rect -6208 -651 -6170 -599
rect -6706 -653 -6650 -651
rect -6626 -653 -6570 -651
rect -6546 -653 -6490 -651
rect -6466 -653 -6410 -651
rect -6386 -653 -6330 -651
rect -6306 -653 -6250 -651
rect -6226 -653 -6170 -651
<< metal3 >>
rect -7582 105 -4707 146
rect -7582 49 -6692 105
rect -6636 49 -6612 105
rect -6556 49 -6532 105
rect -6476 49 -6452 105
rect -6396 49 -6372 105
rect -6316 49 -6292 105
rect -6236 49 -4707 105
rect -7582 6 -4707 49
rect -6155 -202 -6085 -195
rect -6155 -258 -6148 -202
rect -6092 -258 -6085 -202
rect -6155 -265 -6085 -258
rect -6150 -412 -6090 -265
rect -5567 -412 -5497 -407
rect -6150 -414 -5497 -412
rect -6150 -470 -5560 -414
rect -5504 -470 -5497 -414
rect -6150 -472 -5497 -470
rect -5567 -477 -5497 -472
rect -7582 -597 -4715 -544
rect -7582 -653 -6706 -597
rect -6650 -653 -6626 -597
rect -6570 -653 -6546 -597
rect -6490 -653 -6466 -597
rect -6410 -653 -6386 -597
rect -6330 -653 -6306 -597
rect -6250 -653 -6226 -597
rect -6170 -653 -4715 -597
rect -7582 -684 -4715 -653
<< labels >>
flabel metal1 s -4588 62 -4588 62 3 FreeSans 400 0 0 0 VOUTH
flabel metal1 s -4602 -652 -4602 -652 3 FreeSans 400 0 0 0 VOUTL
flabel metal2 s -6826 -242 -6826 -242 7 FreeSans 400 0 0 0 R_L
flabel metal1 s -5418 26 -5418 26 3 FreeSans 400 0 0 0 DX_BUF
flabel metal2 s -6814 -148 -6814 -148 7 FreeSans 400 0 0 0 R_H
flabel metal2 s -7456 -326 -7456 -326 7 FreeSans 400 0 0 0 DX
flabel metal2 s -7466 -440 -7466 -440 7 FreeSans 400 0 0 0 VREFL
flabel metal2 s -7446 -2 -7446 -2 5 FreeSans 400 0 0 0 VREFH
flabel metal3 s -7582 -684 -7552 -544 7 FreeSans 600 0 0 0 VSS
flabel metal3 s -7582 6 -7552 146 7 FreeSans 600 0 0 0 VCC
<< end >>
